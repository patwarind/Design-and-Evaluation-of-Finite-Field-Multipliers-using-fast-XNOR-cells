`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Nitin D. Patwari
// 
// Create Date: 20.01.2022 22:23:39
// Design Name: 
// Module Name: CA_233bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CA_233bit(
    a,
    b,
    y
    );

input [232:0] a;
input [232:0] b;

output [464:0] y;



assign y[0] = (a[0] & b[0]);
assign y[1] = (a[1] & b[0])^(a[0] & b[1]);
assign y[2] = (a[2] & b[0])^(a[1] & b[1])^(a[0] & b[2]);
assign y[3] = (a[3] & b[0])^(a[2] & b[1])^(a[1] & b[2])^(a[0] & b[3]);
assign y[4] = (a[4] & b[0])^(a[3] & b[1])^(a[2] & b[2])^(a[1] & b[3])^(a[0] & b[4]);
assign y[5] = (a[5] & b[0])^(a[4] & b[1])^(a[3] & b[2])^(a[2] & b[3])^(a[1] & b[4])^(a[0] & b[5]);
assign y[6] = (a[6] & b[0])^(a[5] & b[1])^(a[4] & b[2])^(a[3] & b[3])^(a[2] & b[4])^(a[1] & b[5])^(a[0] & b[6]);
assign y[7] = (a[7] & b[0])^(a[6] & b[1])^(a[5] & b[2])^(a[4] & b[3])^(a[3] & b[4])^(a[2] & b[5])^(a[1] & b[6])^(a[0] & b[7]);
assign y[8] = (a[8] & b[0])^(a[7] & b[1])^(a[6] & b[2])^(a[5] & b[3])^(a[4] & b[4])^(a[3] & b[5])^(a[2] & b[6])^(a[1] & b[7])^(a[0] & b[8]);
assign y[9] = (a[9] & b[0])^(a[8] & b[1])^(a[7] & b[2])^(a[6] & b[3])^(a[5] & b[4])^(a[4] & b[5])^(a[3] & b[6])^(a[2] & b[7])^(a[1] & b[8])^(a[0] & b[9]);
assign y[10] = (a[10] & b[0])^(a[9] & b[1])^(a[8] & b[2])^(a[7] & b[3])^(a[6] & b[4])^(a[5] & b[5])^(a[4] & b[6])^(a[3] & b[7])^(a[2] & b[8])^(a[1] & b[9])^(a[0] & b[10]);
assign y[11] = (a[11] & b[0])^(a[10] & b[1])^(a[9] & b[2])^(a[8] & b[3])^(a[7] & b[4])^(a[6] & b[5])^(a[5] & b[6])^(a[4] & b[7])^(a[3] & b[8])^(a[2] & b[9])^(a[1] & b[10])^(a[0] & b[11]);
assign y[12] = (a[12] & b[0])^(a[11] & b[1])^(a[10] & b[2])^(a[9] & b[3])^(a[8] & b[4])^(a[7] & b[5])^(a[6] & b[6])^(a[5] & b[7])^(a[4] & b[8])^(a[3] & b[9])^(a[2] & b[10])^(a[1] & b[11])^(a[0] & b[12]);
assign y[13] = (a[13] & b[0])^(a[12] & b[1])^(a[11] & b[2])^(a[10] & b[3])^(a[9] & b[4])^(a[8] & b[5])^(a[7] & b[6])^(a[6] & b[7])^(a[5] & b[8])^(a[4] & b[9])^(a[3] & b[10])^(a[2] & b[11])^(a[1] & b[12])^(a[0] & b[13]);
assign y[14] = (a[14] & b[0])^(a[13] & b[1])^(a[12] & b[2])^(a[11] & b[3])^(a[10] & b[4])^(a[9] & b[5])^(a[8] & b[6])^(a[7] & b[7])^(a[6] & b[8])^(a[5] & b[9])^(a[4] & b[10])^(a[3] & b[11])^(a[2] & b[12])^(a[1] & b[13])^(a[0] & b[14]);
assign y[15] = (a[15] & b[0])^(a[14] & b[1])^(a[13] & b[2])^(a[12] & b[3])^(a[11] & b[4])^(a[10] & b[5])^(a[9] & b[6])^(a[8] & b[7])^(a[7] & b[8])^(a[6] & b[9])^(a[5] & b[10])^(a[4] & b[11])^(a[3] & b[12])^(a[2] & b[13])^(a[1] & b[14])^(a[0] & b[15]);
assign y[16] = (a[16] & b[0])^(a[15] & b[1])^(a[14] & b[2])^(a[13] & b[3])^(a[12] & b[4])^(a[11] & b[5])^(a[10] & b[6])^(a[9] & b[7])^(a[8] & b[8])^(a[7] & b[9])^(a[6] & b[10])^(a[5] & b[11])^(a[4] & b[12])^(a[3] & b[13])^(a[2] & b[14])^(a[1] & b[15])^(a[0] & b[16]);
assign y[17] = (a[17] & b[0])^(a[16] & b[1])^(a[15] & b[2])^(a[14] & b[3])^(a[13] & b[4])^(a[12] & b[5])^(a[11] & b[6])^(a[10] & b[7])^(a[9] & b[8])^(a[8] & b[9])^(a[7] & b[10])^(a[6] & b[11])^(a[5] & b[12])^(a[4] & b[13])^(a[3] & b[14])^(a[2] & b[15])^(a[1] & b[16])^(a[0] & b[17]);
assign y[18] = (a[18] & b[0])^(a[17] & b[1])^(a[16] & b[2])^(a[15] & b[3])^(a[14] & b[4])^(a[13] & b[5])^(a[12] & b[6])^(a[11] & b[7])^(a[10] & b[8])^(a[9] & b[9])^(a[8] & b[10])^(a[7] & b[11])^(a[6] & b[12])^(a[5] & b[13])^(a[4] & b[14])^(a[3] & b[15])^(a[2] & b[16])^(a[1] & b[17])^(a[0] & b[18]);
assign y[19] = (a[19] & b[0])^(a[18] & b[1])^(a[17] & b[2])^(a[16] & b[3])^(a[15] & b[4])^(a[14] & b[5])^(a[13] & b[6])^(a[12] & b[7])^(a[11] & b[8])^(a[10] & b[9])^(a[9] & b[10])^(a[8] & b[11])^(a[7] & b[12])^(a[6] & b[13])^(a[5] & b[14])^(a[4] & b[15])^(a[3] & b[16])^(a[2] & b[17])^(a[1] & b[18])^(a[0] & b[19]);
assign y[20] = (a[20] & b[0])^(a[19] & b[1])^(a[18] & b[2])^(a[17] & b[3])^(a[16] & b[4])^(a[15] & b[5])^(a[14] & b[6])^(a[13] & b[7])^(a[12] & b[8])^(a[11] & b[9])^(a[10] & b[10])^(a[9] & b[11])^(a[8] & b[12])^(a[7] & b[13])^(a[6] & b[14])^(a[5] & b[15])^(a[4] & b[16])^(a[3] & b[17])^(a[2] & b[18])^(a[1] & b[19])^(a[0] & b[20]);
assign y[21] = (a[21] & b[0])^(a[20] & b[1])^(a[19] & b[2])^(a[18] & b[3])^(a[17] & b[4])^(a[16] & b[5])^(a[15] & b[6])^(a[14] & b[7])^(a[13] & b[8])^(a[12] & b[9])^(a[11] & b[10])^(a[10] & b[11])^(a[9] & b[12])^(a[8] & b[13])^(a[7] & b[14])^(a[6] & b[15])^(a[5] & b[16])^(a[4] & b[17])^(a[3] & b[18])^(a[2] & b[19])^(a[1] & b[20])^(a[0] & b[21]);
assign y[22] = (a[22] & b[0])^(a[21] & b[1])^(a[20] & b[2])^(a[19] & b[3])^(a[18] & b[4])^(a[17] & b[5])^(a[16] & b[6])^(a[15] & b[7])^(a[14] & b[8])^(a[13] & b[9])^(a[12] & b[10])^(a[11] & b[11])^(a[10] & b[12])^(a[9] & b[13])^(a[8] & b[14])^(a[7] & b[15])^(a[6] & b[16])^(a[5] & b[17])^(a[4] & b[18])^(a[3] & b[19])^(a[2] & b[20])^(a[1] & b[21])^(a[0] & b[22]);
assign y[23] = (a[23] & b[0])^(a[22] & b[1])^(a[21] & b[2])^(a[20] & b[3])^(a[19] & b[4])^(a[18] & b[5])^(a[17] & b[6])^(a[16] & b[7])^(a[15] & b[8])^(a[14] & b[9])^(a[13] & b[10])^(a[12] & b[11])^(a[11] & b[12])^(a[10] & b[13])^(a[9] & b[14])^(a[8] & b[15])^(a[7] & b[16])^(a[6] & b[17])^(a[5] & b[18])^(a[4] & b[19])^(a[3] & b[20])^(a[2] & b[21])^(a[1] & b[22])^(a[0] & b[23]);
assign y[24] = (a[24] & b[0])^(a[23] & b[1])^(a[22] & b[2])^(a[21] & b[3])^(a[20] & b[4])^(a[19] & b[5])^(a[18] & b[6])^(a[17] & b[7])^(a[16] & b[8])^(a[15] & b[9])^(a[14] & b[10])^(a[13] & b[11])^(a[12] & b[12])^(a[11] & b[13])^(a[10] & b[14])^(a[9] & b[15])^(a[8] & b[16])^(a[7] & b[17])^(a[6] & b[18])^(a[5] & b[19])^(a[4] & b[20])^(a[3] & b[21])^(a[2] & b[22])^(a[1] & b[23])^(a[0] & b[24]);
assign y[25] = (a[25] & b[0])^(a[24] & b[1])^(a[23] & b[2])^(a[22] & b[3])^(a[21] & b[4])^(a[20] & b[5])^(a[19] & b[6])^(a[18] & b[7])^(a[17] & b[8])^(a[16] & b[9])^(a[15] & b[10])^(a[14] & b[11])^(a[13] & b[12])^(a[12] & b[13])^(a[11] & b[14])^(a[10] & b[15])^(a[9] & b[16])^(a[8] & b[17])^(a[7] & b[18])^(a[6] & b[19])^(a[5] & b[20])^(a[4] & b[21])^(a[3] & b[22])^(a[2] & b[23])^(a[1] & b[24])^(a[0] & b[25]);
assign y[26] = (a[26] & b[0])^(a[25] & b[1])^(a[24] & b[2])^(a[23] & b[3])^(a[22] & b[4])^(a[21] & b[5])^(a[20] & b[6])^(a[19] & b[7])^(a[18] & b[8])^(a[17] & b[9])^(a[16] & b[10])^(a[15] & b[11])^(a[14] & b[12])^(a[13] & b[13])^(a[12] & b[14])^(a[11] & b[15])^(a[10] & b[16])^(a[9] & b[17])^(a[8] & b[18])^(a[7] & b[19])^(a[6] & b[20])^(a[5] & b[21])^(a[4] & b[22])^(a[3] & b[23])^(a[2] & b[24])^(a[1] & b[25])^(a[0] & b[26]);
assign y[27] = (a[27] & b[0])^(a[26] & b[1])^(a[25] & b[2])^(a[24] & b[3])^(a[23] & b[4])^(a[22] & b[5])^(a[21] & b[6])^(a[20] & b[7])^(a[19] & b[8])^(a[18] & b[9])^(a[17] & b[10])^(a[16] & b[11])^(a[15] & b[12])^(a[14] & b[13])^(a[13] & b[14])^(a[12] & b[15])^(a[11] & b[16])^(a[10] & b[17])^(a[9] & b[18])^(a[8] & b[19])^(a[7] & b[20])^(a[6] & b[21])^(a[5] & b[22])^(a[4] & b[23])^(a[3] & b[24])^(a[2] & b[25])^(a[1] & b[26])^(a[0] & b[27]);
assign y[28] = (a[28] & b[0])^(a[27] & b[1])^(a[26] & b[2])^(a[25] & b[3])^(a[24] & b[4])^(a[23] & b[5])^(a[22] & b[6])^(a[21] & b[7])^(a[20] & b[8])^(a[19] & b[9])^(a[18] & b[10])^(a[17] & b[11])^(a[16] & b[12])^(a[15] & b[13])^(a[14] & b[14])^(a[13] & b[15])^(a[12] & b[16])^(a[11] & b[17])^(a[10] & b[18])^(a[9] & b[19])^(a[8] & b[20])^(a[7] & b[21])^(a[6] & b[22])^(a[5] & b[23])^(a[4] & b[24])^(a[3] & b[25])^(a[2] & b[26])^(a[1] & b[27])^(a[0] & b[28]);
assign y[29] = (a[29] & b[0])^(a[28] & b[1])^(a[27] & b[2])^(a[26] & b[3])^(a[25] & b[4])^(a[24] & b[5])^(a[23] & b[6])^(a[22] & b[7])^(a[21] & b[8])^(a[20] & b[9])^(a[19] & b[10])^(a[18] & b[11])^(a[17] & b[12])^(a[16] & b[13])^(a[15] & b[14])^(a[14] & b[15])^(a[13] & b[16])^(a[12] & b[17])^(a[11] & b[18])^(a[10] & b[19])^(a[9] & b[20])^(a[8] & b[21])^(a[7] & b[22])^(a[6] & b[23])^(a[5] & b[24])^(a[4] & b[25])^(a[3] & b[26])^(a[2] & b[27])^(a[1] & b[28])^(a[0] & b[29]);
assign y[30] = (a[30] & b[0])^(a[29] & b[1])^(a[28] & b[2])^(a[27] & b[3])^(a[26] & b[4])^(a[25] & b[5])^(a[24] & b[6])^(a[23] & b[7])^(a[22] & b[8])^(a[21] & b[9])^(a[20] & b[10])^(a[19] & b[11])^(a[18] & b[12])^(a[17] & b[13])^(a[16] & b[14])^(a[15] & b[15])^(a[14] & b[16])^(a[13] & b[17])^(a[12] & b[18])^(a[11] & b[19])^(a[10] & b[20])^(a[9] & b[21])^(a[8] & b[22])^(a[7] & b[23])^(a[6] & b[24])^(a[5] & b[25])^(a[4] & b[26])^(a[3] & b[27])^(a[2] & b[28])^(a[1] & b[29])^(a[0] & b[30]);
assign y[31] = (a[31] & b[0])^(a[30] & b[1])^(a[29] & b[2])^(a[28] & b[3])^(a[27] & b[4])^(a[26] & b[5])^(a[25] & b[6])^(a[24] & b[7])^(a[23] & b[8])^(a[22] & b[9])^(a[21] & b[10])^(a[20] & b[11])^(a[19] & b[12])^(a[18] & b[13])^(a[17] & b[14])^(a[16] & b[15])^(a[15] & b[16])^(a[14] & b[17])^(a[13] & b[18])^(a[12] & b[19])^(a[11] & b[20])^(a[10] & b[21])^(a[9] & b[22])^(a[8] & b[23])^(a[7] & b[24])^(a[6] & b[25])^(a[5] & b[26])^(a[4] & b[27])^(a[3] & b[28])^(a[2] & b[29])^(a[1] & b[30])^(a[0] & b[31]);
assign y[32] = (a[32] & b[0])^(a[31] & b[1])^(a[30] & b[2])^(a[29] & b[3])^(a[28] & b[4])^(a[27] & b[5])^(a[26] & b[6])^(a[25] & b[7])^(a[24] & b[8])^(a[23] & b[9])^(a[22] & b[10])^(a[21] & b[11])^(a[20] & b[12])^(a[19] & b[13])^(a[18] & b[14])^(a[17] & b[15])^(a[16] & b[16])^(a[15] & b[17])^(a[14] & b[18])^(a[13] & b[19])^(a[12] & b[20])^(a[11] & b[21])^(a[10] & b[22])^(a[9] & b[23])^(a[8] & b[24])^(a[7] & b[25])^(a[6] & b[26])^(a[5] & b[27])^(a[4] & b[28])^(a[3] & b[29])^(a[2] & b[30])^(a[1] & b[31])^(a[0] & b[32]);
assign y[33] = (a[33] & b[0])^(a[32] & b[1])^(a[31] & b[2])^(a[30] & b[3])^(a[29] & b[4])^(a[28] & b[5])^(a[27] & b[6])^(a[26] & b[7])^(a[25] & b[8])^(a[24] & b[9])^(a[23] & b[10])^(a[22] & b[11])^(a[21] & b[12])^(a[20] & b[13])^(a[19] & b[14])^(a[18] & b[15])^(a[17] & b[16])^(a[16] & b[17])^(a[15] & b[18])^(a[14] & b[19])^(a[13] & b[20])^(a[12] & b[21])^(a[11] & b[22])^(a[10] & b[23])^(a[9] & b[24])^(a[8] & b[25])^(a[7] & b[26])^(a[6] & b[27])^(a[5] & b[28])^(a[4] & b[29])^(a[3] & b[30])^(a[2] & b[31])^(a[1] & b[32])^(a[0] & b[33]);
assign y[34] = (a[34] & b[0])^(a[33] & b[1])^(a[32] & b[2])^(a[31] & b[3])^(a[30] & b[4])^(a[29] & b[5])^(a[28] & b[6])^(a[27] & b[7])^(a[26] & b[8])^(a[25] & b[9])^(a[24] & b[10])^(a[23] & b[11])^(a[22] & b[12])^(a[21] & b[13])^(a[20] & b[14])^(a[19] & b[15])^(a[18] & b[16])^(a[17] & b[17])^(a[16] & b[18])^(a[15] & b[19])^(a[14] & b[20])^(a[13] & b[21])^(a[12] & b[22])^(a[11] & b[23])^(a[10] & b[24])^(a[9] & b[25])^(a[8] & b[26])^(a[7] & b[27])^(a[6] & b[28])^(a[5] & b[29])^(a[4] & b[30])^(a[3] & b[31])^(a[2] & b[32])^(a[1] & b[33])^(a[0] & b[34]);
assign y[35] = (a[35] & b[0])^(a[34] & b[1])^(a[33] & b[2])^(a[32] & b[3])^(a[31] & b[4])^(a[30] & b[5])^(a[29] & b[6])^(a[28] & b[7])^(a[27] & b[8])^(a[26] & b[9])^(a[25] & b[10])^(a[24] & b[11])^(a[23] & b[12])^(a[22] & b[13])^(a[21] & b[14])^(a[20] & b[15])^(a[19] & b[16])^(a[18] & b[17])^(a[17] & b[18])^(a[16] & b[19])^(a[15] & b[20])^(a[14] & b[21])^(a[13] & b[22])^(a[12] & b[23])^(a[11] & b[24])^(a[10] & b[25])^(a[9] & b[26])^(a[8] & b[27])^(a[7] & b[28])^(a[6] & b[29])^(a[5] & b[30])^(a[4] & b[31])^(a[3] & b[32])^(a[2] & b[33])^(a[1] & b[34])^(a[0] & b[35]);
assign y[36] = (a[36] & b[0])^(a[35] & b[1])^(a[34] & b[2])^(a[33] & b[3])^(a[32] & b[4])^(a[31] & b[5])^(a[30] & b[6])^(a[29] & b[7])^(a[28] & b[8])^(a[27] & b[9])^(a[26] & b[10])^(a[25] & b[11])^(a[24] & b[12])^(a[23] & b[13])^(a[22] & b[14])^(a[21] & b[15])^(a[20] & b[16])^(a[19] & b[17])^(a[18] & b[18])^(a[17] & b[19])^(a[16] & b[20])^(a[15] & b[21])^(a[14] & b[22])^(a[13] & b[23])^(a[12] & b[24])^(a[11] & b[25])^(a[10] & b[26])^(a[9] & b[27])^(a[8] & b[28])^(a[7] & b[29])^(a[6] & b[30])^(a[5] & b[31])^(a[4] & b[32])^(a[3] & b[33])^(a[2] & b[34])^(a[1] & b[35])^(a[0] & b[36]);
assign y[37] = (a[37] & b[0])^(a[36] & b[1])^(a[35] & b[2])^(a[34] & b[3])^(a[33] & b[4])^(a[32] & b[5])^(a[31] & b[6])^(a[30] & b[7])^(a[29] & b[8])^(a[28] & b[9])^(a[27] & b[10])^(a[26] & b[11])^(a[25] & b[12])^(a[24] & b[13])^(a[23] & b[14])^(a[22] & b[15])^(a[21] & b[16])^(a[20] & b[17])^(a[19] & b[18])^(a[18] & b[19])^(a[17] & b[20])^(a[16] & b[21])^(a[15] & b[22])^(a[14] & b[23])^(a[13] & b[24])^(a[12] & b[25])^(a[11] & b[26])^(a[10] & b[27])^(a[9] & b[28])^(a[8] & b[29])^(a[7] & b[30])^(a[6] & b[31])^(a[5] & b[32])^(a[4] & b[33])^(a[3] & b[34])^(a[2] & b[35])^(a[1] & b[36])^(a[0] & b[37]);
assign y[38] = (a[38] & b[0])^(a[37] & b[1])^(a[36] & b[2])^(a[35] & b[3])^(a[34] & b[4])^(a[33] & b[5])^(a[32] & b[6])^(a[31] & b[7])^(a[30] & b[8])^(a[29] & b[9])^(a[28] & b[10])^(a[27] & b[11])^(a[26] & b[12])^(a[25] & b[13])^(a[24] & b[14])^(a[23] & b[15])^(a[22] & b[16])^(a[21] & b[17])^(a[20] & b[18])^(a[19] & b[19])^(a[18] & b[20])^(a[17] & b[21])^(a[16] & b[22])^(a[15] & b[23])^(a[14] & b[24])^(a[13] & b[25])^(a[12] & b[26])^(a[11] & b[27])^(a[10] & b[28])^(a[9] & b[29])^(a[8] & b[30])^(a[7] & b[31])^(a[6] & b[32])^(a[5] & b[33])^(a[4] & b[34])^(a[3] & b[35])^(a[2] & b[36])^(a[1] & b[37])^(a[0] & b[38]);
assign y[39] = (a[39] & b[0])^(a[38] & b[1])^(a[37] & b[2])^(a[36] & b[3])^(a[35] & b[4])^(a[34] & b[5])^(a[33] & b[6])^(a[32] & b[7])^(a[31] & b[8])^(a[30] & b[9])^(a[29] & b[10])^(a[28] & b[11])^(a[27] & b[12])^(a[26] & b[13])^(a[25] & b[14])^(a[24] & b[15])^(a[23] & b[16])^(a[22] & b[17])^(a[21] & b[18])^(a[20] & b[19])^(a[19] & b[20])^(a[18] & b[21])^(a[17] & b[22])^(a[16] & b[23])^(a[15] & b[24])^(a[14] & b[25])^(a[13] & b[26])^(a[12] & b[27])^(a[11] & b[28])^(a[10] & b[29])^(a[9] & b[30])^(a[8] & b[31])^(a[7] & b[32])^(a[6] & b[33])^(a[5] & b[34])^(a[4] & b[35])^(a[3] & b[36])^(a[2] & b[37])^(a[1] & b[38])^(a[0] & b[39]);
assign y[40] = (a[40] & b[0])^(a[39] & b[1])^(a[38] & b[2])^(a[37] & b[3])^(a[36] & b[4])^(a[35] & b[5])^(a[34] & b[6])^(a[33] & b[7])^(a[32] & b[8])^(a[31] & b[9])^(a[30] & b[10])^(a[29] & b[11])^(a[28] & b[12])^(a[27] & b[13])^(a[26] & b[14])^(a[25] & b[15])^(a[24] & b[16])^(a[23] & b[17])^(a[22] & b[18])^(a[21] & b[19])^(a[20] & b[20])^(a[19] & b[21])^(a[18] & b[22])^(a[17] & b[23])^(a[16] & b[24])^(a[15] & b[25])^(a[14] & b[26])^(a[13] & b[27])^(a[12] & b[28])^(a[11] & b[29])^(a[10] & b[30])^(a[9] & b[31])^(a[8] & b[32])^(a[7] & b[33])^(a[6] & b[34])^(a[5] & b[35])^(a[4] & b[36])^(a[3] & b[37])^(a[2] & b[38])^(a[1] & b[39])^(a[0] & b[40]);
assign y[41] = (a[41] & b[0])^(a[40] & b[1])^(a[39] & b[2])^(a[38] & b[3])^(a[37] & b[4])^(a[36] & b[5])^(a[35] & b[6])^(a[34] & b[7])^(a[33] & b[8])^(a[32] & b[9])^(a[31] & b[10])^(a[30] & b[11])^(a[29] & b[12])^(a[28] & b[13])^(a[27] & b[14])^(a[26] & b[15])^(a[25] & b[16])^(a[24] & b[17])^(a[23] & b[18])^(a[22] & b[19])^(a[21] & b[20])^(a[20] & b[21])^(a[19] & b[22])^(a[18] & b[23])^(a[17] & b[24])^(a[16] & b[25])^(a[15] & b[26])^(a[14] & b[27])^(a[13] & b[28])^(a[12] & b[29])^(a[11] & b[30])^(a[10] & b[31])^(a[9] & b[32])^(a[8] & b[33])^(a[7] & b[34])^(a[6] & b[35])^(a[5] & b[36])^(a[4] & b[37])^(a[3] & b[38])^(a[2] & b[39])^(a[1] & b[40])^(a[0] & b[41]);
assign y[42] = (a[42] & b[0])^(a[41] & b[1])^(a[40] & b[2])^(a[39] & b[3])^(a[38] & b[4])^(a[37] & b[5])^(a[36] & b[6])^(a[35] & b[7])^(a[34] & b[8])^(a[33] & b[9])^(a[32] & b[10])^(a[31] & b[11])^(a[30] & b[12])^(a[29] & b[13])^(a[28] & b[14])^(a[27] & b[15])^(a[26] & b[16])^(a[25] & b[17])^(a[24] & b[18])^(a[23] & b[19])^(a[22] & b[20])^(a[21] & b[21])^(a[20] & b[22])^(a[19] & b[23])^(a[18] & b[24])^(a[17] & b[25])^(a[16] & b[26])^(a[15] & b[27])^(a[14] & b[28])^(a[13] & b[29])^(a[12] & b[30])^(a[11] & b[31])^(a[10] & b[32])^(a[9] & b[33])^(a[8] & b[34])^(a[7] & b[35])^(a[6] & b[36])^(a[5] & b[37])^(a[4] & b[38])^(a[3] & b[39])^(a[2] & b[40])^(a[1] & b[41])^(a[0] & b[42]);
assign y[43] = (a[43] & b[0])^(a[42] & b[1])^(a[41] & b[2])^(a[40] & b[3])^(a[39] & b[4])^(a[38] & b[5])^(a[37] & b[6])^(a[36] & b[7])^(a[35] & b[8])^(a[34] & b[9])^(a[33] & b[10])^(a[32] & b[11])^(a[31] & b[12])^(a[30] & b[13])^(a[29] & b[14])^(a[28] & b[15])^(a[27] & b[16])^(a[26] & b[17])^(a[25] & b[18])^(a[24] & b[19])^(a[23] & b[20])^(a[22] & b[21])^(a[21] & b[22])^(a[20] & b[23])^(a[19] & b[24])^(a[18] & b[25])^(a[17] & b[26])^(a[16] & b[27])^(a[15] & b[28])^(a[14] & b[29])^(a[13] & b[30])^(a[12] & b[31])^(a[11] & b[32])^(a[10] & b[33])^(a[9] & b[34])^(a[8] & b[35])^(a[7] & b[36])^(a[6] & b[37])^(a[5] & b[38])^(a[4] & b[39])^(a[3] & b[40])^(a[2] & b[41])^(a[1] & b[42])^(a[0] & b[43]);
assign y[44] = (a[44] & b[0])^(a[43] & b[1])^(a[42] & b[2])^(a[41] & b[3])^(a[40] & b[4])^(a[39] & b[5])^(a[38] & b[6])^(a[37] & b[7])^(a[36] & b[8])^(a[35] & b[9])^(a[34] & b[10])^(a[33] & b[11])^(a[32] & b[12])^(a[31] & b[13])^(a[30] & b[14])^(a[29] & b[15])^(a[28] & b[16])^(a[27] & b[17])^(a[26] & b[18])^(a[25] & b[19])^(a[24] & b[20])^(a[23] & b[21])^(a[22] & b[22])^(a[21] & b[23])^(a[20] & b[24])^(a[19] & b[25])^(a[18] & b[26])^(a[17] & b[27])^(a[16] & b[28])^(a[15] & b[29])^(a[14] & b[30])^(a[13] & b[31])^(a[12] & b[32])^(a[11] & b[33])^(a[10] & b[34])^(a[9] & b[35])^(a[8] & b[36])^(a[7] & b[37])^(a[6] & b[38])^(a[5] & b[39])^(a[4] & b[40])^(a[3] & b[41])^(a[2] & b[42])^(a[1] & b[43])^(a[0] & b[44]);
assign y[45] = (a[45] & b[0])^(a[44] & b[1])^(a[43] & b[2])^(a[42] & b[3])^(a[41] & b[4])^(a[40] & b[5])^(a[39] & b[6])^(a[38] & b[7])^(a[37] & b[8])^(a[36] & b[9])^(a[35] & b[10])^(a[34] & b[11])^(a[33] & b[12])^(a[32] & b[13])^(a[31] & b[14])^(a[30] & b[15])^(a[29] & b[16])^(a[28] & b[17])^(a[27] & b[18])^(a[26] & b[19])^(a[25] & b[20])^(a[24] & b[21])^(a[23] & b[22])^(a[22] & b[23])^(a[21] & b[24])^(a[20] & b[25])^(a[19] & b[26])^(a[18] & b[27])^(a[17] & b[28])^(a[16] & b[29])^(a[15] & b[30])^(a[14] & b[31])^(a[13] & b[32])^(a[12] & b[33])^(a[11] & b[34])^(a[10] & b[35])^(a[9] & b[36])^(a[8] & b[37])^(a[7] & b[38])^(a[6] & b[39])^(a[5] & b[40])^(a[4] & b[41])^(a[3] & b[42])^(a[2] & b[43])^(a[1] & b[44])^(a[0] & b[45]);
assign y[46] = (a[46] & b[0])^(a[45] & b[1])^(a[44] & b[2])^(a[43] & b[3])^(a[42] & b[4])^(a[41] & b[5])^(a[40] & b[6])^(a[39] & b[7])^(a[38] & b[8])^(a[37] & b[9])^(a[36] & b[10])^(a[35] & b[11])^(a[34] & b[12])^(a[33] & b[13])^(a[32] & b[14])^(a[31] & b[15])^(a[30] & b[16])^(a[29] & b[17])^(a[28] & b[18])^(a[27] & b[19])^(a[26] & b[20])^(a[25] & b[21])^(a[24] & b[22])^(a[23] & b[23])^(a[22] & b[24])^(a[21] & b[25])^(a[20] & b[26])^(a[19] & b[27])^(a[18] & b[28])^(a[17] & b[29])^(a[16] & b[30])^(a[15] & b[31])^(a[14] & b[32])^(a[13] & b[33])^(a[12] & b[34])^(a[11] & b[35])^(a[10] & b[36])^(a[9] & b[37])^(a[8] & b[38])^(a[7] & b[39])^(a[6] & b[40])^(a[5] & b[41])^(a[4] & b[42])^(a[3] & b[43])^(a[2] & b[44])^(a[1] & b[45])^(a[0] & b[46]);
assign y[47] = (a[47] & b[0])^(a[46] & b[1])^(a[45] & b[2])^(a[44] & b[3])^(a[43] & b[4])^(a[42] & b[5])^(a[41] & b[6])^(a[40] & b[7])^(a[39] & b[8])^(a[38] & b[9])^(a[37] & b[10])^(a[36] & b[11])^(a[35] & b[12])^(a[34] & b[13])^(a[33] & b[14])^(a[32] & b[15])^(a[31] & b[16])^(a[30] & b[17])^(a[29] & b[18])^(a[28] & b[19])^(a[27] & b[20])^(a[26] & b[21])^(a[25] & b[22])^(a[24] & b[23])^(a[23] & b[24])^(a[22] & b[25])^(a[21] & b[26])^(a[20] & b[27])^(a[19] & b[28])^(a[18] & b[29])^(a[17] & b[30])^(a[16] & b[31])^(a[15] & b[32])^(a[14] & b[33])^(a[13] & b[34])^(a[12] & b[35])^(a[11] & b[36])^(a[10] & b[37])^(a[9] & b[38])^(a[8] & b[39])^(a[7] & b[40])^(a[6] & b[41])^(a[5] & b[42])^(a[4] & b[43])^(a[3] & b[44])^(a[2] & b[45])^(a[1] & b[46])^(a[0] & b[47]);
assign y[48] = (a[48] & b[0])^(a[47] & b[1])^(a[46] & b[2])^(a[45] & b[3])^(a[44] & b[4])^(a[43] & b[5])^(a[42] & b[6])^(a[41] & b[7])^(a[40] & b[8])^(a[39] & b[9])^(a[38] & b[10])^(a[37] & b[11])^(a[36] & b[12])^(a[35] & b[13])^(a[34] & b[14])^(a[33] & b[15])^(a[32] & b[16])^(a[31] & b[17])^(a[30] & b[18])^(a[29] & b[19])^(a[28] & b[20])^(a[27] & b[21])^(a[26] & b[22])^(a[25] & b[23])^(a[24] & b[24])^(a[23] & b[25])^(a[22] & b[26])^(a[21] & b[27])^(a[20] & b[28])^(a[19] & b[29])^(a[18] & b[30])^(a[17] & b[31])^(a[16] & b[32])^(a[15] & b[33])^(a[14] & b[34])^(a[13] & b[35])^(a[12] & b[36])^(a[11] & b[37])^(a[10] & b[38])^(a[9] & b[39])^(a[8] & b[40])^(a[7] & b[41])^(a[6] & b[42])^(a[5] & b[43])^(a[4] & b[44])^(a[3] & b[45])^(a[2] & b[46])^(a[1] & b[47])^(a[0] & b[48]);
assign y[49] = (a[49] & b[0])^(a[48] & b[1])^(a[47] & b[2])^(a[46] & b[3])^(a[45] & b[4])^(a[44] & b[5])^(a[43] & b[6])^(a[42] & b[7])^(a[41] & b[8])^(a[40] & b[9])^(a[39] & b[10])^(a[38] & b[11])^(a[37] & b[12])^(a[36] & b[13])^(a[35] & b[14])^(a[34] & b[15])^(a[33] & b[16])^(a[32] & b[17])^(a[31] & b[18])^(a[30] & b[19])^(a[29] & b[20])^(a[28] & b[21])^(a[27] & b[22])^(a[26] & b[23])^(a[25] & b[24])^(a[24] & b[25])^(a[23] & b[26])^(a[22] & b[27])^(a[21] & b[28])^(a[20] & b[29])^(a[19] & b[30])^(a[18] & b[31])^(a[17] & b[32])^(a[16] & b[33])^(a[15] & b[34])^(a[14] & b[35])^(a[13] & b[36])^(a[12] & b[37])^(a[11] & b[38])^(a[10] & b[39])^(a[9] & b[40])^(a[8] & b[41])^(a[7] & b[42])^(a[6] & b[43])^(a[5] & b[44])^(a[4] & b[45])^(a[3] & b[46])^(a[2] & b[47])^(a[1] & b[48])^(a[0] & b[49]);
assign y[50] = (a[50] & b[0])^(a[49] & b[1])^(a[48] & b[2])^(a[47] & b[3])^(a[46] & b[4])^(a[45] & b[5])^(a[44] & b[6])^(a[43] & b[7])^(a[42] & b[8])^(a[41] & b[9])^(a[40] & b[10])^(a[39] & b[11])^(a[38] & b[12])^(a[37] & b[13])^(a[36] & b[14])^(a[35] & b[15])^(a[34] & b[16])^(a[33] & b[17])^(a[32] & b[18])^(a[31] & b[19])^(a[30] & b[20])^(a[29] & b[21])^(a[28] & b[22])^(a[27] & b[23])^(a[26] & b[24])^(a[25] & b[25])^(a[24] & b[26])^(a[23] & b[27])^(a[22] & b[28])^(a[21] & b[29])^(a[20] & b[30])^(a[19] & b[31])^(a[18] & b[32])^(a[17] & b[33])^(a[16] & b[34])^(a[15] & b[35])^(a[14] & b[36])^(a[13] & b[37])^(a[12] & b[38])^(a[11] & b[39])^(a[10] & b[40])^(a[9] & b[41])^(a[8] & b[42])^(a[7] & b[43])^(a[6] & b[44])^(a[5] & b[45])^(a[4] & b[46])^(a[3] & b[47])^(a[2] & b[48])^(a[1] & b[49])^(a[0] & b[50]);
assign y[51] = (a[51] & b[0])^(a[50] & b[1])^(a[49] & b[2])^(a[48] & b[3])^(a[47] & b[4])^(a[46] & b[5])^(a[45] & b[6])^(a[44] & b[7])^(a[43] & b[8])^(a[42] & b[9])^(a[41] & b[10])^(a[40] & b[11])^(a[39] & b[12])^(a[38] & b[13])^(a[37] & b[14])^(a[36] & b[15])^(a[35] & b[16])^(a[34] & b[17])^(a[33] & b[18])^(a[32] & b[19])^(a[31] & b[20])^(a[30] & b[21])^(a[29] & b[22])^(a[28] & b[23])^(a[27] & b[24])^(a[26] & b[25])^(a[25] & b[26])^(a[24] & b[27])^(a[23] & b[28])^(a[22] & b[29])^(a[21] & b[30])^(a[20] & b[31])^(a[19] & b[32])^(a[18] & b[33])^(a[17] & b[34])^(a[16] & b[35])^(a[15] & b[36])^(a[14] & b[37])^(a[13] & b[38])^(a[12] & b[39])^(a[11] & b[40])^(a[10] & b[41])^(a[9] & b[42])^(a[8] & b[43])^(a[7] & b[44])^(a[6] & b[45])^(a[5] & b[46])^(a[4] & b[47])^(a[3] & b[48])^(a[2] & b[49])^(a[1] & b[50])^(a[0] & b[51]);
assign y[52] = (a[52] & b[0])^(a[51] & b[1])^(a[50] & b[2])^(a[49] & b[3])^(a[48] & b[4])^(a[47] & b[5])^(a[46] & b[6])^(a[45] & b[7])^(a[44] & b[8])^(a[43] & b[9])^(a[42] & b[10])^(a[41] & b[11])^(a[40] & b[12])^(a[39] & b[13])^(a[38] & b[14])^(a[37] & b[15])^(a[36] & b[16])^(a[35] & b[17])^(a[34] & b[18])^(a[33] & b[19])^(a[32] & b[20])^(a[31] & b[21])^(a[30] & b[22])^(a[29] & b[23])^(a[28] & b[24])^(a[27] & b[25])^(a[26] & b[26])^(a[25] & b[27])^(a[24] & b[28])^(a[23] & b[29])^(a[22] & b[30])^(a[21] & b[31])^(a[20] & b[32])^(a[19] & b[33])^(a[18] & b[34])^(a[17] & b[35])^(a[16] & b[36])^(a[15] & b[37])^(a[14] & b[38])^(a[13] & b[39])^(a[12] & b[40])^(a[11] & b[41])^(a[10] & b[42])^(a[9] & b[43])^(a[8] & b[44])^(a[7] & b[45])^(a[6] & b[46])^(a[5] & b[47])^(a[4] & b[48])^(a[3] & b[49])^(a[2] & b[50])^(a[1] & b[51])^(a[0] & b[52]);
assign y[53] = (a[53] & b[0])^(a[52] & b[1])^(a[51] & b[2])^(a[50] & b[3])^(a[49] & b[4])^(a[48] & b[5])^(a[47] & b[6])^(a[46] & b[7])^(a[45] & b[8])^(a[44] & b[9])^(a[43] & b[10])^(a[42] & b[11])^(a[41] & b[12])^(a[40] & b[13])^(a[39] & b[14])^(a[38] & b[15])^(a[37] & b[16])^(a[36] & b[17])^(a[35] & b[18])^(a[34] & b[19])^(a[33] & b[20])^(a[32] & b[21])^(a[31] & b[22])^(a[30] & b[23])^(a[29] & b[24])^(a[28] & b[25])^(a[27] & b[26])^(a[26] & b[27])^(a[25] & b[28])^(a[24] & b[29])^(a[23] & b[30])^(a[22] & b[31])^(a[21] & b[32])^(a[20] & b[33])^(a[19] & b[34])^(a[18] & b[35])^(a[17] & b[36])^(a[16] & b[37])^(a[15] & b[38])^(a[14] & b[39])^(a[13] & b[40])^(a[12] & b[41])^(a[11] & b[42])^(a[10] & b[43])^(a[9] & b[44])^(a[8] & b[45])^(a[7] & b[46])^(a[6] & b[47])^(a[5] & b[48])^(a[4] & b[49])^(a[3] & b[50])^(a[2] & b[51])^(a[1] & b[52])^(a[0] & b[53]);
assign y[54] = (a[54] & b[0])^(a[53] & b[1])^(a[52] & b[2])^(a[51] & b[3])^(a[50] & b[4])^(a[49] & b[5])^(a[48] & b[6])^(a[47] & b[7])^(a[46] & b[8])^(a[45] & b[9])^(a[44] & b[10])^(a[43] & b[11])^(a[42] & b[12])^(a[41] & b[13])^(a[40] & b[14])^(a[39] & b[15])^(a[38] & b[16])^(a[37] & b[17])^(a[36] & b[18])^(a[35] & b[19])^(a[34] & b[20])^(a[33] & b[21])^(a[32] & b[22])^(a[31] & b[23])^(a[30] & b[24])^(a[29] & b[25])^(a[28] & b[26])^(a[27] & b[27])^(a[26] & b[28])^(a[25] & b[29])^(a[24] & b[30])^(a[23] & b[31])^(a[22] & b[32])^(a[21] & b[33])^(a[20] & b[34])^(a[19] & b[35])^(a[18] & b[36])^(a[17] & b[37])^(a[16] & b[38])^(a[15] & b[39])^(a[14] & b[40])^(a[13] & b[41])^(a[12] & b[42])^(a[11] & b[43])^(a[10] & b[44])^(a[9] & b[45])^(a[8] & b[46])^(a[7] & b[47])^(a[6] & b[48])^(a[5] & b[49])^(a[4] & b[50])^(a[3] & b[51])^(a[2] & b[52])^(a[1] & b[53])^(a[0] & b[54]);
assign y[55] = (a[55] & b[0])^(a[54] & b[1])^(a[53] & b[2])^(a[52] & b[3])^(a[51] & b[4])^(a[50] & b[5])^(a[49] & b[6])^(a[48] & b[7])^(a[47] & b[8])^(a[46] & b[9])^(a[45] & b[10])^(a[44] & b[11])^(a[43] & b[12])^(a[42] & b[13])^(a[41] & b[14])^(a[40] & b[15])^(a[39] & b[16])^(a[38] & b[17])^(a[37] & b[18])^(a[36] & b[19])^(a[35] & b[20])^(a[34] & b[21])^(a[33] & b[22])^(a[32] & b[23])^(a[31] & b[24])^(a[30] & b[25])^(a[29] & b[26])^(a[28] & b[27])^(a[27] & b[28])^(a[26] & b[29])^(a[25] & b[30])^(a[24] & b[31])^(a[23] & b[32])^(a[22] & b[33])^(a[21] & b[34])^(a[20] & b[35])^(a[19] & b[36])^(a[18] & b[37])^(a[17] & b[38])^(a[16] & b[39])^(a[15] & b[40])^(a[14] & b[41])^(a[13] & b[42])^(a[12] & b[43])^(a[11] & b[44])^(a[10] & b[45])^(a[9] & b[46])^(a[8] & b[47])^(a[7] & b[48])^(a[6] & b[49])^(a[5] & b[50])^(a[4] & b[51])^(a[3] & b[52])^(a[2] & b[53])^(a[1] & b[54])^(a[0] & b[55]);
assign y[56] = (a[56] & b[0])^(a[55] & b[1])^(a[54] & b[2])^(a[53] & b[3])^(a[52] & b[4])^(a[51] & b[5])^(a[50] & b[6])^(a[49] & b[7])^(a[48] & b[8])^(a[47] & b[9])^(a[46] & b[10])^(a[45] & b[11])^(a[44] & b[12])^(a[43] & b[13])^(a[42] & b[14])^(a[41] & b[15])^(a[40] & b[16])^(a[39] & b[17])^(a[38] & b[18])^(a[37] & b[19])^(a[36] & b[20])^(a[35] & b[21])^(a[34] & b[22])^(a[33] & b[23])^(a[32] & b[24])^(a[31] & b[25])^(a[30] & b[26])^(a[29] & b[27])^(a[28] & b[28])^(a[27] & b[29])^(a[26] & b[30])^(a[25] & b[31])^(a[24] & b[32])^(a[23] & b[33])^(a[22] & b[34])^(a[21] & b[35])^(a[20] & b[36])^(a[19] & b[37])^(a[18] & b[38])^(a[17] & b[39])^(a[16] & b[40])^(a[15] & b[41])^(a[14] & b[42])^(a[13] & b[43])^(a[12] & b[44])^(a[11] & b[45])^(a[10] & b[46])^(a[9] & b[47])^(a[8] & b[48])^(a[7] & b[49])^(a[6] & b[50])^(a[5] & b[51])^(a[4] & b[52])^(a[3] & b[53])^(a[2] & b[54])^(a[1] & b[55])^(a[0] & b[56]);
assign y[57] = (a[57] & b[0])^(a[56] & b[1])^(a[55] & b[2])^(a[54] & b[3])^(a[53] & b[4])^(a[52] & b[5])^(a[51] & b[6])^(a[50] & b[7])^(a[49] & b[8])^(a[48] & b[9])^(a[47] & b[10])^(a[46] & b[11])^(a[45] & b[12])^(a[44] & b[13])^(a[43] & b[14])^(a[42] & b[15])^(a[41] & b[16])^(a[40] & b[17])^(a[39] & b[18])^(a[38] & b[19])^(a[37] & b[20])^(a[36] & b[21])^(a[35] & b[22])^(a[34] & b[23])^(a[33] & b[24])^(a[32] & b[25])^(a[31] & b[26])^(a[30] & b[27])^(a[29] & b[28])^(a[28] & b[29])^(a[27] & b[30])^(a[26] & b[31])^(a[25] & b[32])^(a[24] & b[33])^(a[23] & b[34])^(a[22] & b[35])^(a[21] & b[36])^(a[20] & b[37])^(a[19] & b[38])^(a[18] & b[39])^(a[17] & b[40])^(a[16] & b[41])^(a[15] & b[42])^(a[14] & b[43])^(a[13] & b[44])^(a[12] & b[45])^(a[11] & b[46])^(a[10] & b[47])^(a[9] & b[48])^(a[8] & b[49])^(a[7] & b[50])^(a[6] & b[51])^(a[5] & b[52])^(a[4] & b[53])^(a[3] & b[54])^(a[2] & b[55])^(a[1] & b[56])^(a[0] & b[57]);
assign y[58] = (a[58] & b[0])^(a[57] & b[1])^(a[56] & b[2])^(a[55] & b[3])^(a[54] & b[4])^(a[53] & b[5])^(a[52] & b[6])^(a[51] & b[7])^(a[50] & b[8])^(a[49] & b[9])^(a[48] & b[10])^(a[47] & b[11])^(a[46] & b[12])^(a[45] & b[13])^(a[44] & b[14])^(a[43] & b[15])^(a[42] & b[16])^(a[41] & b[17])^(a[40] & b[18])^(a[39] & b[19])^(a[38] & b[20])^(a[37] & b[21])^(a[36] & b[22])^(a[35] & b[23])^(a[34] & b[24])^(a[33] & b[25])^(a[32] & b[26])^(a[31] & b[27])^(a[30] & b[28])^(a[29] & b[29])^(a[28] & b[30])^(a[27] & b[31])^(a[26] & b[32])^(a[25] & b[33])^(a[24] & b[34])^(a[23] & b[35])^(a[22] & b[36])^(a[21] & b[37])^(a[20] & b[38])^(a[19] & b[39])^(a[18] & b[40])^(a[17] & b[41])^(a[16] & b[42])^(a[15] & b[43])^(a[14] & b[44])^(a[13] & b[45])^(a[12] & b[46])^(a[11] & b[47])^(a[10] & b[48])^(a[9] & b[49])^(a[8] & b[50])^(a[7] & b[51])^(a[6] & b[52])^(a[5] & b[53])^(a[4] & b[54])^(a[3] & b[55])^(a[2] & b[56])^(a[1] & b[57])^(a[0] & b[58]);
assign y[59] = (a[59] & b[0])^(a[58] & b[1])^(a[57] & b[2])^(a[56] & b[3])^(a[55] & b[4])^(a[54] & b[5])^(a[53] & b[6])^(a[52] & b[7])^(a[51] & b[8])^(a[50] & b[9])^(a[49] & b[10])^(a[48] & b[11])^(a[47] & b[12])^(a[46] & b[13])^(a[45] & b[14])^(a[44] & b[15])^(a[43] & b[16])^(a[42] & b[17])^(a[41] & b[18])^(a[40] & b[19])^(a[39] & b[20])^(a[38] & b[21])^(a[37] & b[22])^(a[36] & b[23])^(a[35] & b[24])^(a[34] & b[25])^(a[33] & b[26])^(a[32] & b[27])^(a[31] & b[28])^(a[30] & b[29])^(a[29] & b[30])^(a[28] & b[31])^(a[27] & b[32])^(a[26] & b[33])^(a[25] & b[34])^(a[24] & b[35])^(a[23] & b[36])^(a[22] & b[37])^(a[21] & b[38])^(a[20] & b[39])^(a[19] & b[40])^(a[18] & b[41])^(a[17] & b[42])^(a[16] & b[43])^(a[15] & b[44])^(a[14] & b[45])^(a[13] & b[46])^(a[12] & b[47])^(a[11] & b[48])^(a[10] & b[49])^(a[9] & b[50])^(a[8] & b[51])^(a[7] & b[52])^(a[6] & b[53])^(a[5] & b[54])^(a[4] & b[55])^(a[3] & b[56])^(a[2] & b[57])^(a[1] & b[58])^(a[0] & b[59]);
assign y[60] = (a[60] & b[0])^(a[59] & b[1])^(a[58] & b[2])^(a[57] & b[3])^(a[56] & b[4])^(a[55] & b[5])^(a[54] & b[6])^(a[53] & b[7])^(a[52] & b[8])^(a[51] & b[9])^(a[50] & b[10])^(a[49] & b[11])^(a[48] & b[12])^(a[47] & b[13])^(a[46] & b[14])^(a[45] & b[15])^(a[44] & b[16])^(a[43] & b[17])^(a[42] & b[18])^(a[41] & b[19])^(a[40] & b[20])^(a[39] & b[21])^(a[38] & b[22])^(a[37] & b[23])^(a[36] & b[24])^(a[35] & b[25])^(a[34] & b[26])^(a[33] & b[27])^(a[32] & b[28])^(a[31] & b[29])^(a[30] & b[30])^(a[29] & b[31])^(a[28] & b[32])^(a[27] & b[33])^(a[26] & b[34])^(a[25] & b[35])^(a[24] & b[36])^(a[23] & b[37])^(a[22] & b[38])^(a[21] & b[39])^(a[20] & b[40])^(a[19] & b[41])^(a[18] & b[42])^(a[17] & b[43])^(a[16] & b[44])^(a[15] & b[45])^(a[14] & b[46])^(a[13] & b[47])^(a[12] & b[48])^(a[11] & b[49])^(a[10] & b[50])^(a[9] & b[51])^(a[8] & b[52])^(a[7] & b[53])^(a[6] & b[54])^(a[5] & b[55])^(a[4] & b[56])^(a[3] & b[57])^(a[2] & b[58])^(a[1] & b[59])^(a[0] & b[60]);
assign y[61] = (a[61] & b[0])^(a[60] & b[1])^(a[59] & b[2])^(a[58] & b[3])^(a[57] & b[4])^(a[56] & b[5])^(a[55] & b[6])^(a[54] & b[7])^(a[53] & b[8])^(a[52] & b[9])^(a[51] & b[10])^(a[50] & b[11])^(a[49] & b[12])^(a[48] & b[13])^(a[47] & b[14])^(a[46] & b[15])^(a[45] & b[16])^(a[44] & b[17])^(a[43] & b[18])^(a[42] & b[19])^(a[41] & b[20])^(a[40] & b[21])^(a[39] & b[22])^(a[38] & b[23])^(a[37] & b[24])^(a[36] & b[25])^(a[35] & b[26])^(a[34] & b[27])^(a[33] & b[28])^(a[32] & b[29])^(a[31] & b[30])^(a[30] & b[31])^(a[29] & b[32])^(a[28] & b[33])^(a[27] & b[34])^(a[26] & b[35])^(a[25] & b[36])^(a[24] & b[37])^(a[23] & b[38])^(a[22] & b[39])^(a[21] & b[40])^(a[20] & b[41])^(a[19] & b[42])^(a[18] & b[43])^(a[17] & b[44])^(a[16] & b[45])^(a[15] & b[46])^(a[14] & b[47])^(a[13] & b[48])^(a[12] & b[49])^(a[11] & b[50])^(a[10] & b[51])^(a[9] & b[52])^(a[8] & b[53])^(a[7] & b[54])^(a[6] & b[55])^(a[5] & b[56])^(a[4] & b[57])^(a[3] & b[58])^(a[2] & b[59])^(a[1] & b[60])^(a[0] & b[61]);
assign y[62] = (a[62] & b[0])^(a[61] & b[1])^(a[60] & b[2])^(a[59] & b[3])^(a[58] & b[4])^(a[57] & b[5])^(a[56] & b[6])^(a[55] & b[7])^(a[54] & b[8])^(a[53] & b[9])^(a[52] & b[10])^(a[51] & b[11])^(a[50] & b[12])^(a[49] & b[13])^(a[48] & b[14])^(a[47] & b[15])^(a[46] & b[16])^(a[45] & b[17])^(a[44] & b[18])^(a[43] & b[19])^(a[42] & b[20])^(a[41] & b[21])^(a[40] & b[22])^(a[39] & b[23])^(a[38] & b[24])^(a[37] & b[25])^(a[36] & b[26])^(a[35] & b[27])^(a[34] & b[28])^(a[33] & b[29])^(a[32] & b[30])^(a[31] & b[31])^(a[30] & b[32])^(a[29] & b[33])^(a[28] & b[34])^(a[27] & b[35])^(a[26] & b[36])^(a[25] & b[37])^(a[24] & b[38])^(a[23] & b[39])^(a[22] & b[40])^(a[21] & b[41])^(a[20] & b[42])^(a[19] & b[43])^(a[18] & b[44])^(a[17] & b[45])^(a[16] & b[46])^(a[15] & b[47])^(a[14] & b[48])^(a[13] & b[49])^(a[12] & b[50])^(a[11] & b[51])^(a[10] & b[52])^(a[9] & b[53])^(a[8] & b[54])^(a[7] & b[55])^(a[6] & b[56])^(a[5] & b[57])^(a[4] & b[58])^(a[3] & b[59])^(a[2] & b[60])^(a[1] & b[61])^(a[0] & b[62]);
assign y[63] = (a[63] & b[0])^(a[62] & b[1])^(a[61] & b[2])^(a[60] & b[3])^(a[59] & b[4])^(a[58] & b[5])^(a[57] & b[6])^(a[56] & b[7])^(a[55] & b[8])^(a[54] & b[9])^(a[53] & b[10])^(a[52] & b[11])^(a[51] & b[12])^(a[50] & b[13])^(a[49] & b[14])^(a[48] & b[15])^(a[47] & b[16])^(a[46] & b[17])^(a[45] & b[18])^(a[44] & b[19])^(a[43] & b[20])^(a[42] & b[21])^(a[41] & b[22])^(a[40] & b[23])^(a[39] & b[24])^(a[38] & b[25])^(a[37] & b[26])^(a[36] & b[27])^(a[35] & b[28])^(a[34] & b[29])^(a[33] & b[30])^(a[32] & b[31])^(a[31] & b[32])^(a[30] & b[33])^(a[29] & b[34])^(a[28] & b[35])^(a[27] & b[36])^(a[26] & b[37])^(a[25] & b[38])^(a[24] & b[39])^(a[23] & b[40])^(a[22] & b[41])^(a[21] & b[42])^(a[20] & b[43])^(a[19] & b[44])^(a[18] & b[45])^(a[17] & b[46])^(a[16] & b[47])^(a[15] & b[48])^(a[14] & b[49])^(a[13] & b[50])^(a[12] & b[51])^(a[11] & b[52])^(a[10] & b[53])^(a[9] & b[54])^(a[8] & b[55])^(a[7] & b[56])^(a[6] & b[57])^(a[5] & b[58])^(a[4] & b[59])^(a[3] & b[60])^(a[2] & b[61])^(a[1] & b[62])^(a[0] & b[63]);
assign y[64] = (a[64] & b[0])^(a[63] & b[1])^(a[62] & b[2])^(a[61] & b[3])^(a[60] & b[4])^(a[59] & b[5])^(a[58] & b[6])^(a[57] & b[7])^(a[56] & b[8])^(a[55] & b[9])^(a[54] & b[10])^(a[53] & b[11])^(a[52] & b[12])^(a[51] & b[13])^(a[50] & b[14])^(a[49] & b[15])^(a[48] & b[16])^(a[47] & b[17])^(a[46] & b[18])^(a[45] & b[19])^(a[44] & b[20])^(a[43] & b[21])^(a[42] & b[22])^(a[41] & b[23])^(a[40] & b[24])^(a[39] & b[25])^(a[38] & b[26])^(a[37] & b[27])^(a[36] & b[28])^(a[35] & b[29])^(a[34] & b[30])^(a[33] & b[31])^(a[32] & b[32])^(a[31] & b[33])^(a[30] & b[34])^(a[29] & b[35])^(a[28] & b[36])^(a[27] & b[37])^(a[26] & b[38])^(a[25] & b[39])^(a[24] & b[40])^(a[23] & b[41])^(a[22] & b[42])^(a[21] & b[43])^(a[20] & b[44])^(a[19] & b[45])^(a[18] & b[46])^(a[17] & b[47])^(a[16] & b[48])^(a[15] & b[49])^(a[14] & b[50])^(a[13] & b[51])^(a[12] & b[52])^(a[11] & b[53])^(a[10] & b[54])^(a[9] & b[55])^(a[8] & b[56])^(a[7] & b[57])^(a[6] & b[58])^(a[5] & b[59])^(a[4] & b[60])^(a[3] & b[61])^(a[2] & b[62])^(a[1] & b[63])^(a[0] & b[64]);
assign y[65] = (a[65] & b[0])^(a[64] & b[1])^(a[63] & b[2])^(a[62] & b[3])^(a[61] & b[4])^(a[60] & b[5])^(a[59] & b[6])^(a[58] & b[7])^(a[57] & b[8])^(a[56] & b[9])^(a[55] & b[10])^(a[54] & b[11])^(a[53] & b[12])^(a[52] & b[13])^(a[51] & b[14])^(a[50] & b[15])^(a[49] & b[16])^(a[48] & b[17])^(a[47] & b[18])^(a[46] & b[19])^(a[45] & b[20])^(a[44] & b[21])^(a[43] & b[22])^(a[42] & b[23])^(a[41] & b[24])^(a[40] & b[25])^(a[39] & b[26])^(a[38] & b[27])^(a[37] & b[28])^(a[36] & b[29])^(a[35] & b[30])^(a[34] & b[31])^(a[33] & b[32])^(a[32] & b[33])^(a[31] & b[34])^(a[30] & b[35])^(a[29] & b[36])^(a[28] & b[37])^(a[27] & b[38])^(a[26] & b[39])^(a[25] & b[40])^(a[24] & b[41])^(a[23] & b[42])^(a[22] & b[43])^(a[21] & b[44])^(a[20] & b[45])^(a[19] & b[46])^(a[18] & b[47])^(a[17] & b[48])^(a[16] & b[49])^(a[15] & b[50])^(a[14] & b[51])^(a[13] & b[52])^(a[12] & b[53])^(a[11] & b[54])^(a[10] & b[55])^(a[9] & b[56])^(a[8] & b[57])^(a[7] & b[58])^(a[6] & b[59])^(a[5] & b[60])^(a[4] & b[61])^(a[3] & b[62])^(a[2] & b[63])^(a[1] & b[64])^(a[0] & b[65]);
assign y[66] = (a[66] & b[0])^(a[65] & b[1])^(a[64] & b[2])^(a[63] & b[3])^(a[62] & b[4])^(a[61] & b[5])^(a[60] & b[6])^(a[59] & b[7])^(a[58] & b[8])^(a[57] & b[9])^(a[56] & b[10])^(a[55] & b[11])^(a[54] & b[12])^(a[53] & b[13])^(a[52] & b[14])^(a[51] & b[15])^(a[50] & b[16])^(a[49] & b[17])^(a[48] & b[18])^(a[47] & b[19])^(a[46] & b[20])^(a[45] & b[21])^(a[44] & b[22])^(a[43] & b[23])^(a[42] & b[24])^(a[41] & b[25])^(a[40] & b[26])^(a[39] & b[27])^(a[38] & b[28])^(a[37] & b[29])^(a[36] & b[30])^(a[35] & b[31])^(a[34] & b[32])^(a[33] & b[33])^(a[32] & b[34])^(a[31] & b[35])^(a[30] & b[36])^(a[29] & b[37])^(a[28] & b[38])^(a[27] & b[39])^(a[26] & b[40])^(a[25] & b[41])^(a[24] & b[42])^(a[23] & b[43])^(a[22] & b[44])^(a[21] & b[45])^(a[20] & b[46])^(a[19] & b[47])^(a[18] & b[48])^(a[17] & b[49])^(a[16] & b[50])^(a[15] & b[51])^(a[14] & b[52])^(a[13] & b[53])^(a[12] & b[54])^(a[11] & b[55])^(a[10] & b[56])^(a[9] & b[57])^(a[8] & b[58])^(a[7] & b[59])^(a[6] & b[60])^(a[5] & b[61])^(a[4] & b[62])^(a[3] & b[63])^(a[2] & b[64])^(a[1] & b[65])^(a[0] & b[66]);
assign y[67] = (a[67] & b[0])^(a[66] & b[1])^(a[65] & b[2])^(a[64] & b[3])^(a[63] & b[4])^(a[62] & b[5])^(a[61] & b[6])^(a[60] & b[7])^(a[59] & b[8])^(a[58] & b[9])^(a[57] & b[10])^(a[56] & b[11])^(a[55] & b[12])^(a[54] & b[13])^(a[53] & b[14])^(a[52] & b[15])^(a[51] & b[16])^(a[50] & b[17])^(a[49] & b[18])^(a[48] & b[19])^(a[47] & b[20])^(a[46] & b[21])^(a[45] & b[22])^(a[44] & b[23])^(a[43] & b[24])^(a[42] & b[25])^(a[41] & b[26])^(a[40] & b[27])^(a[39] & b[28])^(a[38] & b[29])^(a[37] & b[30])^(a[36] & b[31])^(a[35] & b[32])^(a[34] & b[33])^(a[33] & b[34])^(a[32] & b[35])^(a[31] & b[36])^(a[30] & b[37])^(a[29] & b[38])^(a[28] & b[39])^(a[27] & b[40])^(a[26] & b[41])^(a[25] & b[42])^(a[24] & b[43])^(a[23] & b[44])^(a[22] & b[45])^(a[21] & b[46])^(a[20] & b[47])^(a[19] & b[48])^(a[18] & b[49])^(a[17] & b[50])^(a[16] & b[51])^(a[15] & b[52])^(a[14] & b[53])^(a[13] & b[54])^(a[12] & b[55])^(a[11] & b[56])^(a[10] & b[57])^(a[9] & b[58])^(a[8] & b[59])^(a[7] & b[60])^(a[6] & b[61])^(a[5] & b[62])^(a[4] & b[63])^(a[3] & b[64])^(a[2] & b[65])^(a[1] & b[66])^(a[0] & b[67]);
assign y[68] = (a[68] & b[0])^(a[67] & b[1])^(a[66] & b[2])^(a[65] & b[3])^(a[64] & b[4])^(a[63] & b[5])^(a[62] & b[6])^(a[61] & b[7])^(a[60] & b[8])^(a[59] & b[9])^(a[58] & b[10])^(a[57] & b[11])^(a[56] & b[12])^(a[55] & b[13])^(a[54] & b[14])^(a[53] & b[15])^(a[52] & b[16])^(a[51] & b[17])^(a[50] & b[18])^(a[49] & b[19])^(a[48] & b[20])^(a[47] & b[21])^(a[46] & b[22])^(a[45] & b[23])^(a[44] & b[24])^(a[43] & b[25])^(a[42] & b[26])^(a[41] & b[27])^(a[40] & b[28])^(a[39] & b[29])^(a[38] & b[30])^(a[37] & b[31])^(a[36] & b[32])^(a[35] & b[33])^(a[34] & b[34])^(a[33] & b[35])^(a[32] & b[36])^(a[31] & b[37])^(a[30] & b[38])^(a[29] & b[39])^(a[28] & b[40])^(a[27] & b[41])^(a[26] & b[42])^(a[25] & b[43])^(a[24] & b[44])^(a[23] & b[45])^(a[22] & b[46])^(a[21] & b[47])^(a[20] & b[48])^(a[19] & b[49])^(a[18] & b[50])^(a[17] & b[51])^(a[16] & b[52])^(a[15] & b[53])^(a[14] & b[54])^(a[13] & b[55])^(a[12] & b[56])^(a[11] & b[57])^(a[10] & b[58])^(a[9] & b[59])^(a[8] & b[60])^(a[7] & b[61])^(a[6] & b[62])^(a[5] & b[63])^(a[4] & b[64])^(a[3] & b[65])^(a[2] & b[66])^(a[1] & b[67])^(a[0] & b[68]);
assign y[69] = (a[69] & b[0])^(a[68] & b[1])^(a[67] & b[2])^(a[66] & b[3])^(a[65] & b[4])^(a[64] & b[5])^(a[63] & b[6])^(a[62] & b[7])^(a[61] & b[8])^(a[60] & b[9])^(a[59] & b[10])^(a[58] & b[11])^(a[57] & b[12])^(a[56] & b[13])^(a[55] & b[14])^(a[54] & b[15])^(a[53] & b[16])^(a[52] & b[17])^(a[51] & b[18])^(a[50] & b[19])^(a[49] & b[20])^(a[48] & b[21])^(a[47] & b[22])^(a[46] & b[23])^(a[45] & b[24])^(a[44] & b[25])^(a[43] & b[26])^(a[42] & b[27])^(a[41] & b[28])^(a[40] & b[29])^(a[39] & b[30])^(a[38] & b[31])^(a[37] & b[32])^(a[36] & b[33])^(a[35] & b[34])^(a[34] & b[35])^(a[33] & b[36])^(a[32] & b[37])^(a[31] & b[38])^(a[30] & b[39])^(a[29] & b[40])^(a[28] & b[41])^(a[27] & b[42])^(a[26] & b[43])^(a[25] & b[44])^(a[24] & b[45])^(a[23] & b[46])^(a[22] & b[47])^(a[21] & b[48])^(a[20] & b[49])^(a[19] & b[50])^(a[18] & b[51])^(a[17] & b[52])^(a[16] & b[53])^(a[15] & b[54])^(a[14] & b[55])^(a[13] & b[56])^(a[12] & b[57])^(a[11] & b[58])^(a[10] & b[59])^(a[9] & b[60])^(a[8] & b[61])^(a[7] & b[62])^(a[6] & b[63])^(a[5] & b[64])^(a[4] & b[65])^(a[3] & b[66])^(a[2] & b[67])^(a[1] & b[68])^(a[0] & b[69]);
assign y[70] = (a[70] & b[0])^(a[69] & b[1])^(a[68] & b[2])^(a[67] & b[3])^(a[66] & b[4])^(a[65] & b[5])^(a[64] & b[6])^(a[63] & b[7])^(a[62] & b[8])^(a[61] & b[9])^(a[60] & b[10])^(a[59] & b[11])^(a[58] & b[12])^(a[57] & b[13])^(a[56] & b[14])^(a[55] & b[15])^(a[54] & b[16])^(a[53] & b[17])^(a[52] & b[18])^(a[51] & b[19])^(a[50] & b[20])^(a[49] & b[21])^(a[48] & b[22])^(a[47] & b[23])^(a[46] & b[24])^(a[45] & b[25])^(a[44] & b[26])^(a[43] & b[27])^(a[42] & b[28])^(a[41] & b[29])^(a[40] & b[30])^(a[39] & b[31])^(a[38] & b[32])^(a[37] & b[33])^(a[36] & b[34])^(a[35] & b[35])^(a[34] & b[36])^(a[33] & b[37])^(a[32] & b[38])^(a[31] & b[39])^(a[30] & b[40])^(a[29] & b[41])^(a[28] & b[42])^(a[27] & b[43])^(a[26] & b[44])^(a[25] & b[45])^(a[24] & b[46])^(a[23] & b[47])^(a[22] & b[48])^(a[21] & b[49])^(a[20] & b[50])^(a[19] & b[51])^(a[18] & b[52])^(a[17] & b[53])^(a[16] & b[54])^(a[15] & b[55])^(a[14] & b[56])^(a[13] & b[57])^(a[12] & b[58])^(a[11] & b[59])^(a[10] & b[60])^(a[9] & b[61])^(a[8] & b[62])^(a[7] & b[63])^(a[6] & b[64])^(a[5] & b[65])^(a[4] & b[66])^(a[3] & b[67])^(a[2] & b[68])^(a[1] & b[69])^(a[0] & b[70]);
assign y[71] = (a[71] & b[0])^(a[70] & b[1])^(a[69] & b[2])^(a[68] & b[3])^(a[67] & b[4])^(a[66] & b[5])^(a[65] & b[6])^(a[64] & b[7])^(a[63] & b[8])^(a[62] & b[9])^(a[61] & b[10])^(a[60] & b[11])^(a[59] & b[12])^(a[58] & b[13])^(a[57] & b[14])^(a[56] & b[15])^(a[55] & b[16])^(a[54] & b[17])^(a[53] & b[18])^(a[52] & b[19])^(a[51] & b[20])^(a[50] & b[21])^(a[49] & b[22])^(a[48] & b[23])^(a[47] & b[24])^(a[46] & b[25])^(a[45] & b[26])^(a[44] & b[27])^(a[43] & b[28])^(a[42] & b[29])^(a[41] & b[30])^(a[40] & b[31])^(a[39] & b[32])^(a[38] & b[33])^(a[37] & b[34])^(a[36] & b[35])^(a[35] & b[36])^(a[34] & b[37])^(a[33] & b[38])^(a[32] & b[39])^(a[31] & b[40])^(a[30] & b[41])^(a[29] & b[42])^(a[28] & b[43])^(a[27] & b[44])^(a[26] & b[45])^(a[25] & b[46])^(a[24] & b[47])^(a[23] & b[48])^(a[22] & b[49])^(a[21] & b[50])^(a[20] & b[51])^(a[19] & b[52])^(a[18] & b[53])^(a[17] & b[54])^(a[16] & b[55])^(a[15] & b[56])^(a[14] & b[57])^(a[13] & b[58])^(a[12] & b[59])^(a[11] & b[60])^(a[10] & b[61])^(a[9] & b[62])^(a[8] & b[63])^(a[7] & b[64])^(a[6] & b[65])^(a[5] & b[66])^(a[4] & b[67])^(a[3] & b[68])^(a[2] & b[69])^(a[1] & b[70])^(a[0] & b[71]);
assign y[72] = (a[72] & b[0])^(a[71] & b[1])^(a[70] & b[2])^(a[69] & b[3])^(a[68] & b[4])^(a[67] & b[5])^(a[66] & b[6])^(a[65] & b[7])^(a[64] & b[8])^(a[63] & b[9])^(a[62] & b[10])^(a[61] & b[11])^(a[60] & b[12])^(a[59] & b[13])^(a[58] & b[14])^(a[57] & b[15])^(a[56] & b[16])^(a[55] & b[17])^(a[54] & b[18])^(a[53] & b[19])^(a[52] & b[20])^(a[51] & b[21])^(a[50] & b[22])^(a[49] & b[23])^(a[48] & b[24])^(a[47] & b[25])^(a[46] & b[26])^(a[45] & b[27])^(a[44] & b[28])^(a[43] & b[29])^(a[42] & b[30])^(a[41] & b[31])^(a[40] & b[32])^(a[39] & b[33])^(a[38] & b[34])^(a[37] & b[35])^(a[36] & b[36])^(a[35] & b[37])^(a[34] & b[38])^(a[33] & b[39])^(a[32] & b[40])^(a[31] & b[41])^(a[30] & b[42])^(a[29] & b[43])^(a[28] & b[44])^(a[27] & b[45])^(a[26] & b[46])^(a[25] & b[47])^(a[24] & b[48])^(a[23] & b[49])^(a[22] & b[50])^(a[21] & b[51])^(a[20] & b[52])^(a[19] & b[53])^(a[18] & b[54])^(a[17] & b[55])^(a[16] & b[56])^(a[15] & b[57])^(a[14] & b[58])^(a[13] & b[59])^(a[12] & b[60])^(a[11] & b[61])^(a[10] & b[62])^(a[9] & b[63])^(a[8] & b[64])^(a[7] & b[65])^(a[6] & b[66])^(a[5] & b[67])^(a[4] & b[68])^(a[3] & b[69])^(a[2] & b[70])^(a[1] & b[71])^(a[0] & b[72]);
assign y[73] = (a[73] & b[0])^(a[72] & b[1])^(a[71] & b[2])^(a[70] & b[3])^(a[69] & b[4])^(a[68] & b[5])^(a[67] & b[6])^(a[66] & b[7])^(a[65] & b[8])^(a[64] & b[9])^(a[63] & b[10])^(a[62] & b[11])^(a[61] & b[12])^(a[60] & b[13])^(a[59] & b[14])^(a[58] & b[15])^(a[57] & b[16])^(a[56] & b[17])^(a[55] & b[18])^(a[54] & b[19])^(a[53] & b[20])^(a[52] & b[21])^(a[51] & b[22])^(a[50] & b[23])^(a[49] & b[24])^(a[48] & b[25])^(a[47] & b[26])^(a[46] & b[27])^(a[45] & b[28])^(a[44] & b[29])^(a[43] & b[30])^(a[42] & b[31])^(a[41] & b[32])^(a[40] & b[33])^(a[39] & b[34])^(a[38] & b[35])^(a[37] & b[36])^(a[36] & b[37])^(a[35] & b[38])^(a[34] & b[39])^(a[33] & b[40])^(a[32] & b[41])^(a[31] & b[42])^(a[30] & b[43])^(a[29] & b[44])^(a[28] & b[45])^(a[27] & b[46])^(a[26] & b[47])^(a[25] & b[48])^(a[24] & b[49])^(a[23] & b[50])^(a[22] & b[51])^(a[21] & b[52])^(a[20] & b[53])^(a[19] & b[54])^(a[18] & b[55])^(a[17] & b[56])^(a[16] & b[57])^(a[15] & b[58])^(a[14] & b[59])^(a[13] & b[60])^(a[12] & b[61])^(a[11] & b[62])^(a[10] & b[63])^(a[9] & b[64])^(a[8] & b[65])^(a[7] & b[66])^(a[6] & b[67])^(a[5] & b[68])^(a[4] & b[69])^(a[3] & b[70])^(a[2] & b[71])^(a[1] & b[72])^(a[0] & b[73]);
assign y[74] = (a[74] & b[0])^(a[73] & b[1])^(a[72] & b[2])^(a[71] & b[3])^(a[70] & b[4])^(a[69] & b[5])^(a[68] & b[6])^(a[67] & b[7])^(a[66] & b[8])^(a[65] & b[9])^(a[64] & b[10])^(a[63] & b[11])^(a[62] & b[12])^(a[61] & b[13])^(a[60] & b[14])^(a[59] & b[15])^(a[58] & b[16])^(a[57] & b[17])^(a[56] & b[18])^(a[55] & b[19])^(a[54] & b[20])^(a[53] & b[21])^(a[52] & b[22])^(a[51] & b[23])^(a[50] & b[24])^(a[49] & b[25])^(a[48] & b[26])^(a[47] & b[27])^(a[46] & b[28])^(a[45] & b[29])^(a[44] & b[30])^(a[43] & b[31])^(a[42] & b[32])^(a[41] & b[33])^(a[40] & b[34])^(a[39] & b[35])^(a[38] & b[36])^(a[37] & b[37])^(a[36] & b[38])^(a[35] & b[39])^(a[34] & b[40])^(a[33] & b[41])^(a[32] & b[42])^(a[31] & b[43])^(a[30] & b[44])^(a[29] & b[45])^(a[28] & b[46])^(a[27] & b[47])^(a[26] & b[48])^(a[25] & b[49])^(a[24] & b[50])^(a[23] & b[51])^(a[22] & b[52])^(a[21] & b[53])^(a[20] & b[54])^(a[19] & b[55])^(a[18] & b[56])^(a[17] & b[57])^(a[16] & b[58])^(a[15] & b[59])^(a[14] & b[60])^(a[13] & b[61])^(a[12] & b[62])^(a[11] & b[63])^(a[10] & b[64])^(a[9] & b[65])^(a[8] & b[66])^(a[7] & b[67])^(a[6] & b[68])^(a[5] & b[69])^(a[4] & b[70])^(a[3] & b[71])^(a[2] & b[72])^(a[1] & b[73])^(a[0] & b[74]);
assign y[75] = (a[75] & b[0])^(a[74] & b[1])^(a[73] & b[2])^(a[72] & b[3])^(a[71] & b[4])^(a[70] & b[5])^(a[69] & b[6])^(a[68] & b[7])^(a[67] & b[8])^(a[66] & b[9])^(a[65] & b[10])^(a[64] & b[11])^(a[63] & b[12])^(a[62] & b[13])^(a[61] & b[14])^(a[60] & b[15])^(a[59] & b[16])^(a[58] & b[17])^(a[57] & b[18])^(a[56] & b[19])^(a[55] & b[20])^(a[54] & b[21])^(a[53] & b[22])^(a[52] & b[23])^(a[51] & b[24])^(a[50] & b[25])^(a[49] & b[26])^(a[48] & b[27])^(a[47] & b[28])^(a[46] & b[29])^(a[45] & b[30])^(a[44] & b[31])^(a[43] & b[32])^(a[42] & b[33])^(a[41] & b[34])^(a[40] & b[35])^(a[39] & b[36])^(a[38] & b[37])^(a[37] & b[38])^(a[36] & b[39])^(a[35] & b[40])^(a[34] & b[41])^(a[33] & b[42])^(a[32] & b[43])^(a[31] & b[44])^(a[30] & b[45])^(a[29] & b[46])^(a[28] & b[47])^(a[27] & b[48])^(a[26] & b[49])^(a[25] & b[50])^(a[24] & b[51])^(a[23] & b[52])^(a[22] & b[53])^(a[21] & b[54])^(a[20] & b[55])^(a[19] & b[56])^(a[18] & b[57])^(a[17] & b[58])^(a[16] & b[59])^(a[15] & b[60])^(a[14] & b[61])^(a[13] & b[62])^(a[12] & b[63])^(a[11] & b[64])^(a[10] & b[65])^(a[9] & b[66])^(a[8] & b[67])^(a[7] & b[68])^(a[6] & b[69])^(a[5] & b[70])^(a[4] & b[71])^(a[3] & b[72])^(a[2] & b[73])^(a[1] & b[74])^(a[0] & b[75]);
assign y[76] = (a[76] & b[0])^(a[75] & b[1])^(a[74] & b[2])^(a[73] & b[3])^(a[72] & b[4])^(a[71] & b[5])^(a[70] & b[6])^(a[69] & b[7])^(a[68] & b[8])^(a[67] & b[9])^(a[66] & b[10])^(a[65] & b[11])^(a[64] & b[12])^(a[63] & b[13])^(a[62] & b[14])^(a[61] & b[15])^(a[60] & b[16])^(a[59] & b[17])^(a[58] & b[18])^(a[57] & b[19])^(a[56] & b[20])^(a[55] & b[21])^(a[54] & b[22])^(a[53] & b[23])^(a[52] & b[24])^(a[51] & b[25])^(a[50] & b[26])^(a[49] & b[27])^(a[48] & b[28])^(a[47] & b[29])^(a[46] & b[30])^(a[45] & b[31])^(a[44] & b[32])^(a[43] & b[33])^(a[42] & b[34])^(a[41] & b[35])^(a[40] & b[36])^(a[39] & b[37])^(a[38] & b[38])^(a[37] & b[39])^(a[36] & b[40])^(a[35] & b[41])^(a[34] & b[42])^(a[33] & b[43])^(a[32] & b[44])^(a[31] & b[45])^(a[30] & b[46])^(a[29] & b[47])^(a[28] & b[48])^(a[27] & b[49])^(a[26] & b[50])^(a[25] & b[51])^(a[24] & b[52])^(a[23] & b[53])^(a[22] & b[54])^(a[21] & b[55])^(a[20] & b[56])^(a[19] & b[57])^(a[18] & b[58])^(a[17] & b[59])^(a[16] & b[60])^(a[15] & b[61])^(a[14] & b[62])^(a[13] & b[63])^(a[12] & b[64])^(a[11] & b[65])^(a[10] & b[66])^(a[9] & b[67])^(a[8] & b[68])^(a[7] & b[69])^(a[6] & b[70])^(a[5] & b[71])^(a[4] & b[72])^(a[3] & b[73])^(a[2] & b[74])^(a[1] & b[75])^(a[0] & b[76]);
assign y[77] = (a[77] & b[0])^(a[76] & b[1])^(a[75] & b[2])^(a[74] & b[3])^(a[73] & b[4])^(a[72] & b[5])^(a[71] & b[6])^(a[70] & b[7])^(a[69] & b[8])^(a[68] & b[9])^(a[67] & b[10])^(a[66] & b[11])^(a[65] & b[12])^(a[64] & b[13])^(a[63] & b[14])^(a[62] & b[15])^(a[61] & b[16])^(a[60] & b[17])^(a[59] & b[18])^(a[58] & b[19])^(a[57] & b[20])^(a[56] & b[21])^(a[55] & b[22])^(a[54] & b[23])^(a[53] & b[24])^(a[52] & b[25])^(a[51] & b[26])^(a[50] & b[27])^(a[49] & b[28])^(a[48] & b[29])^(a[47] & b[30])^(a[46] & b[31])^(a[45] & b[32])^(a[44] & b[33])^(a[43] & b[34])^(a[42] & b[35])^(a[41] & b[36])^(a[40] & b[37])^(a[39] & b[38])^(a[38] & b[39])^(a[37] & b[40])^(a[36] & b[41])^(a[35] & b[42])^(a[34] & b[43])^(a[33] & b[44])^(a[32] & b[45])^(a[31] & b[46])^(a[30] & b[47])^(a[29] & b[48])^(a[28] & b[49])^(a[27] & b[50])^(a[26] & b[51])^(a[25] & b[52])^(a[24] & b[53])^(a[23] & b[54])^(a[22] & b[55])^(a[21] & b[56])^(a[20] & b[57])^(a[19] & b[58])^(a[18] & b[59])^(a[17] & b[60])^(a[16] & b[61])^(a[15] & b[62])^(a[14] & b[63])^(a[13] & b[64])^(a[12] & b[65])^(a[11] & b[66])^(a[10] & b[67])^(a[9] & b[68])^(a[8] & b[69])^(a[7] & b[70])^(a[6] & b[71])^(a[5] & b[72])^(a[4] & b[73])^(a[3] & b[74])^(a[2] & b[75])^(a[1] & b[76])^(a[0] & b[77]);
assign y[78] = (a[78] & b[0])^(a[77] & b[1])^(a[76] & b[2])^(a[75] & b[3])^(a[74] & b[4])^(a[73] & b[5])^(a[72] & b[6])^(a[71] & b[7])^(a[70] & b[8])^(a[69] & b[9])^(a[68] & b[10])^(a[67] & b[11])^(a[66] & b[12])^(a[65] & b[13])^(a[64] & b[14])^(a[63] & b[15])^(a[62] & b[16])^(a[61] & b[17])^(a[60] & b[18])^(a[59] & b[19])^(a[58] & b[20])^(a[57] & b[21])^(a[56] & b[22])^(a[55] & b[23])^(a[54] & b[24])^(a[53] & b[25])^(a[52] & b[26])^(a[51] & b[27])^(a[50] & b[28])^(a[49] & b[29])^(a[48] & b[30])^(a[47] & b[31])^(a[46] & b[32])^(a[45] & b[33])^(a[44] & b[34])^(a[43] & b[35])^(a[42] & b[36])^(a[41] & b[37])^(a[40] & b[38])^(a[39] & b[39])^(a[38] & b[40])^(a[37] & b[41])^(a[36] & b[42])^(a[35] & b[43])^(a[34] & b[44])^(a[33] & b[45])^(a[32] & b[46])^(a[31] & b[47])^(a[30] & b[48])^(a[29] & b[49])^(a[28] & b[50])^(a[27] & b[51])^(a[26] & b[52])^(a[25] & b[53])^(a[24] & b[54])^(a[23] & b[55])^(a[22] & b[56])^(a[21] & b[57])^(a[20] & b[58])^(a[19] & b[59])^(a[18] & b[60])^(a[17] & b[61])^(a[16] & b[62])^(a[15] & b[63])^(a[14] & b[64])^(a[13] & b[65])^(a[12] & b[66])^(a[11] & b[67])^(a[10] & b[68])^(a[9] & b[69])^(a[8] & b[70])^(a[7] & b[71])^(a[6] & b[72])^(a[5] & b[73])^(a[4] & b[74])^(a[3] & b[75])^(a[2] & b[76])^(a[1] & b[77])^(a[0] & b[78]);
assign y[79] = (a[79] & b[0])^(a[78] & b[1])^(a[77] & b[2])^(a[76] & b[3])^(a[75] & b[4])^(a[74] & b[5])^(a[73] & b[6])^(a[72] & b[7])^(a[71] & b[8])^(a[70] & b[9])^(a[69] & b[10])^(a[68] & b[11])^(a[67] & b[12])^(a[66] & b[13])^(a[65] & b[14])^(a[64] & b[15])^(a[63] & b[16])^(a[62] & b[17])^(a[61] & b[18])^(a[60] & b[19])^(a[59] & b[20])^(a[58] & b[21])^(a[57] & b[22])^(a[56] & b[23])^(a[55] & b[24])^(a[54] & b[25])^(a[53] & b[26])^(a[52] & b[27])^(a[51] & b[28])^(a[50] & b[29])^(a[49] & b[30])^(a[48] & b[31])^(a[47] & b[32])^(a[46] & b[33])^(a[45] & b[34])^(a[44] & b[35])^(a[43] & b[36])^(a[42] & b[37])^(a[41] & b[38])^(a[40] & b[39])^(a[39] & b[40])^(a[38] & b[41])^(a[37] & b[42])^(a[36] & b[43])^(a[35] & b[44])^(a[34] & b[45])^(a[33] & b[46])^(a[32] & b[47])^(a[31] & b[48])^(a[30] & b[49])^(a[29] & b[50])^(a[28] & b[51])^(a[27] & b[52])^(a[26] & b[53])^(a[25] & b[54])^(a[24] & b[55])^(a[23] & b[56])^(a[22] & b[57])^(a[21] & b[58])^(a[20] & b[59])^(a[19] & b[60])^(a[18] & b[61])^(a[17] & b[62])^(a[16] & b[63])^(a[15] & b[64])^(a[14] & b[65])^(a[13] & b[66])^(a[12] & b[67])^(a[11] & b[68])^(a[10] & b[69])^(a[9] & b[70])^(a[8] & b[71])^(a[7] & b[72])^(a[6] & b[73])^(a[5] & b[74])^(a[4] & b[75])^(a[3] & b[76])^(a[2] & b[77])^(a[1] & b[78])^(a[0] & b[79]);
assign y[80] = (a[80] & b[0])^(a[79] & b[1])^(a[78] & b[2])^(a[77] & b[3])^(a[76] & b[4])^(a[75] & b[5])^(a[74] & b[6])^(a[73] & b[7])^(a[72] & b[8])^(a[71] & b[9])^(a[70] & b[10])^(a[69] & b[11])^(a[68] & b[12])^(a[67] & b[13])^(a[66] & b[14])^(a[65] & b[15])^(a[64] & b[16])^(a[63] & b[17])^(a[62] & b[18])^(a[61] & b[19])^(a[60] & b[20])^(a[59] & b[21])^(a[58] & b[22])^(a[57] & b[23])^(a[56] & b[24])^(a[55] & b[25])^(a[54] & b[26])^(a[53] & b[27])^(a[52] & b[28])^(a[51] & b[29])^(a[50] & b[30])^(a[49] & b[31])^(a[48] & b[32])^(a[47] & b[33])^(a[46] & b[34])^(a[45] & b[35])^(a[44] & b[36])^(a[43] & b[37])^(a[42] & b[38])^(a[41] & b[39])^(a[40] & b[40])^(a[39] & b[41])^(a[38] & b[42])^(a[37] & b[43])^(a[36] & b[44])^(a[35] & b[45])^(a[34] & b[46])^(a[33] & b[47])^(a[32] & b[48])^(a[31] & b[49])^(a[30] & b[50])^(a[29] & b[51])^(a[28] & b[52])^(a[27] & b[53])^(a[26] & b[54])^(a[25] & b[55])^(a[24] & b[56])^(a[23] & b[57])^(a[22] & b[58])^(a[21] & b[59])^(a[20] & b[60])^(a[19] & b[61])^(a[18] & b[62])^(a[17] & b[63])^(a[16] & b[64])^(a[15] & b[65])^(a[14] & b[66])^(a[13] & b[67])^(a[12] & b[68])^(a[11] & b[69])^(a[10] & b[70])^(a[9] & b[71])^(a[8] & b[72])^(a[7] & b[73])^(a[6] & b[74])^(a[5] & b[75])^(a[4] & b[76])^(a[3] & b[77])^(a[2] & b[78])^(a[1] & b[79])^(a[0] & b[80]);
assign y[81] = (a[81] & b[0])^(a[80] & b[1])^(a[79] & b[2])^(a[78] & b[3])^(a[77] & b[4])^(a[76] & b[5])^(a[75] & b[6])^(a[74] & b[7])^(a[73] & b[8])^(a[72] & b[9])^(a[71] & b[10])^(a[70] & b[11])^(a[69] & b[12])^(a[68] & b[13])^(a[67] & b[14])^(a[66] & b[15])^(a[65] & b[16])^(a[64] & b[17])^(a[63] & b[18])^(a[62] & b[19])^(a[61] & b[20])^(a[60] & b[21])^(a[59] & b[22])^(a[58] & b[23])^(a[57] & b[24])^(a[56] & b[25])^(a[55] & b[26])^(a[54] & b[27])^(a[53] & b[28])^(a[52] & b[29])^(a[51] & b[30])^(a[50] & b[31])^(a[49] & b[32])^(a[48] & b[33])^(a[47] & b[34])^(a[46] & b[35])^(a[45] & b[36])^(a[44] & b[37])^(a[43] & b[38])^(a[42] & b[39])^(a[41] & b[40])^(a[40] & b[41])^(a[39] & b[42])^(a[38] & b[43])^(a[37] & b[44])^(a[36] & b[45])^(a[35] & b[46])^(a[34] & b[47])^(a[33] & b[48])^(a[32] & b[49])^(a[31] & b[50])^(a[30] & b[51])^(a[29] & b[52])^(a[28] & b[53])^(a[27] & b[54])^(a[26] & b[55])^(a[25] & b[56])^(a[24] & b[57])^(a[23] & b[58])^(a[22] & b[59])^(a[21] & b[60])^(a[20] & b[61])^(a[19] & b[62])^(a[18] & b[63])^(a[17] & b[64])^(a[16] & b[65])^(a[15] & b[66])^(a[14] & b[67])^(a[13] & b[68])^(a[12] & b[69])^(a[11] & b[70])^(a[10] & b[71])^(a[9] & b[72])^(a[8] & b[73])^(a[7] & b[74])^(a[6] & b[75])^(a[5] & b[76])^(a[4] & b[77])^(a[3] & b[78])^(a[2] & b[79])^(a[1] & b[80])^(a[0] & b[81]);
assign y[82] = (a[82] & b[0])^(a[81] & b[1])^(a[80] & b[2])^(a[79] & b[3])^(a[78] & b[4])^(a[77] & b[5])^(a[76] & b[6])^(a[75] & b[7])^(a[74] & b[8])^(a[73] & b[9])^(a[72] & b[10])^(a[71] & b[11])^(a[70] & b[12])^(a[69] & b[13])^(a[68] & b[14])^(a[67] & b[15])^(a[66] & b[16])^(a[65] & b[17])^(a[64] & b[18])^(a[63] & b[19])^(a[62] & b[20])^(a[61] & b[21])^(a[60] & b[22])^(a[59] & b[23])^(a[58] & b[24])^(a[57] & b[25])^(a[56] & b[26])^(a[55] & b[27])^(a[54] & b[28])^(a[53] & b[29])^(a[52] & b[30])^(a[51] & b[31])^(a[50] & b[32])^(a[49] & b[33])^(a[48] & b[34])^(a[47] & b[35])^(a[46] & b[36])^(a[45] & b[37])^(a[44] & b[38])^(a[43] & b[39])^(a[42] & b[40])^(a[41] & b[41])^(a[40] & b[42])^(a[39] & b[43])^(a[38] & b[44])^(a[37] & b[45])^(a[36] & b[46])^(a[35] & b[47])^(a[34] & b[48])^(a[33] & b[49])^(a[32] & b[50])^(a[31] & b[51])^(a[30] & b[52])^(a[29] & b[53])^(a[28] & b[54])^(a[27] & b[55])^(a[26] & b[56])^(a[25] & b[57])^(a[24] & b[58])^(a[23] & b[59])^(a[22] & b[60])^(a[21] & b[61])^(a[20] & b[62])^(a[19] & b[63])^(a[18] & b[64])^(a[17] & b[65])^(a[16] & b[66])^(a[15] & b[67])^(a[14] & b[68])^(a[13] & b[69])^(a[12] & b[70])^(a[11] & b[71])^(a[10] & b[72])^(a[9] & b[73])^(a[8] & b[74])^(a[7] & b[75])^(a[6] & b[76])^(a[5] & b[77])^(a[4] & b[78])^(a[3] & b[79])^(a[2] & b[80])^(a[1] & b[81])^(a[0] & b[82]);
assign y[83] = (a[83] & b[0])^(a[82] & b[1])^(a[81] & b[2])^(a[80] & b[3])^(a[79] & b[4])^(a[78] & b[5])^(a[77] & b[6])^(a[76] & b[7])^(a[75] & b[8])^(a[74] & b[9])^(a[73] & b[10])^(a[72] & b[11])^(a[71] & b[12])^(a[70] & b[13])^(a[69] & b[14])^(a[68] & b[15])^(a[67] & b[16])^(a[66] & b[17])^(a[65] & b[18])^(a[64] & b[19])^(a[63] & b[20])^(a[62] & b[21])^(a[61] & b[22])^(a[60] & b[23])^(a[59] & b[24])^(a[58] & b[25])^(a[57] & b[26])^(a[56] & b[27])^(a[55] & b[28])^(a[54] & b[29])^(a[53] & b[30])^(a[52] & b[31])^(a[51] & b[32])^(a[50] & b[33])^(a[49] & b[34])^(a[48] & b[35])^(a[47] & b[36])^(a[46] & b[37])^(a[45] & b[38])^(a[44] & b[39])^(a[43] & b[40])^(a[42] & b[41])^(a[41] & b[42])^(a[40] & b[43])^(a[39] & b[44])^(a[38] & b[45])^(a[37] & b[46])^(a[36] & b[47])^(a[35] & b[48])^(a[34] & b[49])^(a[33] & b[50])^(a[32] & b[51])^(a[31] & b[52])^(a[30] & b[53])^(a[29] & b[54])^(a[28] & b[55])^(a[27] & b[56])^(a[26] & b[57])^(a[25] & b[58])^(a[24] & b[59])^(a[23] & b[60])^(a[22] & b[61])^(a[21] & b[62])^(a[20] & b[63])^(a[19] & b[64])^(a[18] & b[65])^(a[17] & b[66])^(a[16] & b[67])^(a[15] & b[68])^(a[14] & b[69])^(a[13] & b[70])^(a[12] & b[71])^(a[11] & b[72])^(a[10] & b[73])^(a[9] & b[74])^(a[8] & b[75])^(a[7] & b[76])^(a[6] & b[77])^(a[5] & b[78])^(a[4] & b[79])^(a[3] & b[80])^(a[2] & b[81])^(a[1] & b[82])^(a[0] & b[83]);
assign y[84] = (a[84] & b[0])^(a[83] & b[1])^(a[82] & b[2])^(a[81] & b[3])^(a[80] & b[4])^(a[79] & b[5])^(a[78] & b[6])^(a[77] & b[7])^(a[76] & b[8])^(a[75] & b[9])^(a[74] & b[10])^(a[73] & b[11])^(a[72] & b[12])^(a[71] & b[13])^(a[70] & b[14])^(a[69] & b[15])^(a[68] & b[16])^(a[67] & b[17])^(a[66] & b[18])^(a[65] & b[19])^(a[64] & b[20])^(a[63] & b[21])^(a[62] & b[22])^(a[61] & b[23])^(a[60] & b[24])^(a[59] & b[25])^(a[58] & b[26])^(a[57] & b[27])^(a[56] & b[28])^(a[55] & b[29])^(a[54] & b[30])^(a[53] & b[31])^(a[52] & b[32])^(a[51] & b[33])^(a[50] & b[34])^(a[49] & b[35])^(a[48] & b[36])^(a[47] & b[37])^(a[46] & b[38])^(a[45] & b[39])^(a[44] & b[40])^(a[43] & b[41])^(a[42] & b[42])^(a[41] & b[43])^(a[40] & b[44])^(a[39] & b[45])^(a[38] & b[46])^(a[37] & b[47])^(a[36] & b[48])^(a[35] & b[49])^(a[34] & b[50])^(a[33] & b[51])^(a[32] & b[52])^(a[31] & b[53])^(a[30] & b[54])^(a[29] & b[55])^(a[28] & b[56])^(a[27] & b[57])^(a[26] & b[58])^(a[25] & b[59])^(a[24] & b[60])^(a[23] & b[61])^(a[22] & b[62])^(a[21] & b[63])^(a[20] & b[64])^(a[19] & b[65])^(a[18] & b[66])^(a[17] & b[67])^(a[16] & b[68])^(a[15] & b[69])^(a[14] & b[70])^(a[13] & b[71])^(a[12] & b[72])^(a[11] & b[73])^(a[10] & b[74])^(a[9] & b[75])^(a[8] & b[76])^(a[7] & b[77])^(a[6] & b[78])^(a[5] & b[79])^(a[4] & b[80])^(a[3] & b[81])^(a[2] & b[82])^(a[1] & b[83])^(a[0] & b[84]);
assign y[85] = (a[85] & b[0])^(a[84] & b[1])^(a[83] & b[2])^(a[82] & b[3])^(a[81] & b[4])^(a[80] & b[5])^(a[79] & b[6])^(a[78] & b[7])^(a[77] & b[8])^(a[76] & b[9])^(a[75] & b[10])^(a[74] & b[11])^(a[73] & b[12])^(a[72] & b[13])^(a[71] & b[14])^(a[70] & b[15])^(a[69] & b[16])^(a[68] & b[17])^(a[67] & b[18])^(a[66] & b[19])^(a[65] & b[20])^(a[64] & b[21])^(a[63] & b[22])^(a[62] & b[23])^(a[61] & b[24])^(a[60] & b[25])^(a[59] & b[26])^(a[58] & b[27])^(a[57] & b[28])^(a[56] & b[29])^(a[55] & b[30])^(a[54] & b[31])^(a[53] & b[32])^(a[52] & b[33])^(a[51] & b[34])^(a[50] & b[35])^(a[49] & b[36])^(a[48] & b[37])^(a[47] & b[38])^(a[46] & b[39])^(a[45] & b[40])^(a[44] & b[41])^(a[43] & b[42])^(a[42] & b[43])^(a[41] & b[44])^(a[40] & b[45])^(a[39] & b[46])^(a[38] & b[47])^(a[37] & b[48])^(a[36] & b[49])^(a[35] & b[50])^(a[34] & b[51])^(a[33] & b[52])^(a[32] & b[53])^(a[31] & b[54])^(a[30] & b[55])^(a[29] & b[56])^(a[28] & b[57])^(a[27] & b[58])^(a[26] & b[59])^(a[25] & b[60])^(a[24] & b[61])^(a[23] & b[62])^(a[22] & b[63])^(a[21] & b[64])^(a[20] & b[65])^(a[19] & b[66])^(a[18] & b[67])^(a[17] & b[68])^(a[16] & b[69])^(a[15] & b[70])^(a[14] & b[71])^(a[13] & b[72])^(a[12] & b[73])^(a[11] & b[74])^(a[10] & b[75])^(a[9] & b[76])^(a[8] & b[77])^(a[7] & b[78])^(a[6] & b[79])^(a[5] & b[80])^(a[4] & b[81])^(a[3] & b[82])^(a[2] & b[83])^(a[1] & b[84])^(a[0] & b[85]);
assign y[86] = (a[86] & b[0])^(a[85] & b[1])^(a[84] & b[2])^(a[83] & b[3])^(a[82] & b[4])^(a[81] & b[5])^(a[80] & b[6])^(a[79] & b[7])^(a[78] & b[8])^(a[77] & b[9])^(a[76] & b[10])^(a[75] & b[11])^(a[74] & b[12])^(a[73] & b[13])^(a[72] & b[14])^(a[71] & b[15])^(a[70] & b[16])^(a[69] & b[17])^(a[68] & b[18])^(a[67] & b[19])^(a[66] & b[20])^(a[65] & b[21])^(a[64] & b[22])^(a[63] & b[23])^(a[62] & b[24])^(a[61] & b[25])^(a[60] & b[26])^(a[59] & b[27])^(a[58] & b[28])^(a[57] & b[29])^(a[56] & b[30])^(a[55] & b[31])^(a[54] & b[32])^(a[53] & b[33])^(a[52] & b[34])^(a[51] & b[35])^(a[50] & b[36])^(a[49] & b[37])^(a[48] & b[38])^(a[47] & b[39])^(a[46] & b[40])^(a[45] & b[41])^(a[44] & b[42])^(a[43] & b[43])^(a[42] & b[44])^(a[41] & b[45])^(a[40] & b[46])^(a[39] & b[47])^(a[38] & b[48])^(a[37] & b[49])^(a[36] & b[50])^(a[35] & b[51])^(a[34] & b[52])^(a[33] & b[53])^(a[32] & b[54])^(a[31] & b[55])^(a[30] & b[56])^(a[29] & b[57])^(a[28] & b[58])^(a[27] & b[59])^(a[26] & b[60])^(a[25] & b[61])^(a[24] & b[62])^(a[23] & b[63])^(a[22] & b[64])^(a[21] & b[65])^(a[20] & b[66])^(a[19] & b[67])^(a[18] & b[68])^(a[17] & b[69])^(a[16] & b[70])^(a[15] & b[71])^(a[14] & b[72])^(a[13] & b[73])^(a[12] & b[74])^(a[11] & b[75])^(a[10] & b[76])^(a[9] & b[77])^(a[8] & b[78])^(a[7] & b[79])^(a[6] & b[80])^(a[5] & b[81])^(a[4] & b[82])^(a[3] & b[83])^(a[2] & b[84])^(a[1] & b[85])^(a[0] & b[86]);
assign y[87] = (a[87] & b[0])^(a[86] & b[1])^(a[85] & b[2])^(a[84] & b[3])^(a[83] & b[4])^(a[82] & b[5])^(a[81] & b[6])^(a[80] & b[7])^(a[79] & b[8])^(a[78] & b[9])^(a[77] & b[10])^(a[76] & b[11])^(a[75] & b[12])^(a[74] & b[13])^(a[73] & b[14])^(a[72] & b[15])^(a[71] & b[16])^(a[70] & b[17])^(a[69] & b[18])^(a[68] & b[19])^(a[67] & b[20])^(a[66] & b[21])^(a[65] & b[22])^(a[64] & b[23])^(a[63] & b[24])^(a[62] & b[25])^(a[61] & b[26])^(a[60] & b[27])^(a[59] & b[28])^(a[58] & b[29])^(a[57] & b[30])^(a[56] & b[31])^(a[55] & b[32])^(a[54] & b[33])^(a[53] & b[34])^(a[52] & b[35])^(a[51] & b[36])^(a[50] & b[37])^(a[49] & b[38])^(a[48] & b[39])^(a[47] & b[40])^(a[46] & b[41])^(a[45] & b[42])^(a[44] & b[43])^(a[43] & b[44])^(a[42] & b[45])^(a[41] & b[46])^(a[40] & b[47])^(a[39] & b[48])^(a[38] & b[49])^(a[37] & b[50])^(a[36] & b[51])^(a[35] & b[52])^(a[34] & b[53])^(a[33] & b[54])^(a[32] & b[55])^(a[31] & b[56])^(a[30] & b[57])^(a[29] & b[58])^(a[28] & b[59])^(a[27] & b[60])^(a[26] & b[61])^(a[25] & b[62])^(a[24] & b[63])^(a[23] & b[64])^(a[22] & b[65])^(a[21] & b[66])^(a[20] & b[67])^(a[19] & b[68])^(a[18] & b[69])^(a[17] & b[70])^(a[16] & b[71])^(a[15] & b[72])^(a[14] & b[73])^(a[13] & b[74])^(a[12] & b[75])^(a[11] & b[76])^(a[10] & b[77])^(a[9] & b[78])^(a[8] & b[79])^(a[7] & b[80])^(a[6] & b[81])^(a[5] & b[82])^(a[4] & b[83])^(a[3] & b[84])^(a[2] & b[85])^(a[1] & b[86])^(a[0] & b[87]);
assign y[88] = (a[88] & b[0])^(a[87] & b[1])^(a[86] & b[2])^(a[85] & b[3])^(a[84] & b[4])^(a[83] & b[5])^(a[82] & b[6])^(a[81] & b[7])^(a[80] & b[8])^(a[79] & b[9])^(a[78] & b[10])^(a[77] & b[11])^(a[76] & b[12])^(a[75] & b[13])^(a[74] & b[14])^(a[73] & b[15])^(a[72] & b[16])^(a[71] & b[17])^(a[70] & b[18])^(a[69] & b[19])^(a[68] & b[20])^(a[67] & b[21])^(a[66] & b[22])^(a[65] & b[23])^(a[64] & b[24])^(a[63] & b[25])^(a[62] & b[26])^(a[61] & b[27])^(a[60] & b[28])^(a[59] & b[29])^(a[58] & b[30])^(a[57] & b[31])^(a[56] & b[32])^(a[55] & b[33])^(a[54] & b[34])^(a[53] & b[35])^(a[52] & b[36])^(a[51] & b[37])^(a[50] & b[38])^(a[49] & b[39])^(a[48] & b[40])^(a[47] & b[41])^(a[46] & b[42])^(a[45] & b[43])^(a[44] & b[44])^(a[43] & b[45])^(a[42] & b[46])^(a[41] & b[47])^(a[40] & b[48])^(a[39] & b[49])^(a[38] & b[50])^(a[37] & b[51])^(a[36] & b[52])^(a[35] & b[53])^(a[34] & b[54])^(a[33] & b[55])^(a[32] & b[56])^(a[31] & b[57])^(a[30] & b[58])^(a[29] & b[59])^(a[28] & b[60])^(a[27] & b[61])^(a[26] & b[62])^(a[25] & b[63])^(a[24] & b[64])^(a[23] & b[65])^(a[22] & b[66])^(a[21] & b[67])^(a[20] & b[68])^(a[19] & b[69])^(a[18] & b[70])^(a[17] & b[71])^(a[16] & b[72])^(a[15] & b[73])^(a[14] & b[74])^(a[13] & b[75])^(a[12] & b[76])^(a[11] & b[77])^(a[10] & b[78])^(a[9] & b[79])^(a[8] & b[80])^(a[7] & b[81])^(a[6] & b[82])^(a[5] & b[83])^(a[4] & b[84])^(a[3] & b[85])^(a[2] & b[86])^(a[1] & b[87])^(a[0] & b[88]);
assign y[89] = (a[89] & b[0])^(a[88] & b[1])^(a[87] & b[2])^(a[86] & b[3])^(a[85] & b[4])^(a[84] & b[5])^(a[83] & b[6])^(a[82] & b[7])^(a[81] & b[8])^(a[80] & b[9])^(a[79] & b[10])^(a[78] & b[11])^(a[77] & b[12])^(a[76] & b[13])^(a[75] & b[14])^(a[74] & b[15])^(a[73] & b[16])^(a[72] & b[17])^(a[71] & b[18])^(a[70] & b[19])^(a[69] & b[20])^(a[68] & b[21])^(a[67] & b[22])^(a[66] & b[23])^(a[65] & b[24])^(a[64] & b[25])^(a[63] & b[26])^(a[62] & b[27])^(a[61] & b[28])^(a[60] & b[29])^(a[59] & b[30])^(a[58] & b[31])^(a[57] & b[32])^(a[56] & b[33])^(a[55] & b[34])^(a[54] & b[35])^(a[53] & b[36])^(a[52] & b[37])^(a[51] & b[38])^(a[50] & b[39])^(a[49] & b[40])^(a[48] & b[41])^(a[47] & b[42])^(a[46] & b[43])^(a[45] & b[44])^(a[44] & b[45])^(a[43] & b[46])^(a[42] & b[47])^(a[41] & b[48])^(a[40] & b[49])^(a[39] & b[50])^(a[38] & b[51])^(a[37] & b[52])^(a[36] & b[53])^(a[35] & b[54])^(a[34] & b[55])^(a[33] & b[56])^(a[32] & b[57])^(a[31] & b[58])^(a[30] & b[59])^(a[29] & b[60])^(a[28] & b[61])^(a[27] & b[62])^(a[26] & b[63])^(a[25] & b[64])^(a[24] & b[65])^(a[23] & b[66])^(a[22] & b[67])^(a[21] & b[68])^(a[20] & b[69])^(a[19] & b[70])^(a[18] & b[71])^(a[17] & b[72])^(a[16] & b[73])^(a[15] & b[74])^(a[14] & b[75])^(a[13] & b[76])^(a[12] & b[77])^(a[11] & b[78])^(a[10] & b[79])^(a[9] & b[80])^(a[8] & b[81])^(a[7] & b[82])^(a[6] & b[83])^(a[5] & b[84])^(a[4] & b[85])^(a[3] & b[86])^(a[2] & b[87])^(a[1] & b[88])^(a[0] & b[89]);
assign y[90] = (a[90] & b[0])^(a[89] & b[1])^(a[88] & b[2])^(a[87] & b[3])^(a[86] & b[4])^(a[85] & b[5])^(a[84] & b[6])^(a[83] & b[7])^(a[82] & b[8])^(a[81] & b[9])^(a[80] & b[10])^(a[79] & b[11])^(a[78] & b[12])^(a[77] & b[13])^(a[76] & b[14])^(a[75] & b[15])^(a[74] & b[16])^(a[73] & b[17])^(a[72] & b[18])^(a[71] & b[19])^(a[70] & b[20])^(a[69] & b[21])^(a[68] & b[22])^(a[67] & b[23])^(a[66] & b[24])^(a[65] & b[25])^(a[64] & b[26])^(a[63] & b[27])^(a[62] & b[28])^(a[61] & b[29])^(a[60] & b[30])^(a[59] & b[31])^(a[58] & b[32])^(a[57] & b[33])^(a[56] & b[34])^(a[55] & b[35])^(a[54] & b[36])^(a[53] & b[37])^(a[52] & b[38])^(a[51] & b[39])^(a[50] & b[40])^(a[49] & b[41])^(a[48] & b[42])^(a[47] & b[43])^(a[46] & b[44])^(a[45] & b[45])^(a[44] & b[46])^(a[43] & b[47])^(a[42] & b[48])^(a[41] & b[49])^(a[40] & b[50])^(a[39] & b[51])^(a[38] & b[52])^(a[37] & b[53])^(a[36] & b[54])^(a[35] & b[55])^(a[34] & b[56])^(a[33] & b[57])^(a[32] & b[58])^(a[31] & b[59])^(a[30] & b[60])^(a[29] & b[61])^(a[28] & b[62])^(a[27] & b[63])^(a[26] & b[64])^(a[25] & b[65])^(a[24] & b[66])^(a[23] & b[67])^(a[22] & b[68])^(a[21] & b[69])^(a[20] & b[70])^(a[19] & b[71])^(a[18] & b[72])^(a[17] & b[73])^(a[16] & b[74])^(a[15] & b[75])^(a[14] & b[76])^(a[13] & b[77])^(a[12] & b[78])^(a[11] & b[79])^(a[10] & b[80])^(a[9] & b[81])^(a[8] & b[82])^(a[7] & b[83])^(a[6] & b[84])^(a[5] & b[85])^(a[4] & b[86])^(a[3] & b[87])^(a[2] & b[88])^(a[1] & b[89])^(a[0] & b[90]);
assign y[91] = (a[91] & b[0])^(a[90] & b[1])^(a[89] & b[2])^(a[88] & b[3])^(a[87] & b[4])^(a[86] & b[5])^(a[85] & b[6])^(a[84] & b[7])^(a[83] & b[8])^(a[82] & b[9])^(a[81] & b[10])^(a[80] & b[11])^(a[79] & b[12])^(a[78] & b[13])^(a[77] & b[14])^(a[76] & b[15])^(a[75] & b[16])^(a[74] & b[17])^(a[73] & b[18])^(a[72] & b[19])^(a[71] & b[20])^(a[70] & b[21])^(a[69] & b[22])^(a[68] & b[23])^(a[67] & b[24])^(a[66] & b[25])^(a[65] & b[26])^(a[64] & b[27])^(a[63] & b[28])^(a[62] & b[29])^(a[61] & b[30])^(a[60] & b[31])^(a[59] & b[32])^(a[58] & b[33])^(a[57] & b[34])^(a[56] & b[35])^(a[55] & b[36])^(a[54] & b[37])^(a[53] & b[38])^(a[52] & b[39])^(a[51] & b[40])^(a[50] & b[41])^(a[49] & b[42])^(a[48] & b[43])^(a[47] & b[44])^(a[46] & b[45])^(a[45] & b[46])^(a[44] & b[47])^(a[43] & b[48])^(a[42] & b[49])^(a[41] & b[50])^(a[40] & b[51])^(a[39] & b[52])^(a[38] & b[53])^(a[37] & b[54])^(a[36] & b[55])^(a[35] & b[56])^(a[34] & b[57])^(a[33] & b[58])^(a[32] & b[59])^(a[31] & b[60])^(a[30] & b[61])^(a[29] & b[62])^(a[28] & b[63])^(a[27] & b[64])^(a[26] & b[65])^(a[25] & b[66])^(a[24] & b[67])^(a[23] & b[68])^(a[22] & b[69])^(a[21] & b[70])^(a[20] & b[71])^(a[19] & b[72])^(a[18] & b[73])^(a[17] & b[74])^(a[16] & b[75])^(a[15] & b[76])^(a[14] & b[77])^(a[13] & b[78])^(a[12] & b[79])^(a[11] & b[80])^(a[10] & b[81])^(a[9] & b[82])^(a[8] & b[83])^(a[7] & b[84])^(a[6] & b[85])^(a[5] & b[86])^(a[4] & b[87])^(a[3] & b[88])^(a[2] & b[89])^(a[1] & b[90])^(a[0] & b[91]);
assign y[92] = (a[92] & b[0])^(a[91] & b[1])^(a[90] & b[2])^(a[89] & b[3])^(a[88] & b[4])^(a[87] & b[5])^(a[86] & b[6])^(a[85] & b[7])^(a[84] & b[8])^(a[83] & b[9])^(a[82] & b[10])^(a[81] & b[11])^(a[80] & b[12])^(a[79] & b[13])^(a[78] & b[14])^(a[77] & b[15])^(a[76] & b[16])^(a[75] & b[17])^(a[74] & b[18])^(a[73] & b[19])^(a[72] & b[20])^(a[71] & b[21])^(a[70] & b[22])^(a[69] & b[23])^(a[68] & b[24])^(a[67] & b[25])^(a[66] & b[26])^(a[65] & b[27])^(a[64] & b[28])^(a[63] & b[29])^(a[62] & b[30])^(a[61] & b[31])^(a[60] & b[32])^(a[59] & b[33])^(a[58] & b[34])^(a[57] & b[35])^(a[56] & b[36])^(a[55] & b[37])^(a[54] & b[38])^(a[53] & b[39])^(a[52] & b[40])^(a[51] & b[41])^(a[50] & b[42])^(a[49] & b[43])^(a[48] & b[44])^(a[47] & b[45])^(a[46] & b[46])^(a[45] & b[47])^(a[44] & b[48])^(a[43] & b[49])^(a[42] & b[50])^(a[41] & b[51])^(a[40] & b[52])^(a[39] & b[53])^(a[38] & b[54])^(a[37] & b[55])^(a[36] & b[56])^(a[35] & b[57])^(a[34] & b[58])^(a[33] & b[59])^(a[32] & b[60])^(a[31] & b[61])^(a[30] & b[62])^(a[29] & b[63])^(a[28] & b[64])^(a[27] & b[65])^(a[26] & b[66])^(a[25] & b[67])^(a[24] & b[68])^(a[23] & b[69])^(a[22] & b[70])^(a[21] & b[71])^(a[20] & b[72])^(a[19] & b[73])^(a[18] & b[74])^(a[17] & b[75])^(a[16] & b[76])^(a[15] & b[77])^(a[14] & b[78])^(a[13] & b[79])^(a[12] & b[80])^(a[11] & b[81])^(a[10] & b[82])^(a[9] & b[83])^(a[8] & b[84])^(a[7] & b[85])^(a[6] & b[86])^(a[5] & b[87])^(a[4] & b[88])^(a[3] & b[89])^(a[2] & b[90])^(a[1] & b[91])^(a[0] & b[92]);
assign y[93] = (a[93] & b[0])^(a[92] & b[1])^(a[91] & b[2])^(a[90] & b[3])^(a[89] & b[4])^(a[88] & b[5])^(a[87] & b[6])^(a[86] & b[7])^(a[85] & b[8])^(a[84] & b[9])^(a[83] & b[10])^(a[82] & b[11])^(a[81] & b[12])^(a[80] & b[13])^(a[79] & b[14])^(a[78] & b[15])^(a[77] & b[16])^(a[76] & b[17])^(a[75] & b[18])^(a[74] & b[19])^(a[73] & b[20])^(a[72] & b[21])^(a[71] & b[22])^(a[70] & b[23])^(a[69] & b[24])^(a[68] & b[25])^(a[67] & b[26])^(a[66] & b[27])^(a[65] & b[28])^(a[64] & b[29])^(a[63] & b[30])^(a[62] & b[31])^(a[61] & b[32])^(a[60] & b[33])^(a[59] & b[34])^(a[58] & b[35])^(a[57] & b[36])^(a[56] & b[37])^(a[55] & b[38])^(a[54] & b[39])^(a[53] & b[40])^(a[52] & b[41])^(a[51] & b[42])^(a[50] & b[43])^(a[49] & b[44])^(a[48] & b[45])^(a[47] & b[46])^(a[46] & b[47])^(a[45] & b[48])^(a[44] & b[49])^(a[43] & b[50])^(a[42] & b[51])^(a[41] & b[52])^(a[40] & b[53])^(a[39] & b[54])^(a[38] & b[55])^(a[37] & b[56])^(a[36] & b[57])^(a[35] & b[58])^(a[34] & b[59])^(a[33] & b[60])^(a[32] & b[61])^(a[31] & b[62])^(a[30] & b[63])^(a[29] & b[64])^(a[28] & b[65])^(a[27] & b[66])^(a[26] & b[67])^(a[25] & b[68])^(a[24] & b[69])^(a[23] & b[70])^(a[22] & b[71])^(a[21] & b[72])^(a[20] & b[73])^(a[19] & b[74])^(a[18] & b[75])^(a[17] & b[76])^(a[16] & b[77])^(a[15] & b[78])^(a[14] & b[79])^(a[13] & b[80])^(a[12] & b[81])^(a[11] & b[82])^(a[10] & b[83])^(a[9] & b[84])^(a[8] & b[85])^(a[7] & b[86])^(a[6] & b[87])^(a[5] & b[88])^(a[4] & b[89])^(a[3] & b[90])^(a[2] & b[91])^(a[1] & b[92])^(a[0] & b[93]);
assign y[94] = (a[94] & b[0])^(a[93] & b[1])^(a[92] & b[2])^(a[91] & b[3])^(a[90] & b[4])^(a[89] & b[5])^(a[88] & b[6])^(a[87] & b[7])^(a[86] & b[8])^(a[85] & b[9])^(a[84] & b[10])^(a[83] & b[11])^(a[82] & b[12])^(a[81] & b[13])^(a[80] & b[14])^(a[79] & b[15])^(a[78] & b[16])^(a[77] & b[17])^(a[76] & b[18])^(a[75] & b[19])^(a[74] & b[20])^(a[73] & b[21])^(a[72] & b[22])^(a[71] & b[23])^(a[70] & b[24])^(a[69] & b[25])^(a[68] & b[26])^(a[67] & b[27])^(a[66] & b[28])^(a[65] & b[29])^(a[64] & b[30])^(a[63] & b[31])^(a[62] & b[32])^(a[61] & b[33])^(a[60] & b[34])^(a[59] & b[35])^(a[58] & b[36])^(a[57] & b[37])^(a[56] & b[38])^(a[55] & b[39])^(a[54] & b[40])^(a[53] & b[41])^(a[52] & b[42])^(a[51] & b[43])^(a[50] & b[44])^(a[49] & b[45])^(a[48] & b[46])^(a[47] & b[47])^(a[46] & b[48])^(a[45] & b[49])^(a[44] & b[50])^(a[43] & b[51])^(a[42] & b[52])^(a[41] & b[53])^(a[40] & b[54])^(a[39] & b[55])^(a[38] & b[56])^(a[37] & b[57])^(a[36] & b[58])^(a[35] & b[59])^(a[34] & b[60])^(a[33] & b[61])^(a[32] & b[62])^(a[31] & b[63])^(a[30] & b[64])^(a[29] & b[65])^(a[28] & b[66])^(a[27] & b[67])^(a[26] & b[68])^(a[25] & b[69])^(a[24] & b[70])^(a[23] & b[71])^(a[22] & b[72])^(a[21] & b[73])^(a[20] & b[74])^(a[19] & b[75])^(a[18] & b[76])^(a[17] & b[77])^(a[16] & b[78])^(a[15] & b[79])^(a[14] & b[80])^(a[13] & b[81])^(a[12] & b[82])^(a[11] & b[83])^(a[10] & b[84])^(a[9] & b[85])^(a[8] & b[86])^(a[7] & b[87])^(a[6] & b[88])^(a[5] & b[89])^(a[4] & b[90])^(a[3] & b[91])^(a[2] & b[92])^(a[1] & b[93])^(a[0] & b[94]);
assign y[95] = (a[95] & b[0])^(a[94] & b[1])^(a[93] & b[2])^(a[92] & b[3])^(a[91] & b[4])^(a[90] & b[5])^(a[89] & b[6])^(a[88] & b[7])^(a[87] & b[8])^(a[86] & b[9])^(a[85] & b[10])^(a[84] & b[11])^(a[83] & b[12])^(a[82] & b[13])^(a[81] & b[14])^(a[80] & b[15])^(a[79] & b[16])^(a[78] & b[17])^(a[77] & b[18])^(a[76] & b[19])^(a[75] & b[20])^(a[74] & b[21])^(a[73] & b[22])^(a[72] & b[23])^(a[71] & b[24])^(a[70] & b[25])^(a[69] & b[26])^(a[68] & b[27])^(a[67] & b[28])^(a[66] & b[29])^(a[65] & b[30])^(a[64] & b[31])^(a[63] & b[32])^(a[62] & b[33])^(a[61] & b[34])^(a[60] & b[35])^(a[59] & b[36])^(a[58] & b[37])^(a[57] & b[38])^(a[56] & b[39])^(a[55] & b[40])^(a[54] & b[41])^(a[53] & b[42])^(a[52] & b[43])^(a[51] & b[44])^(a[50] & b[45])^(a[49] & b[46])^(a[48] & b[47])^(a[47] & b[48])^(a[46] & b[49])^(a[45] & b[50])^(a[44] & b[51])^(a[43] & b[52])^(a[42] & b[53])^(a[41] & b[54])^(a[40] & b[55])^(a[39] & b[56])^(a[38] & b[57])^(a[37] & b[58])^(a[36] & b[59])^(a[35] & b[60])^(a[34] & b[61])^(a[33] & b[62])^(a[32] & b[63])^(a[31] & b[64])^(a[30] & b[65])^(a[29] & b[66])^(a[28] & b[67])^(a[27] & b[68])^(a[26] & b[69])^(a[25] & b[70])^(a[24] & b[71])^(a[23] & b[72])^(a[22] & b[73])^(a[21] & b[74])^(a[20] & b[75])^(a[19] & b[76])^(a[18] & b[77])^(a[17] & b[78])^(a[16] & b[79])^(a[15] & b[80])^(a[14] & b[81])^(a[13] & b[82])^(a[12] & b[83])^(a[11] & b[84])^(a[10] & b[85])^(a[9] & b[86])^(a[8] & b[87])^(a[7] & b[88])^(a[6] & b[89])^(a[5] & b[90])^(a[4] & b[91])^(a[3] & b[92])^(a[2] & b[93])^(a[1] & b[94])^(a[0] & b[95]);
assign y[96] = (a[96] & b[0])^(a[95] & b[1])^(a[94] & b[2])^(a[93] & b[3])^(a[92] & b[4])^(a[91] & b[5])^(a[90] & b[6])^(a[89] & b[7])^(a[88] & b[8])^(a[87] & b[9])^(a[86] & b[10])^(a[85] & b[11])^(a[84] & b[12])^(a[83] & b[13])^(a[82] & b[14])^(a[81] & b[15])^(a[80] & b[16])^(a[79] & b[17])^(a[78] & b[18])^(a[77] & b[19])^(a[76] & b[20])^(a[75] & b[21])^(a[74] & b[22])^(a[73] & b[23])^(a[72] & b[24])^(a[71] & b[25])^(a[70] & b[26])^(a[69] & b[27])^(a[68] & b[28])^(a[67] & b[29])^(a[66] & b[30])^(a[65] & b[31])^(a[64] & b[32])^(a[63] & b[33])^(a[62] & b[34])^(a[61] & b[35])^(a[60] & b[36])^(a[59] & b[37])^(a[58] & b[38])^(a[57] & b[39])^(a[56] & b[40])^(a[55] & b[41])^(a[54] & b[42])^(a[53] & b[43])^(a[52] & b[44])^(a[51] & b[45])^(a[50] & b[46])^(a[49] & b[47])^(a[48] & b[48])^(a[47] & b[49])^(a[46] & b[50])^(a[45] & b[51])^(a[44] & b[52])^(a[43] & b[53])^(a[42] & b[54])^(a[41] & b[55])^(a[40] & b[56])^(a[39] & b[57])^(a[38] & b[58])^(a[37] & b[59])^(a[36] & b[60])^(a[35] & b[61])^(a[34] & b[62])^(a[33] & b[63])^(a[32] & b[64])^(a[31] & b[65])^(a[30] & b[66])^(a[29] & b[67])^(a[28] & b[68])^(a[27] & b[69])^(a[26] & b[70])^(a[25] & b[71])^(a[24] & b[72])^(a[23] & b[73])^(a[22] & b[74])^(a[21] & b[75])^(a[20] & b[76])^(a[19] & b[77])^(a[18] & b[78])^(a[17] & b[79])^(a[16] & b[80])^(a[15] & b[81])^(a[14] & b[82])^(a[13] & b[83])^(a[12] & b[84])^(a[11] & b[85])^(a[10] & b[86])^(a[9] & b[87])^(a[8] & b[88])^(a[7] & b[89])^(a[6] & b[90])^(a[5] & b[91])^(a[4] & b[92])^(a[3] & b[93])^(a[2] & b[94])^(a[1] & b[95])^(a[0] & b[96]);
assign y[97] = (a[97] & b[0])^(a[96] & b[1])^(a[95] & b[2])^(a[94] & b[3])^(a[93] & b[4])^(a[92] & b[5])^(a[91] & b[6])^(a[90] & b[7])^(a[89] & b[8])^(a[88] & b[9])^(a[87] & b[10])^(a[86] & b[11])^(a[85] & b[12])^(a[84] & b[13])^(a[83] & b[14])^(a[82] & b[15])^(a[81] & b[16])^(a[80] & b[17])^(a[79] & b[18])^(a[78] & b[19])^(a[77] & b[20])^(a[76] & b[21])^(a[75] & b[22])^(a[74] & b[23])^(a[73] & b[24])^(a[72] & b[25])^(a[71] & b[26])^(a[70] & b[27])^(a[69] & b[28])^(a[68] & b[29])^(a[67] & b[30])^(a[66] & b[31])^(a[65] & b[32])^(a[64] & b[33])^(a[63] & b[34])^(a[62] & b[35])^(a[61] & b[36])^(a[60] & b[37])^(a[59] & b[38])^(a[58] & b[39])^(a[57] & b[40])^(a[56] & b[41])^(a[55] & b[42])^(a[54] & b[43])^(a[53] & b[44])^(a[52] & b[45])^(a[51] & b[46])^(a[50] & b[47])^(a[49] & b[48])^(a[48] & b[49])^(a[47] & b[50])^(a[46] & b[51])^(a[45] & b[52])^(a[44] & b[53])^(a[43] & b[54])^(a[42] & b[55])^(a[41] & b[56])^(a[40] & b[57])^(a[39] & b[58])^(a[38] & b[59])^(a[37] & b[60])^(a[36] & b[61])^(a[35] & b[62])^(a[34] & b[63])^(a[33] & b[64])^(a[32] & b[65])^(a[31] & b[66])^(a[30] & b[67])^(a[29] & b[68])^(a[28] & b[69])^(a[27] & b[70])^(a[26] & b[71])^(a[25] & b[72])^(a[24] & b[73])^(a[23] & b[74])^(a[22] & b[75])^(a[21] & b[76])^(a[20] & b[77])^(a[19] & b[78])^(a[18] & b[79])^(a[17] & b[80])^(a[16] & b[81])^(a[15] & b[82])^(a[14] & b[83])^(a[13] & b[84])^(a[12] & b[85])^(a[11] & b[86])^(a[10] & b[87])^(a[9] & b[88])^(a[8] & b[89])^(a[7] & b[90])^(a[6] & b[91])^(a[5] & b[92])^(a[4] & b[93])^(a[3] & b[94])^(a[2] & b[95])^(a[1] & b[96])^(a[0] & b[97]);
assign y[98] = (a[98] & b[0])^(a[97] & b[1])^(a[96] & b[2])^(a[95] & b[3])^(a[94] & b[4])^(a[93] & b[5])^(a[92] & b[6])^(a[91] & b[7])^(a[90] & b[8])^(a[89] & b[9])^(a[88] & b[10])^(a[87] & b[11])^(a[86] & b[12])^(a[85] & b[13])^(a[84] & b[14])^(a[83] & b[15])^(a[82] & b[16])^(a[81] & b[17])^(a[80] & b[18])^(a[79] & b[19])^(a[78] & b[20])^(a[77] & b[21])^(a[76] & b[22])^(a[75] & b[23])^(a[74] & b[24])^(a[73] & b[25])^(a[72] & b[26])^(a[71] & b[27])^(a[70] & b[28])^(a[69] & b[29])^(a[68] & b[30])^(a[67] & b[31])^(a[66] & b[32])^(a[65] & b[33])^(a[64] & b[34])^(a[63] & b[35])^(a[62] & b[36])^(a[61] & b[37])^(a[60] & b[38])^(a[59] & b[39])^(a[58] & b[40])^(a[57] & b[41])^(a[56] & b[42])^(a[55] & b[43])^(a[54] & b[44])^(a[53] & b[45])^(a[52] & b[46])^(a[51] & b[47])^(a[50] & b[48])^(a[49] & b[49])^(a[48] & b[50])^(a[47] & b[51])^(a[46] & b[52])^(a[45] & b[53])^(a[44] & b[54])^(a[43] & b[55])^(a[42] & b[56])^(a[41] & b[57])^(a[40] & b[58])^(a[39] & b[59])^(a[38] & b[60])^(a[37] & b[61])^(a[36] & b[62])^(a[35] & b[63])^(a[34] & b[64])^(a[33] & b[65])^(a[32] & b[66])^(a[31] & b[67])^(a[30] & b[68])^(a[29] & b[69])^(a[28] & b[70])^(a[27] & b[71])^(a[26] & b[72])^(a[25] & b[73])^(a[24] & b[74])^(a[23] & b[75])^(a[22] & b[76])^(a[21] & b[77])^(a[20] & b[78])^(a[19] & b[79])^(a[18] & b[80])^(a[17] & b[81])^(a[16] & b[82])^(a[15] & b[83])^(a[14] & b[84])^(a[13] & b[85])^(a[12] & b[86])^(a[11] & b[87])^(a[10] & b[88])^(a[9] & b[89])^(a[8] & b[90])^(a[7] & b[91])^(a[6] & b[92])^(a[5] & b[93])^(a[4] & b[94])^(a[3] & b[95])^(a[2] & b[96])^(a[1] & b[97])^(a[0] & b[98]);
assign y[99] = (a[99] & b[0])^(a[98] & b[1])^(a[97] & b[2])^(a[96] & b[3])^(a[95] & b[4])^(a[94] & b[5])^(a[93] & b[6])^(a[92] & b[7])^(a[91] & b[8])^(a[90] & b[9])^(a[89] & b[10])^(a[88] & b[11])^(a[87] & b[12])^(a[86] & b[13])^(a[85] & b[14])^(a[84] & b[15])^(a[83] & b[16])^(a[82] & b[17])^(a[81] & b[18])^(a[80] & b[19])^(a[79] & b[20])^(a[78] & b[21])^(a[77] & b[22])^(a[76] & b[23])^(a[75] & b[24])^(a[74] & b[25])^(a[73] & b[26])^(a[72] & b[27])^(a[71] & b[28])^(a[70] & b[29])^(a[69] & b[30])^(a[68] & b[31])^(a[67] & b[32])^(a[66] & b[33])^(a[65] & b[34])^(a[64] & b[35])^(a[63] & b[36])^(a[62] & b[37])^(a[61] & b[38])^(a[60] & b[39])^(a[59] & b[40])^(a[58] & b[41])^(a[57] & b[42])^(a[56] & b[43])^(a[55] & b[44])^(a[54] & b[45])^(a[53] & b[46])^(a[52] & b[47])^(a[51] & b[48])^(a[50] & b[49])^(a[49] & b[50])^(a[48] & b[51])^(a[47] & b[52])^(a[46] & b[53])^(a[45] & b[54])^(a[44] & b[55])^(a[43] & b[56])^(a[42] & b[57])^(a[41] & b[58])^(a[40] & b[59])^(a[39] & b[60])^(a[38] & b[61])^(a[37] & b[62])^(a[36] & b[63])^(a[35] & b[64])^(a[34] & b[65])^(a[33] & b[66])^(a[32] & b[67])^(a[31] & b[68])^(a[30] & b[69])^(a[29] & b[70])^(a[28] & b[71])^(a[27] & b[72])^(a[26] & b[73])^(a[25] & b[74])^(a[24] & b[75])^(a[23] & b[76])^(a[22] & b[77])^(a[21] & b[78])^(a[20] & b[79])^(a[19] & b[80])^(a[18] & b[81])^(a[17] & b[82])^(a[16] & b[83])^(a[15] & b[84])^(a[14] & b[85])^(a[13] & b[86])^(a[12] & b[87])^(a[11] & b[88])^(a[10] & b[89])^(a[9] & b[90])^(a[8] & b[91])^(a[7] & b[92])^(a[6] & b[93])^(a[5] & b[94])^(a[4] & b[95])^(a[3] & b[96])^(a[2] & b[97])^(a[1] & b[98])^(a[0] & b[99]);
assign y[100] = (a[100] & b[0])^(a[99] & b[1])^(a[98] & b[2])^(a[97] & b[3])^(a[96] & b[4])^(a[95] & b[5])^(a[94] & b[6])^(a[93] & b[7])^(a[92] & b[8])^(a[91] & b[9])^(a[90] & b[10])^(a[89] & b[11])^(a[88] & b[12])^(a[87] & b[13])^(a[86] & b[14])^(a[85] & b[15])^(a[84] & b[16])^(a[83] & b[17])^(a[82] & b[18])^(a[81] & b[19])^(a[80] & b[20])^(a[79] & b[21])^(a[78] & b[22])^(a[77] & b[23])^(a[76] & b[24])^(a[75] & b[25])^(a[74] & b[26])^(a[73] & b[27])^(a[72] & b[28])^(a[71] & b[29])^(a[70] & b[30])^(a[69] & b[31])^(a[68] & b[32])^(a[67] & b[33])^(a[66] & b[34])^(a[65] & b[35])^(a[64] & b[36])^(a[63] & b[37])^(a[62] & b[38])^(a[61] & b[39])^(a[60] & b[40])^(a[59] & b[41])^(a[58] & b[42])^(a[57] & b[43])^(a[56] & b[44])^(a[55] & b[45])^(a[54] & b[46])^(a[53] & b[47])^(a[52] & b[48])^(a[51] & b[49])^(a[50] & b[50])^(a[49] & b[51])^(a[48] & b[52])^(a[47] & b[53])^(a[46] & b[54])^(a[45] & b[55])^(a[44] & b[56])^(a[43] & b[57])^(a[42] & b[58])^(a[41] & b[59])^(a[40] & b[60])^(a[39] & b[61])^(a[38] & b[62])^(a[37] & b[63])^(a[36] & b[64])^(a[35] & b[65])^(a[34] & b[66])^(a[33] & b[67])^(a[32] & b[68])^(a[31] & b[69])^(a[30] & b[70])^(a[29] & b[71])^(a[28] & b[72])^(a[27] & b[73])^(a[26] & b[74])^(a[25] & b[75])^(a[24] & b[76])^(a[23] & b[77])^(a[22] & b[78])^(a[21] & b[79])^(a[20] & b[80])^(a[19] & b[81])^(a[18] & b[82])^(a[17] & b[83])^(a[16] & b[84])^(a[15] & b[85])^(a[14] & b[86])^(a[13] & b[87])^(a[12] & b[88])^(a[11] & b[89])^(a[10] & b[90])^(a[9] & b[91])^(a[8] & b[92])^(a[7] & b[93])^(a[6] & b[94])^(a[5] & b[95])^(a[4] & b[96])^(a[3] & b[97])^(a[2] & b[98])^(a[1] & b[99])^(a[0] & b[100]);
assign y[101] = (a[101] & b[0])^(a[100] & b[1])^(a[99] & b[2])^(a[98] & b[3])^(a[97] & b[4])^(a[96] & b[5])^(a[95] & b[6])^(a[94] & b[7])^(a[93] & b[8])^(a[92] & b[9])^(a[91] & b[10])^(a[90] & b[11])^(a[89] & b[12])^(a[88] & b[13])^(a[87] & b[14])^(a[86] & b[15])^(a[85] & b[16])^(a[84] & b[17])^(a[83] & b[18])^(a[82] & b[19])^(a[81] & b[20])^(a[80] & b[21])^(a[79] & b[22])^(a[78] & b[23])^(a[77] & b[24])^(a[76] & b[25])^(a[75] & b[26])^(a[74] & b[27])^(a[73] & b[28])^(a[72] & b[29])^(a[71] & b[30])^(a[70] & b[31])^(a[69] & b[32])^(a[68] & b[33])^(a[67] & b[34])^(a[66] & b[35])^(a[65] & b[36])^(a[64] & b[37])^(a[63] & b[38])^(a[62] & b[39])^(a[61] & b[40])^(a[60] & b[41])^(a[59] & b[42])^(a[58] & b[43])^(a[57] & b[44])^(a[56] & b[45])^(a[55] & b[46])^(a[54] & b[47])^(a[53] & b[48])^(a[52] & b[49])^(a[51] & b[50])^(a[50] & b[51])^(a[49] & b[52])^(a[48] & b[53])^(a[47] & b[54])^(a[46] & b[55])^(a[45] & b[56])^(a[44] & b[57])^(a[43] & b[58])^(a[42] & b[59])^(a[41] & b[60])^(a[40] & b[61])^(a[39] & b[62])^(a[38] & b[63])^(a[37] & b[64])^(a[36] & b[65])^(a[35] & b[66])^(a[34] & b[67])^(a[33] & b[68])^(a[32] & b[69])^(a[31] & b[70])^(a[30] & b[71])^(a[29] & b[72])^(a[28] & b[73])^(a[27] & b[74])^(a[26] & b[75])^(a[25] & b[76])^(a[24] & b[77])^(a[23] & b[78])^(a[22] & b[79])^(a[21] & b[80])^(a[20] & b[81])^(a[19] & b[82])^(a[18] & b[83])^(a[17] & b[84])^(a[16] & b[85])^(a[15] & b[86])^(a[14] & b[87])^(a[13] & b[88])^(a[12] & b[89])^(a[11] & b[90])^(a[10] & b[91])^(a[9] & b[92])^(a[8] & b[93])^(a[7] & b[94])^(a[6] & b[95])^(a[5] & b[96])^(a[4] & b[97])^(a[3] & b[98])^(a[2] & b[99])^(a[1] & b[100])^(a[0] & b[101]);
assign y[102] = (a[102] & b[0])^(a[101] & b[1])^(a[100] & b[2])^(a[99] & b[3])^(a[98] & b[4])^(a[97] & b[5])^(a[96] & b[6])^(a[95] & b[7])^(a[94] & b[8])^(a[93] & b[9])^(a[92] & b[10])^(a[91] & b[11])^(a[90] & b[12])^(a[89] & b[13])^(a[88] & b[14])^(a[87] & b[15])^(a[86] & b[16])^(a[85] & b[17])^(a[84] & b[18])^(a[83] & b[19])^(a[82] & b[20])^(a[81] & b[21])^(a[80] & b[22])^(a[79] & b[23])^(a[78] & b[24])^(a[77] & b[25])^(a[76] & b[26])^(a[75] & b[27])^(a[74] & b[28])^(a[73] & b[29])^(a[72] & b[30])^(a[71] & b[31])^(a[70] & b[32])^(a[69] & b[33])^(a[68] & b[34])^(a[67] & b[35])^(a[66] & b[36])^(a[65] & b[37])^(a[64] & b[38])^(a[63] & b[39])^(a[62] & b[40])^(a[61] & b[41])^(a[60] & b[42])^(a[59] & b[43])^(a[58] & b[44])^(a[57] & b[45])^(a[56] & b[46])^(a[55] & b[47])^(a[54] & b[48])^(a[53] & b[49])^(a[52] & b[50])^(a[51] & b[51])^(a[50] & b[52])^(a[49] & b[53])^(a[48] & b[54])^(a[47] & b[55])^(a[46] & b[56])^(a[45] & b[57])^(a[44] & b[58])^(a[43] & b[59])^(a[42] & b[60])^(a[41] & b[61])^(a[40] & b[62])^(a[39] & b[63])^(a[38] & b[64])^(a[37] & b[65])^(a[36] & b[66])^(a[35] & b[67])^(a[34] & b[68])^(a[33] & b[69])^(a[32] & b[70])^(a[31] & b[71])^(a[30] & b[72])^(a[29] & b[73])^(a[28] & b[74])^(a[27] & b[75])^(a[26] & b[76])^(a[25] & b[77])^(a[24] & b[78])^(a[23] & b[79])^(a[22] & b[80])^(a[21] & b[81])^(a[20] & b[82])^(a[19] & b[83])^(a[18] & b[84])^(a[17] & b[85])^(a[16] & b[86])^(a[15] & b[87])^(a[14] & b[88])^(a[13] & b[89])^(a[12] & b[90])^(a[11] & b[91])^(a[10] & b[92])^(a[9] & b[93])^(a[8] & b[94])^(a[7] & b[95])^(a[6] & b[96])^(a[5] & b[97])^(a[4] & b[98])^(a[3] & b[99])^(a[2] & b[100])^(a[1] & b[101])^(a[0] & b[102]);
assign y[103] = (a[103] & b[0])^(a[102] & b[1])^(a[101] & b[2])^(a[100] & b[3])^(a[99] & b[4])^(a[98] & b[5])^(a[97] & b[6])^(a[96] & b[7])^(a[95] & b[8])^(a[94] & b[9])^(a[93] & b[10])^(a[92] & b[11])^(a[91] & b[12])^(a[90] & b[13])^(a[89] & b[14])^(a[88] & b[15])^(a[87] & b[16])^(a[86] & b[17])^(a[85] & b[18])^(a[84] & b[19])^(a[83] & b[20])^(a[82] & b[21])^(a[81] & b[22])^(a[80] & b[23])^(a[79] & b[24])^(a[78] & b[25])^(a[77] & b[26])^(a[76] & b[27])^(a[75] & b[28])^(a[74] & b[29])^(a[73] & b[30])^(a[72] & b[31])^(a[71] & b[32])^(a[70] & b[33])^(a[69] & b[34])^(a[68] & b[35])^(a[67] & b[36])^(a[66] & b[37])^(a[65] & b[38])^(a[64] & b[39])^(a[63] & b[40])^(a[62] & b[41])^(a[61] & b[42])^(a[60] & b[43])^(a[59] & b[44])^(a[58] & b[45])^(a[57] & b[46])^(a[56] & b[47])^(a[55] & b[48])^(a[54] & b[49])^(a[53] & b[50])^(a[52] & b[51])^(a[51] & b[52])^(a[50] & b[53])^(a[49] & b[54])^(a[48] & b[55])^(a[47] & b[56])^(a[46] & b[57])^(a[45] & b[58])^(a[44] & b[59])^(a[43] & b[60])^(a[42] & b[61])^(a[41] & b[62])^(a[40] & b[63])^(a[39] & b[64])^(a[38] & b[65])^(a[37] & b[66])^(a[36] & b[67])^(a[35] & b[68])^(a[34] & b[69])^(a[33] & b[70])^(a[32] & b[71])^(a[31] & b[72])^(a[30] & b[73])^(a[29] & b[74])^(a[28] & b[75])^(a[27] & b[76])^(a[26] & b[77])^(a[25] & b[78])^(a[24] & b[79])^(a[23] & b[80])^(a[22] & b[81])^(a[21] & b[82])^(a[20] & b[83])^(a[19] & b[84])^(a[18] & b[85])^(a[17] & b[86])^(a[16] & b[87])^(a[15] & b[88])^(a[14] & b[89])^(a[13] & b[90])^(a[12] & b[91])^(a[11] & b[92])^(a[10] & b[93])^(a[9] & b[94])^(a[8] & b[95])^(a[7] & b[96])^(a[6] & b[97])^(a[5] & b[98])^(a[4] & b[99])^(a[3] & b[100])^(a[2] & b[101])^(a[1] & b[102])^(a[0] & b[103]);
assign y[104] = (a[104] & b[0])^(a[103] & b[1])^(a[102] & b[2])^(a[101] & b[3])^(a[100] & b[4])^(a[99] & b[5])^(a[98] & b[6])^(a[97] & b[7])^(a[96] & b[8])^(a[95] & b[9])^(a[94] & b[10])^(a[93] & b[11])^(a[92] & b[12])^(a[91] & b[13])^(a[90] & b[14])^(a[89] & b[15])^(a[88] & b[16])^(a[87] & b[17])^(a[86] & b[18])^(a[85] & b[19])^(a[84] & b[20])^(a[83] & b[21])^(a[82] & b[22])^(a[81] & b[23])^(a[80] & b[24])^(a[79] & b[25])^(a[78] & b[26])^(a[77] & b[27])^(a[76] & b[28])^(a[75] & b[29])^(a[74] & b[30])^(a[73] & b[31])^(a[72] & b[32])^(a[71] & b[33])^(a[70] & b[34])^(a[69] & b[35])^(a[68] & b[36])^(a[67] & b[37])^(a[66] & b[38])^(a[65] & b[39])^(a[64] & b[40])^(a[63] & b[41])^(a[62] & b[42])^(a[61] & b[43])^(a[60] & b[44])^(a[59] & b[45])^(a[58] & b[46])^(a[57] & b[47])^(a[56] & b[48])^(a[55] & b[49])^(a[54] & b[50])^(a[53] & b[51])^(a[52] & b[52])^(a[51] & b[53])^(a[50] & b[54])^(a[49] & b[55])^(a[48] & b[56])^(a[47] & b[57])^(a[46] & b[58])^(a[45] & b[59])^(a[44] & b[60])^(a[43] & b[61])^(a[42] & b[62])^(a[41] & b[63])^(a[40] & b[64])^(a[39] & b[65])^(a[38] & b[66])^(a[37] & b[67])^(a[36] & b[68])^(a[35] & b[69])^(a[34] & b[70])^(a[33] & b[71])^(a[32] & b[72])^(a[31] & b[73])^(a[30] & b[74])^(a[29] & b[75])^(a[28] & b[76])^(a[27] & b[77])^(a[26] & b[78])^(a[25] & b[79])^(a[24] & b[80])^(a[23] & b[81])^(a[22] & b[82])^(a[21] & b[83])^(a[20] & b[84])^(a[19] & b[85])^(a[18] & b[86])^(a[17] & b[87])^(a[16] & b[88])^(a[15] & b[89])^(a[14] & b[90])^(a[13] & b[91])^(a[12] & b[92])^(a[11] & b[93])^(a[10] & b[94])^(a[9] & b[95])^(a[8] & b[96])^(a[7] & b[97])^(a[6] & b[98])^(a[5] & b[99])^(a[4] & b[100])^(a[3] & b[101])^(a[2] & b[102])^(a[1] & b[103])^(a[0] & b[104]);
assign y[105] = (a[105] & b[0])^(a[104] & b[1])^(a[103] & b[2])^(a[102] & b[3])^(a[101] & b[4])^(a[100] & b[5])^(a[99] & b[6])^(a[98] & b[7])^(a[97] & b[8])^(a[96] & b[9])^(a[95] & b[10])^(a[94] & b[11])^(a[93] & b[12])^(a[92] & b[13])^(a[91] & b[14])^(a[90] & b[15])^(a[89] & b[16])^(a[88] & b[17])^(a[87] & b[18])^(a[86] & b[19])^(a[85] & b[20])^(a[84] & b[21])^(a[83] & b[22])^(a[82] & b[23])^(a[81] & b[24])^(a[80] & b[25])^(a[79] & b[26])^(a[78] & b[27])^(a[77] & b[28])^(a[76] & b[29])^(a[75] & b[30])^(a[74] & b[31])^(a[73] & b[32])^(a[72] & b[33])^(a[71] & b[34])^(a[70] & b[35])^(a[69] & b[36])^(a[68] & b[37])^(a[67] & b[38])^(a[66] & b[39])^(a[65] & b[40])^(a[64] & b[41])^(a[63] & b[42])^(a[62] & b[43])^(a[61] & b[44])^(a[60] & b[45])^(a[59] & b[46])^(a[58] & b[47])^(a[57] & b[48])^(a[56] & b[49])^(a[55] & b[50])^(a[54] & b[51])^(a[53] & b[52])^(a[52] & b[53])^(a[51] & b[54])^(a[50] & b[55])^(a[49] & b[56])^(a[48] & b[57])^(a[47] & b[58])^(a[46] & b[59])^(a[45] & b[60])^(a[44] & b[61])^(a[43] & b[62])^(a[42] & b[63])^(a[41] & b[64])^(a[40] & b[65])^(a[39] & b[66])^(a[38] & b[67])^(a[37] & b[68])^(a[36] & b[69])^(a[35] & b[70])^(a[34] & b[71])^(a[33] & b[72])^(a[32] & b[73])^(a[31] & b[74])^(a[30] & b[75])^(a[29] & b[76])^(a[28] & b[77])^(a[27] & b[78])^(a[26] & b[79])^(a[25] & b[80])^(a[24] & b[81])^(a[23] & b[82])^(a[22] & b[83])^(a[21] & b[84])^(a[20] & b[85])^(a[19] & b[86])^(a[18] & b[87])^(a[17] & b[88])^(a[16] & b[89])^(a[15] & b[90])^(a[14] & b[91])^(a[13] & b[92])^(a[12] & b[93])^(a[11] & b[94])^(a[10] & b[95])^(a[9] & b[96])^(a[8] & b[97])^(a[7] & b[98])^(a[6] & b[99])^(a[5] & b[100])^(a[4] & b[101])^(a[3] & b[102])^(a[2] & b[103])^(a[1] & b[104])^(a[0] & b[105]);
assign y[106] = (a[106] & b[0])^(a[105] & b[1])^(a[104] & b[2])^(a[103] & b[3])^(a[102] & b[4])^(a[101] & b[5])^(a[100] & b[6])^(a[99] & b[7])^(a[98] & b[8])^(a[97] & b[9])^(a[96] & b[10])^(a[95] & b[11])^(a[94] & b[12])^(a[93] & b[13])^(a[92] & b[14])^(a[91] & b[15])^(a[90] & b[16])^(a[89] & b[17])^(a[88] & b[18])^(a[87] & b[19])^(a[86] & b[20])^(a[85] & b[21])^(a[84] & b[22])^(a[83] & b[23])^(a[82] & b[24])^(a[81] & b[25])^(a[80] & b[26])^(a[79] & b[27])^(a[78] & b[28])^(a[77] & b[29])^(a[76] & b[30])^(a[75] & b[31])^(a[74] & b[32])^(a[73] & b[33])^(a[72] & b[34])^(a[71] & b[35])^(a[70] & b[36])^(a[69] & b[37])^(a[68] & b[38])^(a[67] & b[39])^(a[66] & b[40])^(a[65] & b[41])^(a[64] & b[42])^(a[63] & b[43])^(a[62] & b[44])^(a[61] & b[45])^(a[60] & b[46])^(a[59] & b[47])^(a[58] & b[48])^(a[57] & b[49])^(a[56] & b[50])^(a[55] & b[51])^(a[54] & b[52])^(a[53] & b[53])^(a[52] & b[54])^(a[51] & b[55])^(a[50] & b[56])^(a[49] & b[57])^(a[48] & b[58])^(a[47] & b[59])^(a[46] & b[60])^(a[45] & b[61])^(a[44] & b[62])^(a[43] & b[63])^(a[42] & b[64])^(a[41] & b[65])^(a[40] & b[66])^(a[39] & b[67])^(a[38] & b[68])^(a[37] & b[69])^(a[36] & b[70])^(a[35] & b[71])^(a[34] & b[72])^(a[33] & b[73])^(a[32] & b[74])^(a[31] & b[75])^(a[30] & b[76])^(a[29] & b[77])^(a[28] & b[78])^(a[27] & b[79])^(a[26] & b[80])^(a[25] & b[81])^(a[24] & b[82])^(a[23] & b[83])^(a[22] & b[84])^(a[21] & b[85])^(a[20] & b[86])^(a[19] & b[87])^(a[18] & b[88])^(a[17] & b[89])^(a[16] & b[90])^(a[15] & b[91])^(a[14] & b[92])^(a[13] & b[93])^(a[12] & b[94])^(a[11] & b[95])^(a[10] & b[96])^(a[9] & b[97])^(a[8] & b[98])^(a[7] & b[99])^(a[6] & b[100])^(a[5] & b[101])^(a[4] & b[102])^(a[3] & b[103])^(a[2] & b[104])^(a[1] & b[105])^(a[0] & b[106]);
assign y[107] = (a[107] & b[0])^(a[106] & b[1])^(a[105] & b[2])^(a[104] & b[3])^(a[103] & b[4])^(a[102] & b[5])^(a[101] & b[6])^(a[100] & b[7])^(a[99] & b[8])^(a[98] & b[9])^(a[97] & b[10])^(a[96] & b[11])^(a[95] & b[12])^(a[94] & b[13])^(a[93] & b[14])^(a[92] & b[15])^(a[91] & b[16])^(a[90] & b[17])^(a[89] & b[18])^(a[88] & b[19])^(a[87] & b[20])^(a[86] & b[21])^(a[85] & b[22])^(a[84] & b[23])^(a[83] & b[24])^(a[82] & b[25])^(a[81] & b[26])^(a[80] & b[27])^(a[79] & b[28])^(a[78] & b[29])^(a[77] & b[30])^(a[76] & b[31])^(a[75] & b[32])^(a[74] & b[33])^(a[73] & b[34])^(a[72] & b[35])^(a[71] & b[36])^(a[70] & b[37])^(a[69] & b[38])^(a[68] & b[39])^(a[67] & b[40])^(a[66] & b[41])^(a[65] & b[42])^(a[64] & b[43])^(a[63] & b[44])^(a[62] & b[45])^(a[61] & b[46])^(a[60] & b[47])^(a[59] & b[48])^(a[58] & b[49])^(a[57] & b[50])^(a[56] & b[51])^(a[55] & b[52])^(a[54] & b[53])^(a[53] & b[54])^(a[52] & b[55])^(a[51] & b[56])^(a[50] & b[57])^(a[49] & b[58])^(a[48] & b[59])^(a[47] & b[60])^(a[46] & b[61])^(a[45] & b[62])^(a[44] & b[63])^(a[43] & b[64])^(a[42] & b[65])^(a[41] & b[66])^(a[40] & b[67])^(a[39] & b[68])^(a[38] & b[69])^(a[37] & b[70])^(a[36] & b[71])^(a[35] & b[72])^(a[34] & b[73])^(a[33] & b[74])^(a[32] & b[75])^(a[31] & b[76])^(a[30] & b[77])^(a[29] & b[78])^(a[28] & b[79])^(a[27] & b[80])^(a[26] & b[81])^(a[25] & b[82])^(a[24] & b[83])^(a[23] & b[84])^(a[22] & b[85])^(a[21] & b[86])^(a[20] & b[87])^(a[19] & b[88])^(a[18] & b[89])^(a[17] & b[90])^(a[16] & b[91])^(a[15] & b[92])^(a[14] & b[93])^(a[13] & b[94])^(a[12] & b[95])^(a[11] & b[96])^(a[10] & b[97])^(a[9] & b[98])^(a[8] & b[99])^(a[7] & b[100])^(a[6] & b[101])^(a[5] & b[102])^(a[4] & b[103])^(a[3] & b[104])^(a[2] & b[105])^(a[1] & b[106])^(a[0] & b[107]);
assign y[108] = (a[108] & b[0])^(a[107] & b[1])^(a[106] & b[2])^(a[105] & b[3])^(a[104] & b[4])^(a[103] & b[5])^(a[102] & b[6])^(a[101] & b[7])^(a[100] & b[8])^(a[99] & b[9])^(a[98] & b[10])^(a[97] & b[11])^(a[96] & b[12])^(a[95] & b[13])^(a[94] & b[14])^(a[93] & b[15])^(a[92] & b[16])^(a[91] & b[17])^(a[90] & b[18])^(a[89] & b[19])^(a[88] & b[20])^(a[87] & b[21])^(a[86] & b[22])^(a[85] & b[23])^(a[84] & b[24])^(a[83] & b[25])^(a[82] & b[26])^(a[81] & b[27])^(a[80] & b[28])^(a[79] & b[29])^(a[78] & b[30])^(a[77] & b[31])^(a[76] & b[32])^(a[75] & b[33])^(a[74] & b[34])^(a[73] & b[35])^(a[72] & b[36])^(a[71] & b[37])^(a[70] & b[38])^(a[69] & b[39])^(a[68] & b[40])^(a[67] & b[41])^(a[66] & b[42])^(a[65] & b[43])^(a[64] & b[44])^(a[63] & b[45])^(a[62] & b[46])^(a[61] & b[47])^(a[60] & b[48])^(a[59] & b[49])^(a[58] & b[50])^(a[57] & b[51])^(a[56] & b[52])^(a[55] & b[53])^(a[54] & b[54])^(a[53] & b[55])^(a[52] & b[56])^(a[51] & b[57])^(a[50] & b[58])^(a[49] & b[59])^(a[48] & b[60])^(a[47] & b[61])^(a[46] & b[62])^(a[45] & b[63])^(a[44] & b[64])^(a[43] & b[65])^(a[42] & b[66])^(a[41] & b[67])^(a[40] & b[68])^(a[39] & b[69])^(a[38] & b[70])^(a[37] & b[71])^(a[36] & b[72])^(a[35] & b[73])^(a[34] & b[74])^(a[33] & b[75])^(a[32] & b[76])^(a[31] & b[77])^(a[30] & b[78])^(a[29] & b[79])^(a[28] & b[80])^(a[27] & b[81])^(a[26] & b[82])^(a[25] & b[83])^(a[24] & b[84])^(a[23] & b[85])^(a[22] & b[86])^(a[21] & b[87])^(a[20] & b[88])^(a[19] & b[89])^(a[18] & b[90])^(a[17] & b[91])^(a[16] & b[92])^(a[15] & b[93])^(a[14] & b[94])^(a[13] & b[95])^(a[12] & b[96])^(a[11] & b[97])^(a[10] & b[98])^(a[9] & b[99])^(a[8] & b[100])^(a[7] & b[101])^(a[6] & b[102])^(a[5] & b[103])^(a[4] & b[104])^(a[3] & b[105])^(a[2] & b[106])^(a[1] & b[107])^(a[0] & b[108]);
assign y[109] = (a[109] & b[0])^(a[108] & b[1])^(a[107] & b[2])^(a[106] & b[3])^(a[105] & b[4])^(a[104] & b[5])^(a[103] & b[6])^(a[102] & b[7])^(a[101] & b[8])^(a[100] & b[9])^(a[99] & b[10])^(a[98] & b[11])^(a[97] & b[12])^(a[96] & b[13])^(a[95] & b[14])^(a[94] & b[15])^(a[93] & b[16])^(a[92] & b[17])^(a[91] & b[18])^(a[90] & b[19])^(a[89] & b[20])^(a[88] & b[21])^(a[87] & b[22])^(a[86] & b[23])^(a[85] & b[24])^(a[84] & b[25])^(a[83] & b[26])^(a[82] & b[27])^(a[81] & b[28])^(a[80] & b[29])^(a[79] & b[30])^(a[78] & b[31])^(a[77] & b[32])^(a[76] & b[33])^(a[75] & b[34])^(a[74] & b[35])^(a[73] & b[36])^(a[72] & b[37])^(a[71] & b[38])^(a[70] & b[39])^(a[69] & b[40])^(a[68] & b[41])^(a[67] & b[42])^(a[66] & b[43])^(a[65] & b[44])^(a[64] & b[45])^(a[63] & b[46])^(a[62] & b[47])^(a[61] & b[48])^(a[60] & b[49])^(a[59] & b[50])^(a[58] & b[51])^(a[57] & b[52])^(a[56] & b[53])^(a[55] & b[54])^(a[54] & b[55])^(a[53] & b[56])^(a[52] & b[57])^(a[51] & b[58])^(a[50] & b[59])^(a[49] & b[60])^(a[48] & b[61])^(a[47] & b[62])^(a[46] & b[63])^(a[45] & b[64])^(a[44] & b[65])^(a[43] & b[66])^(a[42] & b[67])^(a[41] & b[68])^(a[40] & b[69])^(a[39] & b[70])^(a[38] & b[71])^(a[37] & b[72])^(a[36] & b[73])^(a[35] & b[74])^(a[34] & b[75])^(a[33] & b[76])^(a[32] & b[77])^(a[31] & b[78])^(a[30] & b[79])^(a[29] & b[80])^(a[28] & b[81])^(a[27] & b[82])^(a[26] & b[83])^(a[25] & b[84])^(a[24] & b[85])^(a[23] & b[86])^(a[22] & b[87])^(a[21] & b[88])^(a[20] & b[89])^(a[19] & b[90])^(a[18] & b[91])^(a[17] & b[92])^(a[16] & b[93])^(a[15] & b[94])^(a[14] & b[95])^(a[13] & b[96])^(a[12] & b[97])^(a[11] & b[98])^(a[10] & b[99])^(a[9] & b[100])^(a[8] & b[101])^(a[7] & b[102])^(a[6] & b[103])^(a[5] & b[104])^(a[4] & b[105])^(a[3] & b[106])^(a[2] & b[107])^(a[1] & b[108])^(a[0] & b[109]);
assign y[110] = (a[110] & b[0])^(a[109] & b[1])^(a[108] & b[2])^(a[107] & b[3])^(a[106] & b[4])^(a[105] & b[5])^(a[104] & b[6])^(a[103] & b[7])^(a[102] & b[8])^(a[101] & b[9])^(a[100] & b[10])^(a[99] & b[11])^(a[98] & b[12])^(a[97] & b[13])^(a[96] & b[14])^(a[95] & b[15])^(a[94] & b[16])^(a[93] & b[17])^(a[92] & b[18])^(a[91] & b[19])^(a[90] & b[20])^(a[89] & b[21])^(a[88] & b[22])^(a[87] & b[23])^(a[86] & b[24])^(a[85] & b[25])^(a[84] & b[26])^(a[83] & b[27])^(a[82] & b[28])^(a[81] & b[29])^(a[80] & b[30])^(a[79] & b[31])^(a[78] & b[32])^(a[77] & b[33])^(a[76] & b[34])^(a[75] & b[35])^(a[74] & b[36])^(a[73] & b[37])^(a[72] & b[38])^(a[71] & b[39])^(a[70] & b[40])^(a[69] & b[41])^(a[68] & b[42])^(a[67] & b[43])^(a[66] & b[44])^(a[65] & b[45])^(a[64] & b[46])^(a[63] & b[47])^(a[62] & b[48])^(a[61] & b[49])^(a[60] & b[50])^(a[59] & b[51])^(a[58] & b[52])^(a[57] & b[53])^(a[56] & b[54])^(a[55] & b[55])^(a[54] & b[56])^(a[53] & b[57])^(a[52] & b[58])^(a[51] & b[59])^(a[50] & b[60])^(a[49] & b[61])^(a[48] & b[62])^(a[47] & b[63])^(a[46] & b[64])^(a[45] & b[65])^(a[44] & b[66])^(a[43] & b[67])^(a[42] & b[68])^(a[41] & b[69])^(a[40] & b[70])^(a[39] & b[71])^(a[38] & b[72])^(a[37] & b[73])^(a[36] & b[74])^(a[35] & b[75])^(a[34] & b[76])^(a[33] & b[77])^(a[32] & b[78])^(a[31] & b[79])^(a[30] & b[80])^(a[29] & b[81])^(a[28] & b[82])^(a[27] & b[83])^(a[26] & b[84])^(a[25] & b[85])^(a[24] & b[86])^(a[23] & b[87])^(a[22] & b[88])^(a[21] & b[89])^(a[20] & b[90])^(a[19] & b[91])^(a[18] & b[92])^(a[17] & b[93])^(a[16] & b[94])^(a[15] & b[95])^(a[14] & b[96])^(a[13] & b[97])^(a[12] & b[98])^(a[11] & b[99])^(a[10] & b[100])^(a[9] & b[101])^(a[8] & b[102])^(a[7] & b[103])^(a[6] & b[104])^(a[5] & b[105])^(a[4] & b[106])^(a[3] & b[107])^(a[2] & b[108])^(a[1] & b[109])^(a[0] & b[110]);
assign y[111] = (a[111] & b[0])^(a[110] & b[1])^(a[109] & b[2])^(a[108] & b[3])^(a[107] & b[4])^(a[106] & b[5])^(a[105] & b[6])^(a[104] & b[7])^(a[103] & b[8])^(a[102] & b[9])^(a[101] & b[10])^(a[100] & b[11])^(a[99] & b[12])^(a[98] & b[13])^(a[97] & b[14])^(a[96] & b[15])^(a[95] & b[16])^(a[94] & b[17])^(a[93] & b[18])^(a[92] & b[19])^(a[91] & b[20])^(a[90] & b[21])^(a[89] & b[22])^(a[88] & b[23])^(a[87] & b[24])^(a[86] & b[25])^(a[85] & b[26])^(a[84] & b[27])^(a[83] & b[28])^(a[82] & b[29])^(a[81] & b[30])^(a[80] & b[31])^(a[79] & b[32])^(a[78] & b[33])^(a[77] & b[34])^(a[76] & b[35])^(a[75] & b[36])^(a[74] & b[37])^(a[73] & b[38])^(a[72] & b[39])^(a[71] & b[40])^(a[70] & b[41])^(a[69] & b[42])^(a[68] & b[43])^(a[67] & b[44])^(a[66] & b[45])^(a[65] & b[46])^(a[64] & b[47])^(a[63] & b[48])^(a[62] & b[49])^(a[61] & b[50])^(a[60] & b[51])^(a[59] & b[52])^(a[58] & b[53])^(a[57] & b[54])^(a[56] & b[55])^(a[55] & b[56])^(a[54] & b[57])^(a[53] & b[58])^(a[52] & b[59])^(a[51] & b[60])^(a[50] & b[61])^(a[49] & b[62])^(a[48] & b[63])^(a[47] & b[64])^(a[46] & b[65])^(a[45] & b[66])^(a[44] & b[67])^(a[43] & b[68])^(a[42] & b[69])^(a[41] & b[70])^(a[40] & b[71])^(a[39] & b[72])^(a[38] & b[73])^(a[37] & b[74])^(a[36] & b[75])^(a[35] & b[76])^(a[34] & b[77])^(a[33] & b[78])^(a[32] & b[79])^(a[31] & b[80])^(a[30] & b[81])^(a[29] & b[82])^(a[28] & b[83])^(a[27] & b[84])^(a[26] & b[85])^(a[25] & b[86])^(a[24] & b[87])^(a[23] & b[88])^(a[22] & b[89])^(a[21] & b[90])^(a[20] & b[91])^(a[19] & b[92])^(a[18] & b[93])^(a[17] & b[94])^(a[16] & b[95])^(a[15] & b[96])^(a[14] & b[97])^(a[13] & b[98])^(a[12] & b[99])^(a[11] & b[100])^(a[10] & b[101])^(a[9] & b[102])^(a[8] & b[103])^(a[7] & b[104])^(a[6] & b[105])^(a[5] & b[106])^(a[4] & b[107])^(a[3] & b[108])^(a[2] & b[109])^(a[1] & b[110])^(a[0] & b[111]);
assign y[112] = (a[112] & b[0])^(a[111] & b[1])^(a[110] & b[2])^(a[109] & b[3])^(a[108] & b[4])^(a[107] & b[5])^(a[106] & b[6])^(a[105] & b[7])^(a[104] & b[8])^(a[103] & b[9])^(a[102] & b[10])^(a[101] & b[11])^(a[100] & b[12])^(a[99] & b[13])^(a[98] & b[14])^(a[97] & b[15])^(a[96] & b[16])^(a[95] & b[17])^(a[94] & b[18])^(a[93] & b[19])^(a[92] & b[20])^(a[91] & b[21])^(a[90] & b[22])^(a[89] & b[23])^(a[88] & b[24])^(a[87] & b[25])^(a[86] & b[26])^(a[85] & b[27])^(a[84] & b[28])^(a[83] & b[29])^(a[82] & b[30])^(a[81] & b[31])^(a[80] & b[32])^(a[79] & b[33])^(a[78] & b[34])^(a[77] & b[35])^(a[76] & b[36])^(a[75] & b[37])^(a[74] & b[38])^(a[73] & b[39])^(a[72] & b[40])^(a[71] & b[41])^(a[70] & b[42])^(a[69] & b[43])^(a[68] & b[44])^(a[67] & b[45])^(a[66] & b[46])^(a[65] & b[47])^(a[64] & b[48])^(a[63] & b[49])^(a[62] & b[50])^(a[61] & b[51])^(a[60] & b[52])^(a[59] & b[53])^(a[58] & b[54])^(a[57] & b[55])^(a[56] & b[56])^(a[55] & b[57])^(a[54] & b[58])^(a[53] & b[59])^(a[52] & b[60])^(a[51] & b[61])^(a[50] & b[62])^(a[49] & b[63])^(a[48] & b[64])^(a[47] & b[65])^(a[46] & b[66])^(a[45] & b[67])^(a[44] & b[68])^(a[43] & b[69])^(a[42] & b[70])^(a[41] & b[71])^(a[40] & b[72])^(a[39] & b[73])^(a[38] & b[74])^(a[37] & b[75])^(a[36] & b[76])^(a[35] & b[77])^(a[34] & b[78])^(a[33] & b[79])^(a[32] & b[80])^(a[31] & b[81])^(a[30] & b[82])^(a[29] & b[83])^(a[28] & b[84])^(a[27] & b[85])^(a[26] & b[86])^(a[25] & b[87])^(a[24] & b[88])^(a[23] & b[89])^(a[22] & b[90])^(a[21] & b[91])^(a[20] & b[92])^(a[19] & b[93])^(a[18] & b[94])^(a[17] & b[95])^(a[16] & b[96])^(a[15] & b[97])^(a[14] & b[98])^(a[13] & b[99])^(a[12] & b[100])^(a[11] & b[101])^(a[10] & b[102])^(a[9] & b[103])^(a[8] & b[104])^(a[7] & b[105])^(a[6] & b[106])^(a[5] & b[107])^(a[4] & b[108])^(a[3] & b[109])^(a[2] & b[110])^(a[1] & b[111])^(a[0] & b[112]);
assign y[113] = (a[113] & b[0])^(a[112] & b[1])^(a[111] & b[2])^(a[110] & b[3])^(a[109] & b[4])^(a[108] & b[5])^(a[107] & b[6])^(a[106] & b[7])^(a[105] & b[8])^(a[104] & b[9])^(a[103] & b[10])^(a[102] & b[11])^(a[101] & b[12])^(a[100] & b[13])^(a[99] & b[14])^(a[98] & b[15])^(a[97] & b[16])^(a[96] & b[17])^(a[95] & b[18])^(a[94] & b[19])^(a[93] & b[20])^(a[92] & b[21])^(a[91] & b[22])^(a[90] & b[23])^(a[89] & b[24])^(a[88] & b[25])^(a[87] & b[26])^(a[86] & b[27])^(a[85] & b[28])^(a[84] & b[29])^(a[83] & b[30])^(a[82] & b[31])^(a[81] & b[32])^(a[80] & b[33])^(a[79] & b[34])^(a[78] & b[35])^(a[77] & b[36])^(a[76] & b[37])^(a[75] & b[38])^(a[74] & b[39])^(a[73] & b[40])^(a[72] & b[41])^(a[71] & b[42])^(a[70] & b[43])^(a[69] & b[44])^(a[68] & b[45])^(a[67] & b[46])^(a[66] & b[47])^(a[65] & b[48])^(a[64] & b[49])^(a[63] & b[50])^(a[62] & b[51])^(a[61] & b[52])^(a[60] & b[53])^(a[59] & b[54])^(a[58] & b[55])^(a[57] & b[56])^(a[56] & b[57])^(a[55] & b[58])^(a[54] & b[59])^(a[53] & b[60])^(a[52] & b[61])^(a[51] & b[62])^(a[50] & b[63])^(a[49] & b[64])^(a[48] & b[65])^(a[47] & b[66])^(a[46] & b[67])^(a[45] & b[68])^(a[44] & b[69])^(a[43] & b[70])^(a[42] & b[71])^(a[41] & b[72])^(a[40] & b[73])^(a[39] & b[74])^(a[38] & b[75])^(a[37] & b[76])^(a[36] & b[77])^(a[35] & b[78])^(a[34] & b[79])^(a[33] & b[80])^(a[32] & b[81])^(a[31] & b[82])^(a[30] & b[83])^(a[29] & b[84])^(a[28] & b[85])^(a[27] & b[86])^(a[26] & b[87])^(a[25] & b[88])^(a[24] & b[89])^(a[23] & b[90])^(a[22] & b[91])^(a[21] & b[92])^(a[20] & b[93])^(a[19] & b[94])^(a[18] & b[95])^(a[17] & b[96])^(a[16] & b[97])^(a[15] & b[98])^(a[14] & b[99])^(a[13] & b[100])^(a[12] & b[101])^(a[11] & b[102])^(a[10] & b[103])^(a[9] & b[104])^(a[8] & b[105])^(a[7] & b[106])^(a[6] & b[107])^(a[5] & b[108])^(a[4] & b[109])^(a[3] & b[110])^(a[2] & b[111])^(a[1] & b[112])^(a[0] & b[113]);
assign y[114] = (a[114] & b[0])^(a[113] & b[1])^(a[112] & b[2])^(a[111] & b[3])^(a[110] & b[4])^(a[109] & b[5])^(a[108] & b[6])^(a[107] & b[7])^(a[106] & b[8])^(a[105] & b[9])^(a[104] & b[10])^(a[103] & b[11])^(a[102] & b[12])^(a[101] & b[13])^(a[100] & b[14])^(a[99] & b[15])^(a[98] & b[16])^(a[97] & b[17])^(a[96] & b[18])^(a[95] & b[19])^(a[94] & b[20])^(a[93] & b[21])^(a[92] & b[22])^(a[91] & b[23])^(a[90] & b[24])^(a[89] & b[25])^(a[88] & b[26])^(a[87] & b[27])^(a[86] & b[28])^(a[85] & b[29])^(a[84] & b[30])^(a[83] & b[31])^(a[82] & b[32])^(a[81] & b[33])^(a[80] & b[34])^(a[79] & b[35])^(a[78] & b[36])^(a[77] & b[37])^(a[76] & b[38])^(a[75] & b[39])^(a[74] & b[40])^(a[73] & b[41])^(a[72] & b[42])^(a[71] & b[43])^(a[70] & b[44])^(a[69] & b[45])^(a[68] & b[46])^(a[67] & b[47])^(a[66] & b[48])^(a[65] & b[49])^(a[64] & b[50])^(a[63] & b[51])^(a[62] & b[52])^(a[61] & b[53])^(a[60] & b[54])^(a[59] & b[55])^(a[58] & b[56])^(a[57] & b[57])^(a[56] & b[58])^(a[55] & b[59])^(a[54] & b[60])^(a[53] & b[61])^(a[52] & b[62])^(a[51] & b[63])^(a[50] & b[64])^(a[49] & b[65])^(a[48] & b[66])^(a[47] & b[67])^(a[46] & b[68])^(a[45] & b[69])^(a[44] & b[70])^(a[43] & b[71])^(a[42] & b[72])^(a[41] & b[73])^(a[40] & b[74])^(a[39] & b[75])^(a[38] & b[76])^(a[37] & b[77])^(a[36] & b[78])^(a[35] & b[79])^(a[34] & b[80])^(a[33] & b[81])^(a[32] & b[82])^(a[31] & b[83])^(a[30] & b[84])^(a[29] & b[85])^(a[28] & b[86])^(a[27] & b[87])^(a[26] & b[88])^(a[25] & b[89])^(a[24] & b[90])^(a[23] & b[91])^(a[22] & b[92])^(a[21] & b[93])^(a[20] & b[94])^(a[19] & b[95])^(a[18] & b[96])^(a[17] & b[97])^(a[16] & b[98])^(a[15] & b[99])^(a[14] & b[100])^(a[13] & b[101])^(a[12] & b[102])^(a[11] & b[103])^(a[10] & b[104])^(a[9] & b[105])^(a[8] & b[106])^(a[7] & b[107])^(a[6] & b[108])^(a[5] & b[109])^(a[4] & b[110])^(a[3] & b[111])^(a[2] & b[112])^(a[1] & b[113])^(a[0] & b[114]);
assign y[115] = (a[115] & b[0])^(a[114] & b[1])^(a[113] & b[2])^(a[112] & b[3])^(a[111] & b[4])^(a[110] & b[5])^(a[109] & b[6])^(a[108] & b[7])^(a[107] & b[8])^(a[106] & b[9])^(a[105] & b[10])^(a[104] & b[11])^(a[103] & b[12])^(a[102] & b[13])^(a[101] & b[14])^(a[100] & b[15])^(a[99] & b[16])^(a[98] & b[17])^(a[97] & b[18])^(a[96] & b[19])^(a[95] & b[20])^(a[94] & b[21])^(a[93] & b[22])^(a[92] & b[23])^(a[91] & b[24])^(a[90] & b[25])^(a[89] & b[26])^(a[88] & b[27])^(a[87] & b[28])^(a[86] & b[29])^(a[85] & b[30])^(a[84] & b[31])^(a[83] & b[32])^(a[82] & b[33])^(a[81] & b[34])^(a[80] & b[35])^(a[79] & b[36])^(a[78] & b[37])^(a[77] & b[38])^(a[76] & b[39])^(a[75] & b[40])^(a[74] & b[41])^(a[73] & b[42])^(a[72] & b[43])^(a[71] & b[44])^(a[70] & b[45])^(a[69] & b[46])^(a[68] & b[47])^(a[67] & b[48])^(a[66] & b[49])^(a[65] & b[50])^(a[64] & b[51])^(a[63] & b[52])^(a[62] & b[53])^(a[61] & b[54])^(a[60] & b[55])^(a[59] & b[56])^(a[58] & b[57])^(a[57] & b[58])^(a[56] & b[59])^(a[55] & b[60])^(a[54] & b[61])^(a[53] & b[62])^(a[52] & b[63])^(a[51] & b[64])^(a[50] & b[65])^(a[49] & b[66])^(a[48] & b[67])^(a[47] & b[68])^(a[46] & b[69])^(a[45] & b[70])^(a[44] & b[71])^(a[43] & b[72])^(a[42] & b[73])^(a[41] & b[74])^(a[40] & b[75])^(a[39] & b[76])^(a[38] & b[77])^(a[37] & b[78])^(a[36] & b[79])^(a[35] & b[80])^(a[34] & b[81])^(a[33] & b[82])^(a[32] & b[83])^(a[31] & b[84])^(a[30] & b[85])^(a[29] & b[86])^(a[28] & b[87])^(a[27] & b[88])^(a[26] & b[89])^(a[25] & b[90])^(a[24] & b[91])^(a[23] & b[92])^(a[22] & b[93])^(a[21] & b[94])^(a[20] & b[95])^(a[19] & b[96])^(a[18] & b[97])^(a[17] & b[98])^(a[16] & b[99])^(a[15] & b[100])^(a[14] & b[101])^(a[13] & b[102])^(a[12] & b[103])^(a[11] & b[104])^(a[10] & b[105])^(a[9] & b[106])^(a[8] & b[107])^(a[7] & b[108])^(a[6] & b[109])^(a[5] & b[110])^(a[4] & b[111])^(a[3] & b[112])^(a[2] & b[113])^(a[1] & b[114])^(a[0] & b[115]);
assign y[116] = (a[116] & b[0])^(a[115] & b[1])^(a[114] & b[2])^(a[113] & b[3])^(a[112] & b[4])^(a[111] & b[5])^(a[110] & b[6])^(a[109] & b[7])^(a[108] & b[8])^(a[107] & b[9])^(a[106] & b[10])^(a[105] & b[11])^(a[104] & b[12])^(a[103] & b[13])^(a[102] & b[14])^(a[101] & b[15])^(a[100] & b[16])^(a[99] & b[17])^(a[98] & b[18])^(a[97] & b[19])^(a[96] & b[20])^(a[95] & b[21])^(a[94] & b[22])^(a[93] & b[23])^(a[92] & b[24])^(a[91] & b[25])^(a[90] & b[26])^(a[89] & b[27])^(a[88] & b[28])^(a[87] & b[29])^(a[86] & b[30])^(a[85] & b[31])^(a[84] & b[32])^(a[83] & b[33])^(a[82] & b[34])^(a[81] & b[35])^(a[80] & b[36])^(a[79] & b[37])^(a[78] & b[38])^(a[77] & b[39])^(a[76] & b[40])^(a[75] & b[41])^(a[74] & b[42])^(a[73] & b[43])^(a[72] & b[44])^(a[71] & b[45])^(a[70] & b[46])^(a[69] & b[47])^(a[68] & b[48])^(a[67] & b[49])^(a[66] & b[50])^(a[65] & b[51])^(a[64] & b[52])^(a[63] & b[53])^(a[62] & b[54])^(a[61] & b[55])^(a[60] & b[56])^(a[59] & b[57])^(a[58] & b[58])^(a[57] & b[59])^(a[56] & b[60])^(a[55] & b[61])^(a[54] & b[62])^(a[53] & b[63])^(a[52] & b[64])^(a[51] & b[65])^(a[50] & b[66])^(a[49] & b[67])^(a[48] & b[68])^(a[47] & b[69])^(a[46] & b[70])^(a[45] & b[71])^(a[44] & b[72])^(a[43] & b[73])^(a[42] & b[74])^(a[41] & b[75])^(a[40] & b[76])^(a[39] & b[77])^(a[38] & b[78])^(a[37] & b[79])^(a[36] & b[80])^(a[35] & b[81])^(a[34] & b[82])^(a[33] & b[83])^(a[32] & b[84])^(a[31] & b[85])^(a[30] & b[86])^(a[29] & b[87])^(a[28] & b[88])^(a[27] & b[89])^(a[26] & b[90])^(a[25] & b[91])^(a[24] & b[92])^(a[23] & b[93])^(a[22] & b[94])^(a[21] & b[95])^(a[20] & b[96])^(a[19] & b[97])^(a[18] & b[98])^(a[17] & b[99])^(a[16] & b[100])^(a[15] & b[101])^(a[14] & b[102])^(a[13] & b[103])^(a[12] & b[104])^(a[11] & b[105])^(a[10] & b[106])^(a[9] & b[107])^(a[8] & b[108])^(a[7] & b[109])^(a[6] & b[110])^(a[5] & b[111])^(a[4] & b[112])^(a[3] & b[113])^(a[2] & b[114])^(a[1] & b[115])^(a[0] & b[116]);
assign y[117] = (a[117] & b[0])^(a[116] & b[1])^(a[115] & b[2])^(a[114] & b[3])^(a[113] & b[4])^(a[112] & b[5])^(a[111] & b[6])^(a[110] & b[7])^(a[109] & b[8])^(a[108] & b[9])^(a[107] & b[10])^(a[106] & b[11])^(a[105] & b[12])^(a[104] & b[13])^(a[103] & b[14])^(a[102] & b[15])^(a[101] & b[16])^(a[100] & b[17])^(a[99] & b[18])^(a[98] & b[19])^(a[97] & b[20])^(a[96] & b[21])^(a[95] & b[22])^(a[94] & b[23])^(a[93] & b[24])^(a[92] & b[25])^(a[91] & b[26])^(a[90] & b[27])^(a[89] & b[28])^(a[88] & b[29])^(a[87] & b[30])^(a[86] & b[31])^(a[85] & b[32])^(a[84] & b[33])^(a[83] & b[34])^(a[82] & b[35])^(a[81] & b[36])^(a[80] & b[37])^(a[79] & b[38])^(a[78] & b[39])^(a[77] & b[40])^(a[76] & b[41])^(a[75] & b[42])^(a[74] & b[43])^(a[73] & b[44])^(a[72] & b[45])^(a[71] & b[46])^(a[70] & b[47])^(a[69] & b[48])^(a[68] & b[49])^(a[67] & b[50])^(a[66] & b[51])^(a[65] & b[52])^(a[64] & b[53])^(a[63] & b[54])^(a[62] & b[55])^(a[61] & b[56])^(a[60] & b[57])^(a[59] & b[58])^(a[58] & b[59])^(a[57] & b[60])^(a[56] & b[61])^(a[55] & b[62])^(a[54] & b[63])^(a[53] & b[64])^(a[52] & b[65])^(a[51] & b[66])^(a[50] & b[67])^(a[49] & b[68])^(a[48] & b[69])^(a[47] & b[70])^(a[46] & b[71])^(a[45] & b[72])^(a[44] & b[73])^(a[43] & b[74])^(a[42] & b[75])^(a[41] & b[76])^(a[40] & b[77])^(a[39] & b[78])^(a[38] & b[79])^(a[37] & b[80])^(a[36] & b[81])^(a[35] & b[82])^(a[34] & b[83])^(a[33] & b[84])^(a[32] & b[85])^(a[31] & b[86])^(a[30] & b[87])^(a[29] & b[88])^(a[28] & b[89])^(a[27] & b[90])^(a[26] & b[91])^(a[25] & b[92])^(a[24] & b[93])^(a[23] & b[94])^(a[22] & b[95])^(a[21] & b[96])^(a[20] & b[97])^(a[19] & b[98])^(a[18] & b[99])^(a[17] & b[100])^(a[16] & b[101])^(a[15] & b[102])^(a[14] & b[103])^(a[13] & b[104])^(a[12] & b[105])^(a[11] & b[106])^(a[10] & b[107])^(a[9] & b[108])^(a[8] & b[109])^(a[7] & b[110])^(a[6] & b[111])^(a[5] & b[112])^(a[4] & b[113])^(a[3] & b[114])^(a[2] & b[115])^(a[1] & b[116])^(a[0] & b[117]);
assign y[118] = (a[118] & b[0])^(a[117] & b[1])^(a[116] & b[2])^(a[115] & b[3])^(a[114] & b[4])^(a[113] & b[5])^(a[112] & b[6])^(a[111] & b[7])^(a[110] & b[8])^(a[109] & b[9])^(a[108] & b[10])^(a[107] & b[11])^(a[106] & b[12])^(a[105] & b[13])^(a[104] & b[14])^(a[103] & b[15])^(a[102] & b[16])^(a[101] & b[17])^(a[100] & b[18])^(a[99] & b[19])^(a[98] & b[20])^(a[97] & b[21])^(a[96] & b[22])^(a[95] & b[23])^(a[94] & b[24])^(a[93] & b[25])^(a[92] & b[26])^(a[91] & b[27])^(a[90] & b[28])^(a[89] & b[29])^(a[88] & b[30])^(a[87] & b[31])^(a[86] & b[32])^(a[85] & b[33])^(a[84] & b[34])^(a[83] & b[35])^(a[82] & b[36])^(a[81] & b[37])^(a[80] & b[38])^(a[79] & b[39])^(a[78] & b[40])^(a[77] & b[41])^(a[76] & b[42])^(a[75] & b[43])^(a[74] & b[44])^(a[73] & b[45])^(a[72] & b[46])^(a[71] & b[47])^(a[70] & b[48])^(a[69] & b[49])^(a[68] & b[50])^(a[67] & b[51])^(a[66] & b[52])^(a[65] & b[53])^(a[64] & b[54])^(a[63] & b[55])^(a[62] & b[56])^(a[61] & b[57])^(a[60] & b[58])^(a[59] & b[59])^(a[58] & b[60])^(a[57] & b[61])^(a[56] & b[62])^(a[55] & b[63])^(a[54] & b[64])^(a[53] & b[65])^(a[52] & b[66])^(a[51] & b[67])^(a[50] & b[68])^(a[49] & b[69])^(a[48] & b[70])^(a[47] & b[71])^(a[46] & b[72])^(a[45] & b[73])^(a[44] & b[74])^(a[43] & b[75])^(a[42] & b[76])^(a[41] & b[77])^(a[40] & b[78])^(a[39] & b[79])^(a[38] & b[80])^(a[37] & b[81])^(a[36] & b[82])^(a[35] & b[83])^(a[34] & b[84])^(a[33] & b[85])^(a[32] & b[86])^(a[31] & b[87])^(a[30] & b[88])^(a[29] & b[89])^(a[28] & b[90])^(a[27] & b[91])^(a[26] & b[92])^(a[25] & b[93])^(a[24] & b[94])^(a[23] & b[95])^(a[22] & b[96])^(a[21] & b[97])^(a[20] & b[98])^(a[19] & b[99])^(a[18] & b[100])^(a[17] & b[101])^(a[16] & b[102])^(a[15] & b[103])^(a[14] & b[104])^(a[13] & b[105])^(a[12] & b[106])^(a[11] & b[107])^(a[10] & b[108])^(a[9] & b[109])^(a[8] & b[110])^(a[7] & b[111])^(a[6] & b[112])^(a[5] & b[113])^(a[4] & b[114])^(a[3] & b[115])^(a[2] & b[116])^(a[1] & b[117])^(a[0] & b[118]);
assign y[119] = (a[119] & b[0])^(a[118] & b[1])^(a[117] & b[2])^(a[116] & b[3])^(a[115] & b[4])^(a[114] & b[5])^(a[113] & b[6])^(a[112] & b[7])^(a[111] & b[8])^(a[110] & b[9])^(a[109] & b[10])^(a[108] & b[11])^(a[107] & b[12])^(a[106] & b[13])^(a[105] & b[14])^(a[104] & b[15])^(a[103] & b[16])^(a[102] & b[17])^(a[101] & b[18])^(a[100] & b[19])^(a[99] & b[20])^(a[98] & b[21])^(a[97] & b[22])^(a[96] & b[23])^(a[95] & b[24])^(a[94] & b[25])^(a[93] & b[26])^(a[92] & b[27])^(a[91] & b[28])^(a[90] & b[29])^(a[89] & b[30])^(a[88] & b[31])^(a[87] & b[32])^(a[86] & b[33])^(a[85] & b[34])^(a[84] & b[35])^(a[83] & b[36])^(a[82] & b[37])^(a[81] & b[38])^(a[80] & b[39])^(a[79] & b[40])^(a[78] & b[41])^(a[77] & b[42])^(a[76] & b[43])^(a[75] & b[44])^(a[74] & b[45])^(a[73] & b[46])^(a[72] & b[47])^(a[71] & b[48])^(a[70] & b[49])^(a[69] & b[50])^(a[68] & b[51])^(a[67] & b[52])^(a[66] & b[53])^(a[65] & b[54])^(a[64] & b[55])^(a[63] & b[56])^(a[62] & b[57])^(a[61] & b[58])^(a[60] & b[59])^(a[59] & b[60])^(a[58] & b[61])^(a[57] & b[62])^(a[56] & b[63])^(a[55] & b[64])^(a[54] & b[65])^(a[53] & b[66])^(a[52] & b[67])^(a[51] & b[68])^(a[50] & b[69])^(a[49] & b[70])^(a[48] & b[71])^(a[47] & b[72])^(a[46] & b[73])^(a[45] & b[74])^(a[44] & b[75])^(a[43] & b[76])^(a[42] & b[77])^(a[41] & b[78])^(a[40] & b[79])^(a[39] & b[80])^(a[38] & b[81])^(a[37] & b[82])^(a[36] & b[83])^(a[35] & b[84])^(a[34] & b[85])^(a[33] & b[86])^(a[32] & b[87])^(a[31] & b[88])^(a[30] & b[89])^(a[29] & b[90])^(a[28] & b[91])^(a[27] & b[92])^(a[26] & b[93])^(a[25] & b[94])^(a[24] & b[95])^(a[23] & b[96])^(a[22] & b[97])^(a[21] & b[98])^(a[20] & b[99])^(a[19] & b[100])^(a[18] & b[101])^(a[17] & b[102])^(a[16] & b[103])^(a[15] & b[104])^(a[14] & b[105])^(a[13] & b[106])^(a[12] & b[107])^(a[11] & b[108])^(a[10] & b[109])^(a[9] & b[110])^(a[8] & b[111])^(a[7] & b[112])^(a[6] & b[113])^(a[5] & b[114])^(a[4] & b[115])^(a[3] & b[116])^(a[2] & b[117])^(a[1] & b[118])^(a[0] & b[119]);
assign y[120] = (a[120] & b[0])^(a[119] & b[1])^(a[118] & b[2])^(a[117] & b[3])^(a[116] & b[4])^(a[115] & b[5])^(a[114] & b[6])^(a[113] & b[7])^(a[112] & b[8])^(a[111] & b[9])^(a[110] & b[10])^(a[109] & b[11])^(a[108] & b[12])^(a[107] & b[13])^(a[106] & b[14])^(a[105] & b[15])^(a[104] & b[16])^(a[103] & b[17])^(a[102] & b[18])^(a[101] & b[19])^(a[100] & b[20])^(a[99] & b[21])^(a[98] & b[22])^(a[97] & b[23])^(a[96] & b[24])^(a[95] & b[25])^(a[94] & b[26])^(a[93] & b[27])^(a[92] & b[28])^(a[91] & b[29])^(a[90] & b[30])^(a[89] & b[31])^(a[88] & b[32])^(a[87] & b[33])^(a[86] & b[34])^(a[85] & b[35])^(a[84] & b[36])^(a[83] & b[37])^(a[82] & b[38])^(a[81] & b[39])^(a[80] & b[40])^(a[79] & b[41])^(a[78] & b[42])^(a[77] & b[43])^(a[76] & b[44])^(a[75] & b[45])^(a[74] & b[46])^(a[73] & b[47])^(a[72] & b[48])^(a[71] & b[49])^(a[70] & b[50])^(a[69] & b[51])^(a[68] & b[52])^(a[67] & b[53])^(a[66] & b[54])^(a[65] & b[55])^(a[64] & b[56])^(a[63] & b[57])^(a[62] & b[58])^(a[61] & b[59])^(a[60] & b[60])^(a[59] & b[61])^(a[58] & b[62])^(a[57] & b[63])^(a[56] & b[64])^(a[55] & b[65])^(a[54] & b[66])^(a[53] & b[67])^(a[52] & b[68])^(a[51] & b[69])^(a[50] & b[70])^(a[49] & b[71])^(a[48] & b[72])^(a[47] & b[73])^(a[46] & b[74])^(a[45] & b[75])^(a[44] & b[76])^(a[43] & b[77])^(a[42] & b[78])^(a[41] & b[79])^(a[40] & b[80])^(a[39] & b[81])^(a[38] & b[82])^(a[37] & b[83])^(a[36] & b[84])^(a[35] & b[85])^(a[34] & b[86])^(a[33] & b[87])^(a[32] & b[88])^(a[31] & b[89])^(a[30] & b[90])^(a[29] & b[91])^(a[28] & b[92])^(a[27] & b[93])^(a[26] & b[94])^(a[25] & b[95])^(a[24] & b[96])^(a[23] & b[97])^(a[22] & b[98])^(a[21] & b[99])^(a[20] & b[100])^(a[19] & b[101])^(a[18] & b[102])^(a[17] & b[103])^(a[16] & b[104])^(a[15] & b[105])^(a[14] & b[106])^(a[13] & b[107])^(a[12] & b[108])^(a[11] & b[109])^(a[10] & b[110])^(a[9] & b[111])^(a[8] & b[112])^(a[7] & b[113])^(a[6] & b[114])^(a[5] & b[115])^(a[4] & b[116])^(a[3] & b[117])^(a[2] & b[118])^(a[1] & b[119])^(a[0] & b[120]);
assign y[121] = (a[121] & b[0])^(a[120] & b[1])^(a[119] & b[2])^(a[118] & b[3])^(a[117] & b[4])^(a[116] & b[5])^(a[115] & b[6])^(a[114] & b[7])^(a[113] & b[8])^(a[112] & b[9])^(a[111] & b[10])^(a[110] & b[11])^(a[109] & b[12])^(a[108] & b[13])^(a[107] & b[14])^(a[106] & b[15])^(a[105] & b[16])^(a[104] & b[17])^(a[103] & b[18])^(a[102] & b[19])^(a[101] & b[20])^(a[100] & b[21])^(a[99] & b[22])^(a[98] & b[23])^(a[97] & b[24])^(a[96] & b[25])^(a[95] & b[26])^(a[94] & b[27])^(a[93] & b[28])^(a[92] & b[29])^(a[91] & b[30])^(a[90] & b[31])^(a[89] & b[32])^(a[88] & b[33])^(a[87] & b[34])^(a[86] & b[35])^(a[85] & b[36])^(a[84] & b[37])^(a[83] & b[38])^(a[82] & b[39])^(a[81] & b[40])^(a[80] & b[41])^(a[79] & b[42])^(a[78] & b[43])^(a[77] & b[44])^(a[76] & b[45])^(a[75] & b[46])^(a[74] & b[47])^(a[73] & b[48])^(a[72] & b[49])^(a[71] & b[50])^(a[70] & b[51])^(a[69] & b[52])^(a[68] & b[53])^(a[67] & b[54])^(a[66] & b[55])^(a[65] & b[56])^(a[64] & b[57])^(a[63] & b[58])^(a[62] & b[59])^(a[61] & b[60])^(a[60] & b[61])^(a[59] & b[62])^(a[58] & b[63])^(a[57] & b[64])^(a[56] & b[65])^(a[55] & b[66])^(a[54] & b[67])^(a[53] & b[68])^(a[52] & b[69])^(a[51] & b[70])^(a[50] & b[71])^(a[49] & b[72])^(a[48] & b[73])^(a[47] & b[74])^(a[46] & b[75])^(a[45] & b[76])^(a[44] & b[77])^(a[43] & b[78])^(a[42] & b[79])^(a[41] & b[80])^(a[40] & b[81])^(a[39] & b[82])^(a[38] & b[83])^(a[37] & b[84])^(a[36] & b[85])^(a[35] & b[86])^(a[34] & b[87])^(a[33] & b[88])^(a[32] & b[89])^(a[31] & b[90])^(a[30] & b[91])^(a[29] & b[92])^(a[28] & b[93])^(a[27] & b[94])^(a[26] & b[95])^(a[25] & b[96])^(a[24] & b[97])^(a[23] & b[98])^(a[22] & b[99])^(a[21] & b[100])^(a[20] & b[101])^(a[19] & b[102])^(a[18] & b[103])^(a[17] & b[104])^(a[16] & b[105])^(a[15] & b[106])^(a[14] & b[107])^(a[13] & b[108])^(a[12] & b[109])^(a[11] & b[110])^(a[10] & b[111])^(a[9] & b[112])^(a[8] & b[113])^(a[7] & b[114])^(a[6] & b[115])^(a[5] & b[116])^(a[4] & b[117])^(a[3] & b[118])^(a[2] & b[119])^(a[1] & b[120])^(a[0] & b[121]);
assign y[122] = (a[122] & b[0])^(a[121] & b[1])^(a[120] & b[2])^(a[119] & b[3])^(a[118] & b[4])^(a[117] & b[5])^(a[116] & b[6])^(a[115] & b[7])^(a[114] & b[8])^(a[113] & b[9])^(a[112] & b[10])^(a[111] & b[11])^(a[110] & b[12])^(a[109] & b[13])^(a[108] & b[14])^(a[107] & b[15])^(a[106] & b[16])^(a[105] & b[17])^(a[104] & b[18])^(a[103] & b[19])^(a[102] & b[20])^(a[101] & b[21])^(a[100] & b[22])^(a[99] & b[23])^(a[98] & b[24])^(a[97] & b[25])^(a[96] & b[26])^(a[95] & b[27])^(a[94] & b[28])^(a[93] & b[29])^(a[92] & b[30])^(a[91] & b[31])^(a[90] & b[32])^(a[89] & b[33])^(a[88] & b[34])^(a[87] & b[35])^(a[86] & b[36])^(a[85] & b[37])^(a[84] & b[38])^(a[83] & b[39])^(a[82] & b[40])^(a[81] & b[41])^(a[80] & b[42])^(a[79] & b[43])^(a[78] & b[44])^(a[77] & b[45])^(a[76] & b[46])^(a[75] & b[47])^(a[74] & b[48])^(a[73] & b[49])^(a[72] & b[50])^(a[71] & b[51])^(a[70] & b[52])^(a[69] & b[53])^(a[68] & b[54])^(a[67] & b[55])^(a[66] & b[56])^(a[65] & b[57])^(a[64] & b[58])^(a[63] & b[59])^(a[62] & b[60])^(a[61] & b[61])^(a[60] & b[62])^(a[59] & b[63])^(a[58] & b[64])^(a[57] & b[65])^(a[56] & b[66])^(a[55] & b[67])^(a[54] & b[68])^(a[53] & b[69])^(a[52] & b[70])^(a[51] & b[71])^(a[50] & b[72])^(a[49] & b[73])^(a[48] & b[74])^(a[47] & b[75])^(a[46] & b[76])^(a[45] & b[77])^(a[44] & b[78])^(a[43] & b[79])^(a[42] & b[80])^(a[41] & b[81])^(a[40] & b[82])^(a[39] & b[83])^(a[38] & b[84])^(a[37] & b[85])^(a[36] & b[86])^(a[35] & b[87])^(a[34] & b[88])^(a[33] & b[89])^(a[32] & b[90])^(a[31] & b[91])^(a[30] & b[92])^(a[29] & b[93])^(a[28] & b[94])^(a[27] & b[95])^(a[26] & b[96])^(a[25] & b[97])^(a[24] & b[98])^(a[23] & b[99])^(a[22] & b[100])^(a[21] & b[101])^(a[20] & b[102])^(a[19] & b[103])^(a[18] & b[104])^(a[17] & b[105])^(a[16] & b[106])^(a[15] & b[107])^(a[14] & b[108])^(a[13] & b[109])^(a[12] & b[110])^(a[11] & b[111])^(a[10] & b[112])^(a[9] & b[113])^(a[8] & b[114])^(a[7] & b[115])^(a[6] & b[116])^(a[5] & b[117])^(a[4] & b[118])^(a[3] & b[119])^(a[2] & b[120])^(a[1] & b[121])^(a[0] & b[122]);
assign y[123] = (a[123] & b[0])^(a[122] & b[1])^(a[121] & b[2])^(a[120] & b[3])^(a[119] & b[4])^(a[118] & b[5])^(a[117] & b[6])^(a[116] & b[7])^(a[115] & b[8])^(a[114] & b[9])^(a[113] & b[10])^(a[112] & b[11])^(a[111] & b[12])^(a[110] & b[13])^(a[109] & b[14])^(a[108] & b[15])^(a[107] & b[16])^(a[106] & b[17])^(a[105] & b[18])^(a[104] & b[19])^(a[103] & b[20])^(a[102] & b[21])^(a[101] & b[22])^(a[100] & b[23])^(a[99] & b[24])^(a[98] & b[25])^(a[97] & b[26])^(a[96] & b[27])^(a[95] & b[28])^(a[94] & b[29])^(a[93] & b[30])^(a[92] & b[31])^(a[91] & b[32])^(a[90] & b[33])^(a[89] & b[34])^(a[88] & b[35])^(a[87] & b[36])^(a[86] & b[37])^(a[85] & b[38])^(a[84] & b[39])^(a[83] & b[40])^(a[82] & b[41])^(a[81] & b[42])^(a[80] & b[43])^(a[79] & b[44])^(a[78] & b[45])^(a[77] & b[46])^(a[76] & b[47])^(a[75] & b[48])^(a[74] & b[49])^(a[73] & b[50])^(a[72] & b[51])^(a[71] & b[52])^(a[70] & b[53])^(a[69] & b[54])^(a[68] & b[55])^(a[67] & b[56])^(a[66] & b[57])^(a[65] & b[58])^(a[64] & b[59])^(a[63] & b[60])^(a[62] & b[61])^(a[61] & b[62])^(a[60] & b[63])^(a[59] & b[64])^(a[58] & b[65])^(a[57] & b[66])^(a[56] & b[67])^(a[55] & b[68])^(a[54] & b[69])^(a[53] & b[70])^(a[52] & b[71])^(a[51] & b[72])^(a[50] & b[73])^(a[49] & b[74])^(a[48] & b[75])^(a[47] & b[76])^(a[46] & b[77])^(a[45] & b[78])^(a[44] & b[79])^(a[43] & b[80])^(a[42] & b[81])^(a[41] & b[82])^(a[40] & b[83])^(a[39] & b[84])^(a[38] & b[85])^(a[37] & b[86])^(a[36] & b[87])^(a[35] & b[88])^(a[34] & b[89])^(a[33] & b[90])^(a[32] & b[91])^(a[31] & b[92])^(a[30] & b[93])^(a[29] & b[94])^(a[28] & b[95])^(a[27] & b[96])^(a[26] & b[97])^(a[25] & b[98])^(a[24] & b[99])^(a[23] & b[100])^(a[22] & b[101])^(a[21] & b[102])^(a[20] & b[103])^(a[19] & b[104])^(a[18] & b[105])^(a[17] & b[106])^(a[16] & b[107])^(a[15] & b[108])^(a[14] & b[109])^(a[13] & b[110])^(a[12] & b[111])^(a[11] & b[112])^(a[10] & b[113])^(a[9] & b[114])^(a[8] & b[115])^(a[7] & b[116])^(a[6] & b[117])^(a[5] & b[118])^(a[4] & b[119])^(a[3] & b[120])^(a[2] & b[121])^(a[1] & b[122])^(a[0] & b[123]);
assign y[124] = (a[124] & b[0])^(a[123] & b[1])^(a[122] & b[2])^(a[121] & b[3])^(a[120] & b[4])^(a[119] & b[5])^(a[118] & b[6])^(a[117] & b[7])^(a[116] & b[8])^(a[115] & b[9])^(a[114] & b[10])^(a[113] & b[11])^(a[112] & b[12])^(a[111] & b[13])^(a[110] & b[14])^(a[109] & b[15])^(a[108] & b[16])^(a[107] & b[17])^(a[106] & b[18])^(a[105] & b[19])^(a[104] & b[20])^(a[103] & b[21])^(a[102] & b[22])^(a[101] & b[23])^(a[100] & b[24])^(a[99] & b[25])^(a[98] & b[26])^(a[97] & b[27])^(a[96] & b[28])^(a[95] & b[29])^(a[94] & b[30])^(a[93] & b[31])^(a[92] & b[32])^(a[91] & b[33])^(a[90] & b[34])^(a[89] & b[35])^(a[88] & b[36])^(a[87] & b[37])^(a[86] & b[38])^(a[85] & b[39])^(a[84] & b[40])^(a[83] & b[41])^(a[82] & b[42])^(a[81] & b[43])^(a[80] & b[44])^(a[79] & b[45])^(a[78] & b[46])^(a[77] & b[47])^(a[76] & b[48])^(a[75] & b[49])^(a[74] & b[50])^(a[73] & b[51])^(a[72] & b[52])^(a[71] & b[53])^(a[70] & b[54])^(a[69] & b[55])^(a[68] & b[56])^(a[67] & b[57])^(a[66] & b[58])^(a[65] & b[59])^(a[64] & b[60])^(a[63] & b[61])^(a[62] & b[62])^(a[61] & b[63])^(a[60] & b[64])^(a[59] & b[65])^(a[58] & b[66])^(a[57] & b[67])^(a[56] & b[68])^(a[55] & b[69])^(a[54] & b[70])^(a[53] & b[71])^(a[52] & b[72])^(a[51] & b[73])^(a[50] & b[74])^(a[49] & b[75])^(a[48] & b[76])^(a[47] & b[77])^(a[46] & b[78])^(a[45] & b[79])^(a[44] & b[80])^(a[43] & b[81])^(a[42] & b[82])^(a[41] & b[83])^(a[40] & b[84])^(a[39] & b[85])^(a[38] & b[86])^(a[37] & b[87])^(a[36] & b[88])^(a[35] & b[89])^(a[34] & b[90])^(a[33] & b[91])^(a[32] & b[92])^(a[31] & b[93])^(a[30] & b[94])^(a[29] & b[95])^(a[28] & b[96])^(a[27] & b[97])^(a[26] & b[98])^(a[25] & b[99])^(a[24] & b[100])^(a[23] & b[101])^(a[22] & b[102])^(a[21] & b[103])^(a[20] & b[104])^(a[19] & b[105])^(a[18] & b[106])^(a[17] & b[107])^(a[16] & b[108])^(a[15] & b[109])^(a[14] & b[110])^(a[13] & b[111])^(a[12] & b[112])^(a[11] & b[113])^(a[10] & b[114])^(a[9] & b[115])^(a[8] & b[116])^(a[7] & b[117])^(a[6] & b[118])^(a[5] & b[119])^(a[4] & b[120])^(a[3] & b[121])^(a[2] & b[122])^(a[1] & b[123])^(a[0] & b[124]);
assign y[125] = (a[125] & b[0])^(a[124] & b[1])^(a[123] & b[2])^(a[122] & b[3])^(a[121] & b[4])^(a[120] & b[5])^(a[119] & b[6])^(a[118] & b[7])^(a[117] & b[8])^(a[116] & b[9])^(a[115] & b[10])^(a[114] & b[11])^(a[113] & b[12])^(a[112] & b[13])^(a[111] & b[14])^(a[110] & b[15])^(a[109] & b[16])^(a[108] & b[17])^(a[107] & b[18])^(a[106] & b[19])^(a[105] & b[20])^(a[104] & b[21])^(a[103] & b[22])^(a[102] & b[23])^(a[101] & b[24])^(a[100] & b[25])^(a[99] & b[26])^(a[98] & b[27])^(a[97] & b[28])^(a[96] & b[29])^(a[95] & b[30])^(a[94] & b[31])^(a[93] & b[32])^(a[92] & b[33])^(a[91] & b[34])^(a[90] & b[35])^(a[89] & b[36])^(a[88] & b[37])^(a[87] & b[38])^(a[86] & b[39])^(a[85] & b[40])^(a[84] & b[41])^(a[83] & b[42])^(a[82] & b[43])^(a[81] & b[44])^(a[80] & b[45])^(a[79] & b[46])^(a[78] & b[47])^(a[77] & b[48])^(a[76] & b[49])^(a[75] & b[50])^(a[74] & b[51])^(a[73] & b[52])^(a[72] & b[53])^(a[71] & b[54])^(a[70] & b[55])^(a[69] & b[56])^(a[68] & b[57])^(a[67] & b[58])^(a[66] & b[59])^(a[65] & b[60])^(a[64] & b[61])^(a[63] & b[62])^(a[62] & b[63])^(a[61] & b[64])^(a[60] & b[65])^(a[59] & b[66])^(a[58] & b[67])^(a[57] & b[68])^(a[56] & b[69])^(a[55] & b[70])^(a[54] & b[71])^(a[53] & b[72])^(a[52] & b[73])^(a[51] & b[74])^(a[50] & b[75])^(a[49] & b[76])^(a[48] & b[77])^(a[47] & b[78])^(a[46] & b[79])^(a[45] & b[80])^(a[44] & b[81])^(a[43] & b[82])^(a[42] & b[83])^(a[41] & b[84])^(a[40] & b[85])^(a[39] & b[86])^(a[38] & b[87])^(a[37] & b[88])^(a[36] & b[89])^(a[35] & b[90])^(a[34] & b[91])^(a[33] & b[92])^(a[32] & b[93])^(a[31] & b[94])^(a[30] & b[95])^(a[29] & b[96])^(a[28] & b[97])^(a[27] & b[98])^(a[26] & b[99])^(a[25] & b[100])^(a[24] & b[101])^(a[23] & b[102])^(a[22] & b[103])^(a[21] & b[104])^(a[20] & b[105])^(a[19] & b[106])^(a[18] & b[107])^(a[17] & b[108])^(a[16] & b[109])^(a[15] & b[110])^(a[14] & b[111])^(a[13] & b[112])^(a[12] & b[113])^(a[11] & b[114])^(a[10] & b[115])^(a[9] & b[116])^(a[8] & b[117])^(a[7] & b[118])^(a[6] & b[119])^(a[5] & b[120])^(a[4] & b[121])^(a[3] & b[122])^(a[2] & b[123])^(a[1] & b[124])^(a[0] & b[125]);
assign y[126] = (a[126] & b[0])^(a[125] & b[1])^(a[124] & b[2])^(a[123] & b[3])^(a[122] & b[4])^(a[121] & b[5])^(a[120] & b[6])^(a[119] & b[7])^(a[118] & b[8])^(a[117] & b[9])^(a[116] & b[10])^(a[115] & b[11])^(a[114] & b[12])^(a[113] & b[13])^(a[112] & b[14])^(a[111] & b[15])^(a[110] & b[16])^(a[109] & b[17])^(a[108] & b[18])^(a[107] & b[19])^(a[106] & b[20])^(a[105] & b[21])^(a[104] & b[22])^(a[103] & b[23])^(a[102] & b[24])^(a[101] & b[25])^(a[100] & b[26])^(a[99] & b[27])^(a[98] & b[28])^(a[97] & b[29])^(a[96] & b[30])^(a[95] & b[31])^(a[94] & b[32])^(a[93] & b[33])^(a[92] & b[34])^(a[91] & b[35])^(a[90] & b[36])^(a[89] & b[37])^(a[88] & b[38])^(a[87] & b[39])^(a[86] & b[40])^(a[85] & b[41])^(a[84] & b[42])^(a[83] & b[43])^(a[82] & b[44])^(a[81] & b[45])^(a[80] & b[46])^(a[79] & b[47])^(a[78] & b[48])^(a[77] & b[49])^(a[76] & b[50])^(a[75] & b[51])^(a[74] & b[52])^(a[73] & b[53])^(a[72] & b[54])^(a[71] & b[55])^(a[70] & b[56])^(a[69] & b[57])^(a[68] & b[58])^(a[67] & b[59])^(a[66] & b[60])^(a[65] & b[61])^(a[64] & b[62])^(a[63] & b[63])^(a[62] & b[64])^(a[61] & b[65])^(a[60] & b[66])^(a[59] & b[67])^(a[58] & b[68])^(a[57] & b[69])^(a[56] & b[70])^(a[55] & b[71])^(a[54] & b[72])^(a[53] & b[73])^(a[52] & b[74])^(a[51] & b[75])^(a[50] & b[76])^(a[49] & b[77])^(a[48] & b[78])^(a[47] & b[79])^(a[46] & b[80])^(a[45] & b[81])^(a[44] & b[82])^(a[43] & b[83])^(a[42] & b[84])^(a[41] & b[85])^(a[40] & b[86])^(a[39] & b[87])^(a[38] & b[88])^(a[37] & b[89])^(a[36] & b[90])^(a[35] & b[91])^(a[34] & b[92])^(a[33] & b[93])^(a[32] & b[94])^(a[31] & b[95])^(a[30] & b[96])^(a[29] & b[97])^(a[28] & b[98])^(a[27] & b[99])^(a[26] & b[100])^(a[25] & b[101])^(a[24] & b[102])^(a[23] & b[103])^(a[22] & b[104])^(a[21] & b[105])^(a[20] & b[106])^(a[19] & b[107])^(a[18] & b[108])^(a[17] & b[109])^(a[16] & b[110])^(a[15] & b[111])^(a[14] & b[112])^(a[13] & b[113])^(a[12] & b[114])^(a[11] & b[115])^(a[10] & b[116])^(a[9] & b[117])^(a[8] & b[118])^(a[7] & b[119])^(a[6] & b[120])^(a[5] & b[121])^(a[4] & b[122])^(a[3] & b[123])^(a[2] & b[124])^(a[1] & b[125])^(a[0] & b[126]);
assign y[127] = (a[127] & b[0])^(a[126] & b[1])^(a[125] & b[2])^(a[124] & b[3])^(a[123] & b[4])^(a[122] & b[5])^(a[121] & b[6])^(a[120] & b[7])^(a[119] & b[8])^(a[118] & b[9])^(a[117] & b[10])^(a[116] & b[11])^(a[115] & b[12])^(a[114] & b[13])^(a[113] & b[14])^(a[112] & b[15])^(a[111] & b[16])^(a[110] & b[17])^(a[109] & b[18])^(a[108] & b[19])^(a[107] & b[20])^(a[106] & b[21])^(a[105] & b[22])^(a[104] & b[23])^(a[103] & b[24])^(a[102] & b[25])^(a[101] & b[26])^(a[100] & b[27])^(a[99] & b[28])^(a[98] & b[29])^(a[97] & b[30])^(a[96] & b[31])^(a[95] & b[32])^(a[94] & b[33])^(a[93] & b[34])^(a[92] & b[35])^(a[91] & b[36])^(a[90] & b[37])^(a[89] & b[38])^(a[88] & b[39])^(a[87] & b[40])^(a[86] & b[41])^(a[85] & b[42])^(a[84] & b[43])^(a[83] & b[44])^(a[82] & b[45])^(a[81] & b[46])^(a[80] & b[47])^(a[79] & b[48])^(a[78] & b[49])^(a[77] & b[50])^(a[76] & b[51])^(a[75] & b[52])^(a[74] & b[53])^(a[73] & b[54])^(a[72] & b[55])^(a[71] & b[56])^(a[70] & b[57])^(a[69] & b[58])^(a[68] & b[59])^(a[67] & b[60])^(a[66] & b[61])^(a[65] & b[62])^(a[64] & b[63])^(a[63] & b[64])^(a[62] & b[65])^(a[61] & b[66])^(a[60] & b[67])^(a[59] & b[68])^(a[58] & b[69])^(a[57] & b[70])^(a[56] & b[71])^(a[55] & b[72])^(a[54] & b[73])^(a[53] & b[74])^(a[52] & b[75])^(a[51] & b[76])^(a[50] & b[77])^(a[49] & b[78])^(a[48] & b[79])^(a[47] & b[80])^(a[46] & b[81])^(a[45] & b[82])^(a[44] & b[83])^(a[43] & b[84])^(a[42] & b[85])^(a[41] & b[86])^(a[40] & b[87])^(a[39] & b[88])^(a[38] & b[89])^(a[37] & b[90])^(a[36] & b[91])^(a[35] & b[92])^(a[34] & b[93])^(a[33] & b[94])^(a[32] & b[95])^(a[31] & b[96])^(a[30] & b[97])^(a[29] & b[98])^(a[28] & b[99])^(a[27] & b[100])^(a[26] & b[101])^(a[25] & b[102])^(a[24] & b[103])^(a[23] & b[104])^(a[22] & b[105])^(a[21] & b[106])^(a[20] & b[107])^(a[19] & b[108])^(a[18] & b[109])^(a[17] & b[110])^(a[16] & b[111])^(a[15] & b[112])^(a[14] & b[113])^(a[13] & b[114])^(a[12] & b[115])^(a[11] & b[116])^(a[10] & b[117])^(a[9] & b[118])^(a[8] & b[119])^(a[7] & b[120])^(a[6] & b[121])^(a[5] & b[122])^(a[4] & b[123])^(a[3] & b[124])^(a[2] & b[125])^(a[1] & b[126])^(a[0] & b[127]);
assign y[128] = (a[128] & b[0])^(a[127] & b[1])^(a[126] & b[2])^(a[125] & b[3])^(a[124] & b[4])^(a[123] & b[5])^(a[122] & b[6])^(a[121] & b[7])^(a[120] & b[8])^(a[119] & b[9])^(a[118] & b[10])^(a[117] & b[11])^(a[116] & b[12])^(a[115] & b[13])^(a[114] & b[14])^(a[113] & b[15])^(a[112] & b[16])^(a[111] & b[17])^(a[110] & b[18])^(a[109] & b[19])^(a[108] & b[20])^(a[107] & b[21])^(a[106] & b[22])^(a[105] & b[23])^(a[104] & b[24])^(a[103] & b[25])^(a[102] & b[26])^(a[101] & b[27])^(a[100] & b[28])^(a[99] & b[29])^(a[98] & b[30])^(a[97] & b[31])^(a[96] & b[32])^(a[95] & b[33])^(a[94] & b[34])^(a[93] & b[35])^(a[92] & b[36])^(a[91] & b[37])^(a[90] & b[38])^(a[89] & b[39])^(a[88] & b[40])^(a[87] & b[41])^(a[86] & b[42])^(a[85] & b[43])^(a[84] & b[44])^(a[83] & b[45])^(a[82] & b[46])^(a[81] & b[47])^(a[80] & b[48])^(a[79] & b[49])^(a[78] & b[50])^(a[77] & b[51])^(a[76] & b[52])^(a[75] & b[53])^(a[74] & b[54])^(a[73] & b[55])^(a[72] & b[56])^(a[71] & b[57])^(a[70] & b[58])^(a[69] & b[59])^(a[68] & b[60])^(a[67] & b[61])^(a[66] & b[62])^(a[65] & b[63])^(a[64] & b[64])^(a[63] & b[65])^(a[62] & b[66])^(a[61] & b[67])^(a[60] & b[68])^(a[59] & b[69])^(a[58] & b[70])^(a[57] & b[71])^(a[56] & b[72])^(a[55] & b[73])^(a[54] & b[74])^(a[53] & b[75])^(a[52] & b[76])^(a[51] & b[77])^(a[50] & b[78])^(a[49] & b[79])^(a[48] & b[80])^(a[47] & b[81])^(a[46] & b[82])^(a[45] & b[83])^(a[44] & b[84])^(a[43] & b[85])^(a[42] & b[86])^(a[41] & b[87])^(a[40] & b[88])^(a[39] & b[89])^(a[38] & b[90])^(a[37] & b[91])^(a[36] & b[92])^(a[35] & b[93])^(a[34] & b[94])^(a[33] & b[95])^(a[32] & b[96])^(a[31] & b[97])^(a[30] & b[98])^(a[29] & b[99])^(a[28] & b[100])^(a[27] & b[101])^(a[26] & b[102])^(a[25] & b[103])^(a[24] & b[104])^(a[23] & b[105])^(a[22] & b[106])^(a[21] & b[107])^(a[20] & b[108])^(a[19] & b[109])^(a[18] & b[110])^(a[17] & b[111])^(a[16] & b[112])^(a[15] & b[113])^(a[14] & b[114])^(a[13] & b[115])^(a[12] & b[116])^(a[11] & b[117])^(a[10] & b[118])^(a[9] & b[119])^(a[8] & b[120])^(a[7] & b[121])^(a[6] & b[122])^(a[5] & b[123])^(a[4] & b[124])^(a[3] & b[125])^(a[2] & b[126])^(a[1] & b[127])^(a[0] & b[128]);
assign y[129] = (a[129] & b[0])^(a[128] & b[1])^(a[127] & b[2])^(a[126] & b[3])^(a[125] & b[4])^(a[124] & b[5])^(a[123] & b[6])^(a[122] & b[7])^(a[121] & b[8])^(a[120] & b[9])^(a[119] & b[10])^(a[118] & b[11])^(a[117] & b[12])^(a[116] & b[13])^(a[115] & b[14])^(a[114] & b[15])^(a[113] & b[16])^(a[112] & b[17])^(a[111] & b[18])^(a[110] & b[19])^(a[109] & b[20])^(a[108] & b[21])^(a[107] & b[22])^(a[106] & b[23])^(a[105] & b[24])^(a[104] & b[25])^(a[103] & b[26])^(a[102] & b[27])^(a[101] & b[28])^(a[100] & b[29])^(a[99] & b[30])^(a[98] & b[31])^(a[97] & b[32])^(a[96] & b[33])^(a[95] & b[34])^(a[94] & b[35])^(a[93] & b[36])^(a[92] & b[37])^(a[91] & b[38])^(a[90] & b[39])^(a[89] & b[40])^(a[88] & b[41])^(a[87] & b[42])^(a[86] & b[43])^(a[85] & b[44])^(a[84] & b[45])^(a[83] & b[46])^(a[82] & b[47])^(a[81] & b[48])^(a[80] & b[49])^(a[79] & b[50])^(a[78] & b[51])^(a[77] & b[52])^(a[76] & b[53])^(a[75] & b[54])^(a[74] & b[55])^(a[73] & b[56])^(a[72] & b[57])^(a[71] & b[58])^(a[70] & b[59])^(a[69] & b[60])^(a[68] & b[61])^(a[67] & b[62])^(a[66] & b[63])^(a[65] & b[64])^(a[64] & b[65])^(a[63] & b[66])^(a[62] & b[67])^(a[61] & b[68])^(a[60] & b[69])^(a[59] & b[70])^(a[58] & b[71])^(a[57] & b[72])^(a[56] & b[73])^(a[55] & b[74])^(a[54] & b[75])^(a[53] & b[76])^(a[52] & b[77])^(a[51] & b[78])^(a[50] & b[79])^(a[49] & b[80])^(a[48] & b[81])^(a[47] & b[82])^(a[46] & b[83])^(a[45] & b[84])^(a[44] & b[85])^(a[43] & b[86])^(a[42] & b[87])^(a[41] & b[88])^(a[40] & b[89])^(a[39] & b[90])^(a[38] & b[91])^(a[37] & b[92])^(a[36] & b[93])^(a[35] & b[94])^(a[34] & b[95])^(a[33] & b[96])^(a[32] & b[97])^(a[31] & b[98])^(a[30] & b[99])^(a[29] & b[100])^(a[28] & b[101])^(a[27] & b[102])^(a[26] & b[103])^(a[25] & b[104])^(a[24] & b[105])^(a[23] & b[106])^(a[22] & b[107])^(a[21] & b[108])^(a[20] & b[109])^(a[19] & b[110])^(a[18] & b[111])^(a[17] & b[112])^(a[16] & b[113])^(a[15] & b[114])^(a[14] & b[115])^(a[13] & b[116])^(a[12] & b[117])^(a[11] & b[118])^(a[10] & b[119])^(a[9] & b[120])^(a[8] & b[121])^(a[7] & b[122])^(a[6] & b[123])^(a[5] & b[124])^(a[4] & b[125])^(a[3] & b[126])^(a[2] & b[127])^(a[1] & b[128])^(a[0] & b[129]);
assign y[130] = (a[130] & b[0])^(a[129] & b[1])^(a[128] & b[2])^(a[127] & b[3])^(a[126] & b[4])^(a[125] & b[5])^(a[124] & b[6])^(a[123] & b[7])^(a[122] & b[8])^(a[121] & b[9])^(a[120] & b[10])^(a[119] & b[11])^(a[118] & b[12])^(a[117] & b[13])^(a[116] & b[14])^(a[115] & b[15])^(a[114] & b[16])^(a[113] & b[17])^(a[112] & b[18])^(a[111] & b[19])^(a[110] & b[20])^(a[109] & b[21])^(a[108] & b[22])^(a[107] & b[23])^(a[106] & b[24])^(a[105] & b[25])^(a[104] & b[26])^(a[103] & b[27])^(a[102] & b[28])^(a[101] & b[29])^(a[100] & b[30])^(a[99] & b[31])^(a[98] & b[32])^(a[97] & b[33])^(a[96] & b[34])^(a[95] & b[35])^(a[94] & b[36])^(a[93] & b[37])^(a[92] & b[38])^(a[91] & b[39])^(a[90] & b[40])^(a[89] & b[41])^(a[88] & b[42])^(a[87] & b[43])^(a[86] & b[44])^(a[85] & b[45])^(a[84] & b[46])^(a[83] & b[47])^(a[82] & b[48])^(a[81] & b[49])^(a[80] & b[50])^(a[79] & b[51])^(a[78] & b[52])^(a[77] & b[53])^(a[76] & b[54])^(a[75] & b[55])^(a[74] & b[56])^(a[73] & b[57])^(a[72] & b[58])^(a[71] & b[59])^(a[70] & b[60])^(a[69] & b[61])^(a[68] & b[62])^(a[67] & b[63])^(a[66] & b[64])^(a[65] & b[65])^(a[64] & b[66])^(a[63] & b[67])^(a[62] & b[68])^(a[61] & b[69])^(a[60] & b[70])^(a[59] & b[71])^(a[58] & b[72])^(a[57] & b[73])^(a[56] & b[74])^(a[55] & b[75])^(a[54] & b[76])^(a[53] & b[77])^(a[52] & b[78])^(a[51] & b[79])^(a[50] & b[80])^(a[49] & b[81])^(a[48] & b[82])^(a[47] & b[83])^(a[46] & b[84])^(a[45] & b[85])^(a[44] & b[86])^(a[43] & b[87])^(a[42] & b[88])^(a[41] & b[89])^(a[40] & b[90])^(a[39] & b[91])^(a[38] & b[92])^(a[37] & b[93])^(a[36] & b[94])^(a[35] & b[95])^(a[34] & b[96])^(a[33] & b[97])^(a[32] & b[98])^(a[31] & b[99])^(a[30] & b[100])^(a[29] & b[101])^(a[28] & b[102])^(a[27] & b[103])^(a[26] & b[104])^(a[25] & b[105])^(a[24] & b[106])^(a[23] & b[107])^(a[22] & b[108])^(a[21] & b[109])^(a[20] & b[110])^(a[19] & b[111])^(a[18] & b[112])^(a[17] & b[113])^(a[16] & b[114])^(a[15] & b[115])^(a[14] & b[116])^(a[13] & b[117])^(a[12] & b[118])^(a[11] & b[119])^(a[10] & b[120])^(a[9] & b[121])^(a[8] & b[122])^(a[7] & b[123])^(a[6] & b[124])^(a[5] & b[125])^(a[4] & b[126])^(a[3] & b[127])^(a[2] & b[128])^(a[1] & b[129])^(a[0] & b[130]);
assign y[131] = (a[131] & b[0])^(a[130] & b[1])^(a[129] & b[2])^(a[128] & b[3])^(a[127] & b[4])^(a[126] & b[5])^(a[125] & b[6])^(a[124] & b[7])^(a[123] & b[8])^(a[122] & b[9])^(a[121] & b[10])^(a[120] & b[11])^(a[119] & b[12])^(a[118] & b[13])^(a[117] & b[14])^(a[116] & b[15])^(a[115] & b[16])^(a[114] & b[17])^(a[113] & b[18])^(a[112] & b[19])^(a[111] & b[20])^(a[110] & b[21])^(a[109] & b[22])^(a[108] & b[23])^(a[107] & b[24])^(a[106] & b[25])^(a[105] & b[26])^(a[104] & b[27])^(a[103] & b[28])^(a[102] & b[29])^(a[101] & b[30])^(a[100] & b[31])^(a[99] & b[32])^(a[98] & b[33])^(a[97] & b[34])^(a[96] & b[35])^(a[95] & b[36])^(a[94] & b[37])^(a[93] & b[38])^(a[92] & b[39])^(a[91] & b[40])^(a[90] & b[41])^(a[89] & b[42])^(a[88] & b[43])^(a[87] & b[44])^(a[86] & b[45])^(a[85] & b[46])^(a[84] & b[47])^(a[83] & b[48])^(a[82] & b[49])^(a[81] & b[50])^(a[80] & b[51])^(a[79] & b[52])^(a[78] & b[53])^(a[77] & b[54])^(a[76] & b[55])^(a[75] & b[56])^(a[74] & b[57])^(a[73] & b[58])^(a[72] & b[59])^(a[71] & b[60])^(a[70] & b[61])^(a[69] & b[62])^(a[68] & b[63])^(a[67] & b[64])^(a[66] & b[65])^(a[65] & b[66])^(a[64] & b[67])^(a[63] & b[68])^(a[62] & b[69])^(a[61] & b[70])^(a[60] & b[71])^(a[59] & b[72])^(a[58] & b[73])^(a[57] & b[74])^(a[56] & b[75])^(a[55] & b[76])^(a[54] & b[77])^(a[53] & b[78])^(a[52] & b[79])^(a[51] & b[80])^(a[50] & b[81])^(a[49] & b[82])^(a[48] & b[83])^(a[47] & b[84])^(a[46] & b[85])^(a[45] & b[86])^(a[44] & b[87])^(a[43] & b[88])^(a[42] & b[89])^(a[41] & b[90])^(a[40] & b[91])^(a[39] & b[92])^(a[38] & b[93])^(a[37] & b[94])^(a[36] & b[95])^(a[35] & b[96])^(a[34] & b[97])^(a[33] & b[98])^(a[32] & b[99])^(a[31] & b[100])^(a[30] & b[101])^(a[29] & b[102])^(a[28] & b[103])^(a[27] & b[104])^(a[26] & b[105])^(a[25] & b[106])^(a[24] & b[107])^(a[23] & b[108])^(a[22] & b[109])^(a[21] & b[110])^(a[20] & b[111])^(a[19] & b[112])^(a[18] & b[113])^(a[17] & b[114])^(a[16] & b[115])^(a[15] & b[116])^(a[14] & b[117])^(a[13] & b[118])^(a[12] & b[119])^(a[11] & b[120])^(a[10] & b[121])^(a[9] & b[122])^(a[8] & b[123])^(a[7] & b[124])^(a[6] & b[125])^(a[5] & b[126])^(a[4] & b[127])^(a[3] & b[128])^(a[2] & b[129])^(a[1] & b[130])^(a[0] & b[131]);
assign y[132] = (a[132] & b[0])^(a[131] & b[1])^(a[130] & b[2])^(a[129] & b[3])^(a[128] & b[4])^(a[127] & b[5])^(a[126] & b[6])^(a[125] & b[7])^(a[124] & b[8])^(a[123] & b[9])^(a[122] & b[10])^(a[121] & b[11])^(a[120] & b[12])^(a[119] & b[13])^(a[118] & b[14])^(a[117] & b[15])^(a[116] & b[16])^(a[115] & b[17])^(a[114] & b[18])^(a[113] & b[19])^(a[112] & b[20])^(a[111] & b[21])^(a[110] & b[22])^(a[109] & b[23])^(a[108] & b[24])^(a[107] & b[25])^(a[106] & b[26])^(a[105] & b[27])^(a[104] & b[28])^(a[103] & b[29])^(a[102] & b[30])^(a[101] & b[31])^(a[100] & b[32])^(a[99] & b[33])^(a[98] & b[34])^(a[97] & b[35])^(a[96] & b[36])^(a[95] & b[37])^(a[94] & b[38])^(a[93] & b[39])^(a[92] & b[40])^(a[91] & b[41])^(a[90] & b[42])^(a[89] & b[43])^(a[88] & b[44])^(a[87] & b[45])^(a[86] & b[46])^(a[85] & b[47])^(a[84] & b[48])^(a[83] & b[49])^(a[82] & b[50])^(a[81] & b[51])^(a[80] & b[52])^(a[79] & b[53])^(a[78] & b[54])^(a[77] & b[55])^(a[76] & b[56])^(a[75] & b[57])^(a[74] & b[58])^(a[73] & b[59])^(a[72] & b[60])^(a[71] & b[61])^(a[70] & b[62])^(a[69] & b[63])^(a[68] & b[64])^(a[67] & b[65])^(a[66] & b[66])^(a[65] & b[67])^(a[64] & b[68])^(a[63] & b[69])^(a[62] & b[70])^(a[61] & b[71])^(a[60] & b[72])^(a[59] & b[73])^(a[58] & b[74])^(a[57] & b[75])^(a[56] & b[76])^(a[55] & b[77])^(a[54] & b[78])^(a[53] & b[79])^(a[52] & b[80])^(a[51] & b[81])^(a[50] & b[82])^(a[49] & b[83])^(a[48] & b[84])^(a[47] & b[85])^(a[46] & b[86])^(a[45] & b[87])^(a[44] & b[88])^(a[43] & b[89])^(a[42] & b[90])^(a[41] & b[91])^(a[40] & b[92])^(a[39] & b[93])^(a[38] & b[94])^(a[37] & b[95])^(a[36] & b[96])^(a[35] & b[97])^(a[34] & b[98])^(a[33] & b[99])^(a[32] & b[100])^(a[31] & b[101])^(a[30] & b[102])^(a[29] & b[103])^(a[28] & b[104])^(a[27] & b[105])^(a[26] & b[106])^(a[25] & b[107])^(a[24] & b[108])^(a[23] & b[109])^(a[22] & b[110])^(a[21] & b[111])^(a[20] & b[112])^(a[19] & b[113])^(a[18] & b[114])^(a[17] & b[115])^(a[16] & b[116])^(a[15] & b[117])^(a[14] & b[118])^(a[13] & b[119])^(a[12] & b[120])^(a[11] & b[121])^(a[10] & b[122])^(a[9] & b[123])^(a[8] & b[124])^(a[7] & b[125])^(a[6] & b[126])^(a[5] & b[127])^(a[4] & b[128])^(a[3] & b[129])^(a[2] & b[130])^(a[1] & b[131])^(a[0] & b[132]);
assign y[133] = (a[133] & b[0])^(a[132] & b[1])^(a[131] & b[2])^(a[130] & b[3])^(a[129] & b[4])^(a[128] & b[5])^(a[127] & b[6])^(a[126] & b[7])^(a[125] & b[8])^(a[124] & b[9])^(a[123] & b[10])^(a[122] & b[11])^(a[121] & b[12])^(a[120] & b[13])^(a[119] & b[14])^(a[118] & b[15])^(a[117] & b[16])^(a[116] & b[17])^(a[115] & b[18])^(a[114] & b[19])^(a[113] & b[20])^(a[112] & b[21])^(a[111] & b[22])^(a[110] & b[23])^(a[109] & b[24])^(a[108] & b[25])^(a[107] & b[26])^(a[106] & b[27])^(a[105] & b[28])^(a[104] & b[29])^(a[103] & b[30])^(a[102] & b[31])^(a[101] & b[32])^(a[100] & b[33])^(a[99] & b[34])^(a[98] & b[35])^(a[97] & b[36])^(a[96] & b[37])^(a[95] & b[38])^(a[94] & b[39])^(a[93] & b[40])^(a[92] & b[41])^(a[91] & b[42])^(a[90] & b[43])^(a[89] & b[44])^(a[88] & b[45])^(a[87] & b[46])^(a[86] & b[47])^(a[85] & b[48])^(a[84] & b[49])^(a[83] & b[50])^(a[82] & b[51])^(a[81] & b[52])^(a[80] & b[53])^(a[79] & b[54])^(a[78] & b[55])^(a[77] & b[56])^(a[76] & b[57])^(a[75] & b[58])^(a[74] & b[59])^(a[73] & b[60])^(a[72] & b[61])^(a[71] & b[62])^(a[70] & b[63])^(a[69] & b[64])^(a[68] & b[65])^(a[67] & b[66])^(a[66] & b[67])^(a[65] & b[68])^(a[64] & b[69])^(a[63] & b[70])^(a[62] & b[71])^(a[61] & b[72])^(a[60] & b[73])^(a[59] & b[74])^(a[58] & b[75])^(a[57] & b[76])^(a[56] & b[77])^(a[55] & b[78])^(a[54] & b[79])^(a[53] & b[80])^(a[52] & b[81])^(a[51] & b[82])^(a[50] & b[83])^(a[49] & b[84])^(a[48] & b[85])^(a[47] & b[86])^(a[46] & b[87])^(a[45] & b[88])^(a[44] & b[89])^(a[43] & b[90])^(a[42] & b[91])^(a[41] & b[92])^(a[40] & b[93])^(a[39] & b[94])^(a[38] & b[95])^(a[37] & b[96])^(a[36] & b[97])^(a[35] & b[98])^(a[34] & b[99])^(a[33] & b[100])^(a[32] & b[101])^(a[31] & b[102])^(a[30] & b[103])^(a[29] & b[104])^(a[28] & b[105])^(a[27] & b[106])^(a[26] & b[107])^(a[25] & b[108])^(a[24] & b[109])^(a[23] & b[110])^(a[22] & b[111])^(a[21] & b[112])^(a[20] & b[113])^(a[19] & b[114])^(a[18] & b[115])^(a[17] & b[116])^(a[16] & b[117])^(a[15] & b[118])^(a[14] & b[119])^(a[13] & b[120])^(a[12] & b[121])^(a[11] & b[122])^(a[10] & b[123])^(a[9] & b[124])^(a[8] & b[125])^(a[7] & b[126])^(a[6] & b[127])^(a[5] & b[128])^(a[4] & b[129])^(a[3] & b[130])^(a[2] & b[131])^(a[1] & b[132])^(a[0] & b[133]);
assign y[134] = (a[134] & b[0])^(a[133] & b[1])^(a[132] & b[2])^(a[131] & b[3])^(a[130] & b[4])^(a[129] & b[5])^(a[128] & b[6])^(a[127] & b[7])^(a[126] & b[8])^(a[125] & b[9])^(a[124] & b[10])^(a[123] & b[11])^(a[122] & b[12])^(a[121] & b[13])^(a[120] & b[14])^(a[119] & b[15])^(a[118] & b[16])^(a[117] & b[17])^(a[116] & b[18])^(a[115] & b[19])^(a[114] & b[20])^(a[113] & b[21])^(a[112] & b[22])^(a[111] & b[23])^(a[110] & b[24])^(a[109] & b[25])^(a[108] & b[26])^(a[107] & b[27])^(a[106] & b[28])^(a[105] & b[29])^(a[104] & b[30])^(a[103] & b[31])^(a[102] & b[32])^(a[101] & b[33])^(a[100] & b[34])^(a[99] & b[35])^(a[98] & b[36])^(a[97] & b[37])^(a[96] & b[38])^(a[95] & b[39])^(a[94] & b[40])^(a[93] & b[41])^(a[92] & b[42])^(a[91] & b[43])^(a[90] & b[44])^(a[89] & b[45])^(a[88] & b[46])^(a[87] & b[47])^(a[86] & b[48])^(a[85] & b[49])^(a[84] & b[50])^(a[83] & b[51])^(a[82] & b[52])^(a[81] & b[53])^(a[80] & b[54])^(a[79] & b[55])^(a[78] & b[56])^(a[77] & b[57])^(a[76] & b[58])^(a[75] & b[59])^(a[74] & b[60])^(a[73] & b[61])^(a[72] & b[62])^(a[71] & b[63])^(a[70] & b[64])^(a[69] & b[65])^(a[68] & b[66])^(a[67] & b[67])^(a[66] & b[68])^(a[65] & b[69])^(a[64] & b[70])^(a[63] & b[71])^(a[62] & b[72])^(a[61] & b[73])^(a[60] & b[74])^(a[59] & b[75])^(a[58] & b[76])^(a[57] & b[77])^(a[56] & b[78])^(a[55] & b[79])^(a[54] & b[80])^(a[53] & b[81])^(a[52] & b[82])^(a[51] & b[83])^(a[50] & b[84])^(a[49] & b[85])^(a[48] & b[86])^(a[47] & b[87])^(a[46] & b[88])^(a[45] & b[89])^(a[44] & b[90])^(a[43] & b[91])^(a[42] & b[92])^(a[41] & b[93])^(a[40] & b[94])^(a[39] & b[95])^(a[38] & b[96])^(a[37] & b[97])^(a[36] & b[98])^(a[35] & b[99])^(a[34] & b[100])^(a[33] & b[101])^(a[32] & b[102])^(a[31] & b[103])^(a[30] & b[104])^(a[29] & b[105])^(a[28] & b[106])^(a[27] & b[107])^(a[26] & b[108])^(a[25] & b[109])^(a[24] & b[110])^(a[23] & b[111])^(a[22] & b[112])^(a[21] & b[113])^(a[20] & b[114])^(a[19] & b[115])^(a[18] & b[116])^(a[17] & b[117])^(a[16] & b[118])^(a[15] & b[119])^(a[14] & b[120])^(a[13] & b[121])^(a[12] & b[122])^(a[11] & b[123])^(a[10] & b[124])^(a[9] & b[125])^(a[8] & b[126])^(a[7] & b[127])^(a[6] & b[128])^(a[5] & b[129])^(a[4] & b[130])^(a[3] & b[131])^(a[2] & b[132])^(a[1] & b[133])^(a[0] & b[134]);
assign y[135] = (a[135] & b[0])^(a[134] & b[1])^(a[133] & b[2])^(a[132] & b[3])^(a[131] & b[4])^(a[130] & b[5])^(a[129] & b[6])^(a[128] & b[7])^(a[127] & b[8])^(a[126] & b[9])^(a[125] & b[10])^(a[124] & b[11])^(a[123] & b[12])^(a[122] & b[13])^(a[121] & b[14])^(a[120] & b[15])^(a[119] & b[16])^(a[118] & b[17])^(a[117] & b[18])^(a[116] & b[19])^(a[115] & b[20])^(a[114] & b[21])^(a[113] & b[22])^(a[112] & b[23])^(a[111] & b[24])^(a[110] & b[25])^(a[109] & b[26])^(a[108] & b[27])^(a[107] & b[28])^(a[106] & b[29])^(a[105] & b[30])^(a[104] & b[31])^(a[103] & b[32])^(a[102] & b[33])^(a[101] & b[34])^(a[100] & b[35])^(a[99] & b[36])^(a[98] & b[37])^(a[97] & b[38])^(a[96] & b[39])^(a[95] & b[40])^(a[94] & b[41])^(a[93] & b[42])^(a[92] & b[43])^(a[91] & b[44])^(a[90] & b[45])^(a[89] & b[46])^(a[88] & b[47])^(a[87] & b[48])^(a[86] & b[49])^(a[85] & b[50])^(a[84] & b[51])^(a[83] & b[52])^(a[82] & b[53])^(a[81] & b[54])^(a[80] & b[55])^(a[79] & b[56])^(a[78] & b[57])^(a[77] & b[58])^(a[76] & b[59])^(a[75] & b[60])^(a[74] & b[61])^(a[73] & b[62])^(a[72] & b[63])^(a[71] & b[64])^(a[70] & b[65])^(a[69] & b[66])^(a[68] & b[67])^(a[67] & b[68])^(a[66] & b[69])^(a[65] & b[70])^(a[64] & b[71])^(a[63] & b[72])^(a[62] & b[73])^(a[61] & b[74])^(a[60] & b[75])^(a[59] & b[76])^(a[58] & b[77])^(a[57] & b[78])^(a[56] & b[79])^(a[55] & b[80])^(a[54] & b[81])^(a[53] & b[82])^(a[52] & b[83])^(a[51] & b[84])^(a[50] & b[85])^(a[49] & b[86])^(a[48] & b[87])^(a[47] & b[88])^(a[46] & b[89])^(a[45] & b[90])^(a[44] & b[91])^(a[43] & b[92])^(a[42] & b[93])^(a[41] & b[94])^(a[40] & b[95])^(a[39] & b[96])^(a[38] & b[97])^(a[37] & b[98])^(a[36] & b[99])^(a[35] & b[100])^(a[34] & b[101])^(a[33] & b[102])^(a[32] & b[103])^(a[31] & b[104])^(a[30] & b[105])^(a[29] & b[106])^(a[28] & b[107])^(a[27] & b[108])^(a[26] & b[109])^(a[25] & b[110])^(a[24] & b[111])^(a[23] & b[112])^(a[22] & b[113])^(a[21] & b[114])^(a[20] & b[115])^(a[19] & b[116])^(a[18] & b[117])^(a[17] & b[118])^(a[16] & b[119])^(a[15] & b[120])^(a[14] & b[121])^(a[13] & b[122])^(a[12] & b[123])^(a[11] & b[124])^(a[10] & b[125])^(a[9] & b[126])^(a[8] & b[127])^(a[7] & b[128])^(a[6] & b[129])^(a[5] & b[130])^(a[4] & b[131])^(a[3] & b[132])^(a[2] & b[133])^(a[1] & b[134])^(a[0] & b[135]);
assign y[136] = (a[136] & b[0])^(a[135] & b[1])^(a[134] & b[2])^(a[133] & b[3])^(a[132] & b[4])^(a[131] & b[5])^(a[130] & b[6])^(a[129] & b[7])^(a[128] & b[8])^(a[127] & b[9])^(a[126] & b[10])^(a[125] & b[11])^(a[124] & b[12])^(a[123] & b[13])^(a[122] & b[14])^(a[121] & b[15])^(a[120] & b[16])^(a[119] & b[17])^(a[118] & b[18])^(a[117] & b[19])^(a[116] & b[20])^(a[115] & b[21])^(a[114] & b[22])^(a[113] & b[23])^(a[112] & b[24])^(a[111] & b[25])^(a[110] & b[26])^(a[109] & b[27])^(a[108] & b[28])^(a[107] & b[29])^(a[106] & b[30])^(a[105] & b[31])^(a[104] & b[32])^(a[103] & b[33])^(a[102] & b[34])^(a[101] & b[35])^(a[100] & b[36])^(a[99] & b[37])^(a[98] & b[38])^(a[97] & b[39])^(a[96] & b[40])^(a[95] & b[41])^(a[94] & b[42])^(a[93] & b[43])^(a[92] & b[44])^(a[91] & b[45])^(a[90] & b[46])^(a[89] & b[47])^(a[88] & b[48])^(a[87] & b[49])^(a[86] & b[50])^(a[85] & b[51])^(a[84] & b[52])^(a[83] & b[53])^(a[82] & b[54])^(a[81] & b[55])^(a[80] & b[56])^(a[79] & b[57])^(a[78] & b[58])^(a[77] & b[59])^(a[76] & b[60])^(a[75] & b[61])^(a[74] & b[62])^(a[73] & b[63])^(a[72] & b[64])^(a[71] & b[65])^(a[70] & b[66])^(a[69] & b[67])^(a[68] & b[68])^(a[67] & b[69])^(a[66] & b[70])^(a[65] & b[71])^(a[64] & b[72])^(a[63] & b[73])^(a[62] & b[74])^(a[61] & b[75])^(a[60] & b[76])^(a[59] & b[77])^(a[58] & b[78])^(a[57] & b[79])^(a[56] & b[80])^(a[55] & b[81])^(a[54] & b[82])^(a[53] & b[83])^(a[52] & b[84])^(a[51] & b[85])^(a[50] & b[86])^(a[49] & b[87])^(a[48] & b[88])^(a[47] & b[89])^(a[46] & b[90])^(a[45] & b[91])^(a[44] & b[92])^(a[43] & b[93])^(a[42] & b[94])^(a[41] & b[95])^(a[40] & b[96])^(a[39] & b[97])^(a[38] & b[98])^(a[37] & b[99])^(a[36] & b[100])^(a[35] & b[101])^(a[34] & b[102])^(a[33] & b[103])^(a[32] & b[104])^(a[31] & b[105])^(a[30] & b[106])^(a[29] & b[107])^(a[28] & b[108])^(a[27] & b[109])^(a[26] & b[110])^(a[25] & b[111])^(a[24] & b[112])^(a[23] & b[113])^(a[22] & b[114])^(a[21] & b[115])^(a[20] & b[116])^(a[19] & b[117])^(a[18] & b[118])^(a[17] & b[119])^(a[16] & b[120])^(a[15] & b[121])^(a[14] & b[122])^(a[13] & b[123])^(a[12] & b[124])^(a[11] & b[125])^(a[10] & b[126])^(a[9] & b[127])^(a[8] & b[128])^(a[7] & b[129])^(a[6] & b[130])^(a[5] & b[131])^(a[4] & b[132])^(a[3] & b[133])^(a[2] & b[134])^(a[1] & b[135])^(a[0] & b[136]);
assign y[137] = (a[137] & b[0])^(a[136] & b[1])^(a[135] & b[2])^(a[134] & b[3])^(a[133] & b[4])^(a[132] & b[5])^(a[131] & b[6])^(a[130] & b[7])^(a[129] & b[8])^(a[128] & b[9])^(a[127] & b[10])^(a[126] & b[11])^(a[125] & b[12])^(a[124] & b[13])^(a[123] & b[14])^(a[122] & b[15])^(a[121] & b[16])^(a[120] & b[17])^(a[119] & b[18])^(a[118] & b[19])^(a[117] & b[20])^(a[116] & b[21])^(a[115] & b[22])^(a[114] & b[23])^(a[113] & b[24])^(a[112] & b[25])^(a[111] & b[26])^(a[110] & b[27])^(a[109] & b[28])^(a[108] & b[29])^(a[107] & b[30])^(a[106] & b[31])^(a[105] & b[32])^(a[104] & b[33])^(a[103] & b[34])^(a[102] & b[35])^(a[101] & b[36])^(a[100] & b[37])^(a[99] & b[38])^(a[98] & b[39])^(a[97] & b[40])^(a[96] & b[41])^(a[95] & b[42])^(a[94] & b[43])^(a[93] & b[44])^(a[92] & b[45])^(a[91] & b[46])^(a[90] & b[47])^(a[89] & b[48])^(a[88] & b[49])^(a[87] & b[50])^(a[86] & b[51])^(a[85] & b[52])^(a[84] & b[53])^(a[83] & b[54])^(a[82] & b[55])^(a[81] & b[56])^(a[80] & b[57])^(a[79] & b[58])^(a[78] & b[59])^(a[77] & b[60])^(a[76] & b[61])^(a[75] & b[62])^(a[74] & b[63])^(a[73] & b[64])^(a[72] & b[65])^(a[71] & b[66])^(a[70] & b[67])^(a[69] & b[68])^(a[68] & b[69])^(a[67] & b[70])^(a[66] & b[71])^(a[65] & b[72])^(a[64] & b[73])^(a[63] & b[74])^(a[62] & b[75])^(a[61] & b[76])^(a[60] & b[77])^(a[59] & b[78])^(a[58] & b[79])^(a[57] & b[80])^(a[56] & b[81])^(a[55] & b[82])^(a[54] & b[83])^(a[53] & b[84])^(a[52] & b[85])^(a[51] & b[86])^(a[50] & b[87])^(a[49] & b[88])^(a[48] & b[89])^(a[47] & b[90])^(a[46] & b[91])^(a[45] & b[92])^(a[44] & b[93])^(a[43] & b[94])^(a[42] & b[95])^(a[41] & b[96])^(a[40] & b[97])^(a[39] & b[98])^(a[38] & b[99])^(a[37] & b[100])^(a[36] & b[101])^(a[35] & b[102])^(a[34] & b[103])^(a[33] & b[104])^(a[32] & b[105])^(a[31] & b[106])^(a[30] & b[107])^(a[29] & b[108])^(a[28] & b[109])^(a[27] & b[110])^(a[26] & b[111])^(a[25] & b[112])^(a[24] & b[113])^(a[23] & b[114])^(a[22] & b[115])^(a[21] & b[116])^(a[20] & b[117])^(a[19] & b[118])^(a[18] & b[119])^(a[17] & b[120])^(a[16] & b[121])^(a[15] & b[122])^(a[14] & b[123])^(a[13] & b[124])^(a[12] & b[125])^(a[11] & b[126])^(a[10] & b[127])^(a[9] & b[128])^(a[8] & b[129])^(a[7] & b[130])^(a[6] & b[131])^(a[5] & b[132])^(a[4] & b[133])^(a[3] & b[134])^(a[2] & b[135])^(a[1] & b[136])^(a[0] & b[137]);
assign y[138] = (a[138] & b[0])^(a[137] & b[1])^(a[136] & b[2])^(a[135] & b[3])^(a[134] & b[4])^(a[133] & b[5])^(a[132] & b[6])^(a[131] & b[7])^(a[130] & b[8])^(a[129] & b[9])^(a[128] & b[10])^(a[127] & b[11])^(a[126] & b[12])^(a[125] & b[13])^(a[124] & b[14])^(a[123] & b[15])^(a[122] & b[16])^(a[121] & b[17])^(a[120] & b[18])^(a[119] & b[19])^(a[118] & b[20])^(a[117] & b[21])^(a[116] & b[22])^(a[115] & b[23])^(a[114] & b[24])^(a[113] & b[25])^(a[112] & b[26])^(a[111] & b[27])^(a[110] & b[28])^(a[109] & b[29])^(a[108] & b[30])^(a[107] & b[31])^(a[106] & b[32])^(a[105] & b[33])^(a[104] & b[34])^(a[103] & b[35])^(a[102] & b[36])^(a[101] & b[37])^(a[100] & b[38])^(a[99] & b[39])^(a[98] & b[40])^(a[97] & b[41])^(a[96] & b[42])^(a[95] & b[43])^(a[94] & b[44])^(a[93] & b[45])^(a[92] & b[46])^(a[91] & b[47])^(a[90] & b[48])^(a[89] & b[49])^(a[88] & b[50])^(a[87] & b[51])^(a[86] & b[52])^(a[85] & b[53])^(a[84] & b[54])^(a[83] & b[55])^(a[82] & b[56])^(a[81] & b[57])^(a[80] & b[58])^(a[79] & b[59])^(a[78] & b[60])^(a[77] & b[61])^(a[76] & b[62])^(a[75] & b[63])^(a[74] & b[64])^(a[73] & b[65])^(a[72] & b[66])^(a[71] & b[67])^(a[70] & b[68])^(a[69] & b[69])^(a[68] & b[70])^(a[67] & b[71])^(a[66] & b[72])^(a[65] & b[73])^(a[64] & b[74])^(a[63] & b[75])^(a[62] & b[76])^(a[61] & b[77])^(a[60] & b[78])^(a[59] & b[79])^(a[58] & b[80])^(a[57] & b[81])^(a[56] & b[82])^(a[55] & b[83])^(a[54] & b[84])^(a[53] & b[85])^(a[52] & b[86])^(a[51] & b[87])^(a[50] & b[88])^(a[49] & b[89])^(a[48] & b[90])^(a[47] & b[91])^(a[46] & b[92])^(a[45] & b[93])^(a[44] & b[94])^(a[43] & b[95])^(a[42] & b[96])^(a[41] & b[97])^(a[40] & b[98])^(a[39] & b[99])^(a[38] & b[100])^(a[37] & b[101])^(a[36] & b[102])^(a[35] & b[103])^(a[34] & b[104])^(a[33] & b[105])^(a[32] & b[106])^(a[31] & b[107])^(a[30] & b[108])^(a[29] & b[109])^(a[28] & b[110])^(a[27] & b[111])^(a[26] & b[112])^(a[25] & b[113])^(a[24] & b[114])^(a[23] & b[115])^(a[22] & b[116])^(a[21] & b[117])^(a[20] & b[118])^(a[19] & b[119])^(a[18] & b[120])^(a[17] & b[121])^(a[16] & b[122])^(a[15] & b[123])^(a[14] & b[124])^(a[13] & b[125])^(a[12] & b[126])^(a[11] & b[127])^(a[10] & b[128])^(a[9] & b[129])^(a[8] & b[130])^(a[7] & b[131])^(a[6] & b[132])^(a[5] & b[133])^(a[4] & b[134])^(a[3] & b[135])^(a[2] & b[136])^(a[1] & b[137])^(a[0] & b[138]);
assign y[139] = (a[139] & b[0])^(a[138] & b[1])^(a[137] & b[2])^(a[136] & b[3])^(a[135] & b[4])^(a[134] & b[5])^(a[133] & b[6])^(a[132] & b[7])^(a[131] & b[8])^(a[130] & b[9])^(a[129] & b[10])^(a[128] & b[11])^(a[127] & b[12])^(a[126] & b[13])^(a[125] & b[14])^(a[124] & b[15])^(a[123] & b[16])^(a[122] & b[17])^(a[121] & b[18])^(a[120] & b[19])^(a[119] & b[20])^(a[118] & b[21])^(a[117] & b[22])^(a[116] & b[23])^(a[115] & b[24])^(a[114] & b[25])^(a[113] & b[26])^(a[112] & b[27])^(a[111] & b[28])^(a[110] & b[29])^(a[109] & b[30])^(a[108] & b[31])^(a[107] & b[32])^(a[106] & b[33])^(a[105] & b[34])^(a[104] & b[35])^(a[103] & b[36])^(a[102] & b[37])^(a[101] & b[38])^(a[100] & b[39])^(a[99] & b[40])^(a[98] & b[41])^(a[97] & b[42])^(a[96] & b[43])^(a[95] & b[44])^(a[94] & b[45])^(a[93] & b[46])^(a[92] & b[47])^(a[91] & b[48])^(a[90] & b[49])^(a[89] & b[50])^(a[88] & b[51])^(a[87] & b[52])^(a[86] & b[53])^(a[85] & b[54])^(a[84] & b[55])^(a[83] & b[56])^(a[82] & b[57])^(a[81] & b[58])^(a[80] & b[59])^(a[79] & b[60])^(a[78] & b[61])^(a[77] & b[62])^(a[76] & b[63])^(a[75] & b[64])^(a[74] & b[65])^(a[73] & b[66])^(a[72] & b[67])^(a[71] & b[68])^(a[70] & b[69])^(a[69] & b[70])^(a[68] & b[71])^(a[67] & b[72])^(a[66] & b[73])^(a[65] & b[74])^(a[64] & b[75])^(a[63] & b[76])^(a[62] & b[77])^(a[61] & b[78])^(a[60] & b[79])^(a[59] & b[80])^(a[58] & b[81])^(a[57] & b[82])^(a[56] & b[83])^(a[55] & b[84])^(a[54] & b[85])^(a[53] & b[86])^(a[52] & b[87])^(a[51] & b[88])^(a[50] & b[89])^(a[49] & b[90])^(a[48] & b[91])^(a[47] & b[92])^(a[46] & b[93])^(a[45] & b[94])^(a[44] & b[95])^(a[43] & b[96])^(a[42] & b[97])^(a[41] & b[98])^(a[40] & b[99])^(a[39] & b[100])^(a[38] & b[101])^(a[37] & b[102])^(a[36] & b[103])^(a[35] & b[104])^(a[34] & b[105])^(a[33] & b[106])^(a[32] & b[107])^(a[31] & b[108])^(a[30] & b[109])^(a[29] & b[110])^(a[28] & b[111])^(a[27] & b[112])^(a[26] & b[113])^(a[25] & b[114])^(a[24] & b[115])^(a[23] & b[116])^(a[22] & b[117])^(a[21] & b[118])^(a[20] & b[119])^(a[19] & b[120])^(a[18] & b[121])^(a[17] & b[122])^(a[16] & b[123])^(a[15] & b[124])^(a[14] & b[125])^(a[13] & b[126])^(a[12] & b[127])^(a[11] & b[128])^(a[10] & b[129])^(a[9] & b[130])^(a[8] & b[131])^(a[7] & b[132])^(a[6] & b[133])^(a[5] & b[134])^(a[4] & b[135])^(a[3] & b[136])^(a[2] & b[137])^(a[1] & b[138])^(a[0] & b[139]);
assign y[140] = (a[140] & b[0])^(a[139] & b[1])^(a[138] & b[2])^(a[137] & b[3])^(a[136] & b[4])^(a[135] & b[5])^(a[134] & b[6])^(a[133] & b[7])^(a[132] & b[8])^(a[131] & b[9])^(a[130] & b[10])^(a[129] & b[11])^(a[128] & b[12])^(a[127] & b[13])^(a[126] & b[14])^(a[125] & b[15])^(a[124] & b[16])^(a[123] & b[17])^(a[122] & b[18])^(a[121] & b[19])^(a[120] & b[20])^(a[119] & b[21])^(a[118] & b[22])^(a[117] & b[23])^(a[116] & b[24])^(a[115] & b[25])^(a[114] & b[26])^(a[113] & b[27])^(a[112] & b[28])^(a[111] & b[29])^(a[110] & b[30])^(a[109] & b[31])^(a[108] & b[32])^(a[107] & b[33])^(a[106] & b[34])^(a[105] & b[35])^(a[104] & b[36])^(a[103] & b[37])^(a[102] & b[38])^(a[101] & b[39])^(a[100] & b[40])^(a[99] & b[41])^(a[98] & b[42])^(a[97] & b[43])^(a[96] & b[44])^(a[95] & b[45])^(a[94] & b[46])^(a[93] & b[47])^(a[92] & b[48])^(a[91] & b[49])^(a[90] & b[50])^(a[89] & b[51])^(a[88] & b[52])^(a[87] & b[53])^(a[86] & b[54])^(a[85] & b[55])^(a[84] & b[56])^(a[83] & b[57])^(a[82] & b[58])^(a[81] & b[59])^(a[80] & b[60])^(a[79] & b[61])^(a[78] & b[62])^(a[77] & b[63])^(a[76] & b[64])^(a[75] & b[65])^(a[74] & b[66])^(a[73] & b[67])^(a[72] & b[68])^(a[71] & b[69])^(a[70] & b[70])^(a[69] & b[71])^(a[68] & b[72])^(a[67] & b[73])^(a[66] & b[74])^(a[65] & b[75])^(a[64] & b[76])^(a[63] & b[77])^(a[62] & b[78])^(a[61] & b[79])^(a[60] & b[80])^(a[59] & b[81])^(a[58] & b[82])^(a[57] & b[83])^(a[56] & b[84])^(a[55] & b[85])^(a[54] & b[86])^(a[53] & b[87])^(a[52] & b[88])^(a[51] & b[89])^(a[50] & b[90])^(a[49] & b[91])^(a[48] & b[92])^(a[47] & b[93])^(a[46] & b[94])^(a[45] & b[95])^(a[44] & b[96])^(a[43] & b[97])^(a[42] & b[98])^(a[41] & b[99])^(a[40] & b[100])^(a[39] & b[101])^(a[38] & b[102])^(a[37] & b[103])^(a[36] & b[104])^(a[35] & b[105])^(a[34] & b[106])^(a[33] & b[107])^(a[32] & b[108])^(a[31] & b[109])^(a[30] & b[110])^(a[29] & b[111])^(a[28] & b[112])^(a[27] & b[113])^(a[26] & b[114])^(a[25] & b[115])^(a[24] & b[116])^(a[23] & b[117])^(a[22] & b[118])^(a[21] & b[119])^(a[20] & b[120])^(a[19] & b[121])^(a[18] & b[122])^(a[17] & b[123])^(a[16] & b[124])^(a[15] & b[125])^(a[14] & b[126])^(a[13] & b[127])^(a[12] & b[128])^(a[11] & b[129])^(a[10] & b[130])^(a[9] & b[131])^(a[8] & b[132])^(a[7] & b[133])^(a[6] & b[134])^(a[5] & b[135])^(a[4] & b[136])^(a[3] & b[137])^(a[2] & b[138])^(a[1] & b[139])^(a[0] & b[140]);
assign y[141] = (a[141] & b[0])^(a[140] & b[1])^(a[139] & b[2])^(a[138] & b[3])^(a[137] & b[4])^(a[136] & b[5])^(a[135] & b[6])^(a[134] & b[7])^(a[133] & b[8])^(a[132] & b[9])^(a[131] & b[10])^(a[130] & b[11])^(a[129] & b[12])^(a[128] & b[13])^(a[127] & b[14])^(a[126] & b[15])^(a[125] & b[16])^(a[124] & b[17])^(a[123] & b[18])^(a[122] & b[19])^(a[121] & b[20])^(a[120] & b[21])^(a[119] & b[22])^(a[118] & b[23])^(a[117] & b[24])^(a[116] & b[25])^(a[115] & b[26])^(a[114] & b[27])^(a[113] & b[28])^(a[112] & b[29])^(a[111] & b[30])^(a[110] & b[31])^(a[109] & b[32])^(a[108] & b[33])^(a[107] & b[34])^(a[106] & b[35])^(a[105] & b[36])^(a[104] & b[37])^(a[103] & b[38])^(a[102] & b[39])^(a[101] & b[40])^(a[100] & b[41])^(a[99] & b[42])^(a[98] & b[43])^(a[97] & b[44])^(a[96] & b[45])^(a[95] & b[46])^(a[94] & b[47])^(a[93] & b[48])^(a[92] & b[49])^(a[91] & b[50])^(a[90] & b[51])^(a[89] & b[52])^(a[88] & b[53])^(a[87] & b[54])^(a[86] & b[55])^(a[85] & b[56])^(a[84] & b[57])^(a[83] & b[58])^(a[82] & b[59])^(a[81] & b[60])^(a[80] & b[61])^(a[79] & b[62])^(a[78] & b[63])^(a[77] & b[64])^(a[76] & b[65])^(a[75] & b[66])^(a[74] & b[67])^(a[73] & b[68])^(a[72] & b[69])^(a[71] & b[70])^(a[70] & b[71])^(a[69] & b[72])^(a[68] & b[73])^(a[67] & b[74])^(a[66] & b[75])^(a[65] & b[76])^(a[64] & b[77])^(a[63] & b[78])^(a[62] & b[79])^(a[61] & b[80])^(a[60] & b[81])^(a[59] & b[82])^(a[58] & b[83])^(a[57] & b[84])^(a[56] & b[85])^(a[55] & b[86])^(a[54] & b[87])^(a[53] & b[88])^(a[52] & b[89])^(a[51] & b[90])^(a[50] & b[91])^(a[49] & b[92])^(a[48] & b[93])^(a[47] & b[94])^(a[46] & b[95])^(a[45] & b[96])^(a[44] & b[97])^(a[43] & b[98])^(a[42] & b[99])^(a[41] & b[100])^(a[40] & b[101])^(a[39] & b[102])^(a[38] & b[103])^(a[37] & b[104])^(a[36] & b[105])^(a[35] & b[106])^(a[34] & b[107])^(a[33] & b[108])^(a[32] & b[109])^(a[31] & b[110])^(a[30] & b[111])^(a[29] & b[112])^(a[28] & b[113])^(a[27] & b[114])^(a[26] & b[115])^(a[25] & b[116])^(a[24] & b[117])^(a[23] & b[118])^(a[22] & b[119])^(a[21] & b[120])^(a[20] & b[121])^(a[19] & b[122])^(a[18] & b[123])^(a[17] & b[124])^(a[16] & b[125])^(a[15] & b[126])^(a[14] & b[127])^(a[13] & b[128])^(a[12] & b[129])^(a[11] & b[130])^(a[10] & b[131])^(a[9] & b[132])^(a[8] & b[133])^(a[7] & b[134])^(a[6] & b[135])^(a[5] & b[136])^(a[4] & b[137])^(a[3] & b[138])^(a[2] & b[139])^(a[1] & b[140])^(a[0] & b[141]);
assign y[142] = (a[142] & b[0])^(a[141] & b[1])^(a[140] & b[2])^(a[139] & b[3])^(a[138] & b[4])^(a[137] & b[5])^(a[136] & b[6])^(a[135] & b[7])^(a[134] & b[8])^(a[133] & b[9])^(a[132] & b[10])^(a[131] & b[11])^(a[130] & b[12])^(a[129] & b[13])^(a[128] & b[14])^(a[127] & b[15])^(a[126] & b[16])^(a[125] & b[17])^(a[124] & b[18])^(a[123] & b[19])^(a[122] & b[20])^(a[121] & b[21])^(a[120] & b[22])^(a[119] & b[23])^(a[118] & b[24])^(a[117] & b[25])^(a[116] & b[26])^(a[115] & b[27])^(a[114] & b[28])^(a[113] & b[29])^(a[112] & b[30])^(a[111] & b[31])^(a[110] & b[32])^(a[109] & b[33])^(a[108] & b[34])^(a[107] & b[35])^(a[106] & b[36])^(a[105] & b[37])^(a[104] & b[38])^(a[103] & b[39])^(a[102] & b[40])^(a[101] & b[41])^(a[100] & b[42])^(a[99] & b[43])^(a[98] & b[44])^(a[97] & b[45])^(a[96] & b[46])^(a[95] & b[47])^(a[94] & b[48])^(a[93] & b[49])^(a[92] & b[50])^(a[91] & b[51])^(a[90] & b[52])^(a[89] & b[53])^(a[88] & b[54])^(a[87] & b[55])^(a[86] & b[56])^(a[85] & b[57])^(a[84] & b[58])^(a[83] & b[59])^(a[82] & b[60])^(a[81] & b[61])^(a[80] & b[62])^(a[79] & b[63])^(a[78] & b[64])^(a[77] & b[65])^(a[76] & b[66])^(a[75] & b[67])^(a[74] & b[68])^(a[73] & b[69])^(a[72] & b[70])^(a[71] & b[71])^(a[70] & b[72])^(a[69] & b[73])^(a[68] & b[74])^(a[67] & b[75])^(a[66] & b[76])^(a[65] & b[77])^(a[64] & b[78])^(a[63] & b[79])^(a[62] & b[80])^(a[61] & b[81])^(a[60] & b[82])^(a[59] & b[83])^(a[58] & b[84])^(a[57] & b[85])^(a[56] & b[86])^(a[55] & b[87])^(a[54] & b[88])^(a[53] & b[89])^(a[52] & b[90])^(a[51] & b[91])^(a[50] & b[92])^(a[49] & b[93])^(a[48] & b[94])^(a[47] & b[95])^(a[46] & b[96])^(a[45] & b[97])^(a[44] & b[98])^(a[43] & b[99])^(a[42] & b[100])^(a[41] & b[101])^(a[40] & b[102])^(a[39] & b[103])^(a[38] & b[104])^(a[37] & b[105])^(a[36] & b[106])^(a[35] & b[107])^(a[34] & b[108])^(a[33] & b[109])^(a[32] & b[110])^(a[31] & b[111])^(a[30] & b[112])^(a[29] & b[113])^(a[28] & b[114])^(a[27] & b[115])^(a[26] & b[116])^(a[25] & b[117])^(a[24] & b[118])^(a[23] & b[119])^(a[22] & b[120])^(a[21] & b[121])^(a[20] & b[122])^(a[19] & b[123])^(a[18] & b[124])^(a[17] & b[125])^(a[16] & b[126])^(a[15] & b[127])^(a[14] & b[128])^(a[13] & b[129])^(a[12] & b[130])^(a[11] & b[131])^(a[10] & b[132])^(a[9] & b[133])^(a[8] & b[134])^(a[7] & b[135])^(a[6] & b[136])^(a[5] & b[137])^(a[4] & b[138])^(a[3] & b[139])^(a[2] & b[140])^(a[1] & b[141])^(a[0] & b[142]);
assign y[143] = (a[143] & b[0])^(a[142] & b[1])^(a[141] & b[2])^(a[140] & b[3])^(a[139] & b[4])^(a[138] & b[5])^(a[137] & b[6])^(a[136] & b[7])^(a[135] & b[8])^(a[134] & b[9])^(a[133] & b[10])^(a[132] & b[11])^(a[131] & b[12])^(a[130] & b[13])^(a[129] & b[14])^(a[128] & b[15])^(a[127] & b[16])^(a[126] & b[17])^(a[125] & b[18])^(a[124] & b[19])^(a[123] & b[20])^(a[122] & b[21])^(a[121] & b[22])^(a[120] & b[23])^(a[119] & b[24])^(a[118] & b[25])^(a[117] & b[26])^(a[116] & b[27])^(a[115] & b[28])^(a[114] & b[29])^(a[113] & b[30])^(a[112] & b[31])^(a[111] & b[32])^(a[110] & b[33])^(a[109] & b[34])^(a[108] & b[35])^(a[107] & b[36])^(a[106] & b[37])^(a[105] & b[38])^(a[104] & b[39])^(a[103] & b[40])^(a[102] & b[41])^(a[101] & b[42])^(a[100] & b[43])^(a[99] & b[44])^(a[98] & b[45])^(a[97] & b[46])^(a[96] & b[47])^(a[95] & b[48])^(a[94] & b[49])^(a[93] & b[50])^(a[92] & b[51])^(a[91] & b[52])^(a[90] & b[53])^(a[89] & b[54])^(a[88] & b[55])^(a[87] & b[56])^(a[86] & b[57])^(a[85] & b[58])^(a[84] & b[59])^(a[83] & b[60])^(a[82] & b[61])^(a[81] & b[62])^(a[80] & b[63])^(a[79] & b[64])^(a[78] & b[65])^(a[77] & b[66])^(a[76] & b[67])^(a[75] & b[68])^(a[74] & b[69])^(a[73] & b[70])^(a[72] & b[71])^(a[71] & b[72])^(a[70] & b[73])^(a[69] & b[74])^(a[68] & b[75])^(a[67] & b[76])^(a[66] & b[77])^(a[65] & b[78])^(a[64] & b[79])^(a[63] & b[80])^(a[62] & b[81])^(a[61] & b[82])^(a[60] & b[83])^(a[59] & b[84])^(a[58] & b[85])^(a[57] & b[86])^(a[56] & b[87])^(a[55] & b[88])^(a[54] & b[89])^(a[53] & b[90])^(a[52] & b[91])^(a[51] & b[92])^(a[50] & b[93])^(a[49] & b[94])^(a[48] & b[95])^(a[47] & b[96])^(a[46] & b[97])^(a[45] & b[98])^(a[44] & b[99])^(a[43] & b[100])^(a[42] & b[101])^(a[41] & b[102])^(a[40] & b[103])^(a[39] & b[104])^(a[38] & b[105])^(a[37] & b[106])^(a[36] & b[107])^(a[35] & b[108])^(a[34] & b[109])^(a[33] & b[110])^(a[32] & b[111])^(a[31] & b[112])^(a[30] & b[113])^(a[29] & b[114])^(a[28] & b[115])^(a[27] & b[116])^(a[26] & b[117])^(a[25] & b[118])^(a[24] & b[119])^(a[23] & b[120])^(a[22] & b[121])^(a[21] & b[122])^(a[20] & b[123])^(a[19] & b[124])^(a[18] & b[125])^(a[17] & b[126])^(a[16] & b[127])^(a[15] & b[128])^(a[14] & b[129])^(a[13] & b[130])^(a[12] & b[131])^(a[11] & b[132])^(a[10] & b[133])^(a[9] & b[134])^(a[8] & b[135])^(a[7] & b[136])^(a[6] & b[137])^(a[5] & b[138])^(a[4] & b[139])^(a[3] & b[140])^(a[2] & b[141])^(a[1] & b[142])^(a[0] & b[143]);
assign y[144] = (a[144] & b[0])^(a[143] & b[1])^(a[142] & b[2])^(a[141] & b[3])^(a[140] & b[4])^(a[139] & b[5])^(a[138] & b[6])^(a[137] & b[7])^(a[136] & b[8])^(a[135] & b[9])^(a[134] & b[10])^(a[133] & b[11])^(a[132] & b[12])^(a[131] & b[13])^(a[130] & b[14])^(a[129] & b[15])^(a[128] & b[16])^(a[127] & b[17])^(a[126] & b[18])^(a[125] & b[19])^(a[124] & b[20])^(a[123] & b[21])^(a[122] & b[22])^(a[121] & b[23])^(a[120] & b[24])^(a[119] & b[25])^(a[118] & b[26])^(a[117] & b[27])^(a[116] & b[28])^(a[115] & b[29])^(a[114] & b[30])^(a[113] & b[31])^(a[112] & b[32])^(a[111] & b[33])^(a[110] & b[34])^(a[109] & b[35])^(a[108] & b[36])^(a[107] & b[37])^(a[106] & b[38])^(a[105] & b[39])^(a[104] & b[40])^(a[103] & b[41])^(a[102] & b[42])^(a[101] & b[43])^(a[100] & b[44])^(a[99] & b[45])^(a[98] & b[46])^(a[97] & b[47])^(a[96] & b[48])^(a[95] & b[49])^(a[94] & b[50])^(a[93] & b[51])^(a[92] & b[52])^(a[91] & b[53])^(a[90] & b[54])^(a[89] & b[55])^(a[88] & b[56])^(a[87] & b[57])^(a[86] & b[58])^(a[85] & b[59])^(a[84] & b[60])^(a[83] & b[61])^(a[82] & b[62])^(a[81] & b[63])^(a[80] & b[64])^(a[79] & b[65])^(a[78] & b[66])^(a[77] & b[67])^(a[76] & b[68])^(a[75] & b[69])^(a[74] & b[70])^(a[73] & b[71])^(a[72] & b[72])^(a[71] & b[73])^(a[70] & b[74])^(a[69] & b[75])^(a[68] & b[76])^(a[67] & b[77])^(a[66] & b[78])^(a[65] & b[79])^(a[64] & b[80])^(a[63] & b[81])^(a[62] & b[82])^(a[61] & b[83])^(a[60] & b[84])^(a[59] & b[85])^(a[58] & b[86])^(a[57] & b[87])^(a[56] & b[88])^(a[55] & b[89])^(a[54] & b[90])^(a[53] & b[91])^(a[52] & b[92])^(a[51] & b[93])^(a[50] & b[94])^(a[49] & b[95])^(a[48] & b[96])^(a[47] & b[97])^(a[46] & b[98])^(a[45] & b[99])^(a[44] & b[100])^(a[43] & b[101])^(a[42] & b[102])^(a[41] & b[103])^(a[40] & b[104])^(a[39] & b[105])^(a[38] & b[106])^(a[37] & b[107])^(a[36] & b[108])^(a[35] & b[109])^(a[34] & b[110])^(a[33] & b[111])^(a[32] & b[112])^(a[31] & b[113])^(a[30] & b[114])^(a[29] & b[115])^(a[28] & b[116])^(a[27] & b[117])^(a[26] & b[118])^(a[25] & b[119])^(a[24] & b[120])^(a[23] & b[121])^(a[22] & b[122])^(a[21] & b[123])^(a[20] & b[124])^(a[19] & b[125])^(a[18] & b[126])^(a[17] & b[127])^(a[16] & b[128])^(a[15] & b[129])^(a[14] & b[130])^(a[13] & b[131])^(a[12] & b[132])^(a[11] & b[133])^(a[10] & b[134])^(a[9] & b[135])^(a[8] & b[136])^(a[7] & b[137])^(a[6] & b[138])^(a[5] & b[139])^(a[4] & b[140])^(a[3] & b[141])^(a[2] & b[142])^(a[1] & b[143])^(a[0] & b[144]);
assign y[145] = (a[145] & b[0])^(a[144] & b[1])^(a[143] & b[2])^(a[142] & b[3])^(a[141] & b[4])^(a[140] & b[5])^(a[139] & b[6])^(a[138] & b[7])^(a[137] & b[8])^(a[136] & b[9])^(a[135] & b[10])^(a[134] & b[11])^(a[133] & b[12])^(a[132] & b[13])^(a[131] & b[14])^(a[130] & b[15])^(a[129] & b[16])^(a[128] & b[17])^(a[127] & b[18])^(a[126] & b[19])^(a[125] & b[20])^(a[124] & b[21])^(a[123] & b[22])^(a[122] & b[23])^(a[121] & b[24])^(a[120] & b[25])^(a[119] & b[26])^(a[118] & b[27])^(a[117] & b[28])^(a[116] & b[29])^(a[115] & b[30])^(a[114] & b[31])^(a[113] & b[32])^(a[112] & b[33])^(a[111] & b[34])^(a[110] & b[35])^(a[109] & b[36])^(a[108] & b[37])^(a[107] & b[38])^(a[106] & b[39])^(a[105] & b[40])^(a[104] & b[41])^(a[103] & b[42])^(a[102] & b[43])^(a[101] & b[44])^(a[100] & b[45])^(a[99] & b[46])^(a[98] & b[47])^(a[97] & b[48])^(a[96] & b[49])^(a[95] & b[50])^(a[94] & b[51])^(a[93] & b[52])^(a[92] & b[53])^(a[91] & b[54])^(a[90] & b[55])^(a[89] & b[56])^(a[88] & b[57])^(a[87] & b[58])^(a[86] & b[59])^(a[85] & b[60])^(a[84] & b[61])^(a[83] & b[62])^(a[82] & b[63])^(a[81] & b[64])^(a[80] & b[65])^(a[79] & b[66])^(a[78] & b[67])^(a[77] & b[68])^(a[76] & b[69])^(a[75] & b[70])^(a[74] & b[71])^(a[73] & b[72])^(a[72] & b[73])^(a[71] & b[74])^(a[70] & b[75])^(a[69] & b[76])^(a[68] & b[77])^(a[67] & b[78])^(a[66] & b[79])^(a[65] & b[80])^(a[64] & b[81])^(a[63] & b[82])^(a[62] & b[83])^(a[61] & b[84])^(a[60] & b[85])^(a[59] & b[86])^(a[58] & b[87])^(a[57] & b[88])^(a[56] & b[89])^(a[55] & b[90])^(a[54] & b[91])^(a[53] & b[92])^(a[52] & b[93])^(a[51] & b[94])^(a[50] & b[95])^(a[49] & b[96])^(a[48] & b[97])^(a[47] & b[98])^(a[46] & b[99])^(a[45] & b[100])^(a[44] & b[101])^(a[43] & b[102])^(a[42] & b[103])^(a[41] & b[104])^(a[40] & b[105])^(a[39] & b[106])^(a[38] & b[107])^(a[37] & b[108])^(a[36] & b[109])^(a[35] & b[110])^(a[34] & b[111])^(a[33] & b[112])^(a[32] & b[113])^(a[31] & b[114])^(a[30] & b[115])^(a[29] & b[116])^(a[28] & b[117])^(a[27] & b[118])^(a[26] & b[119])^(a[25] & b[120])^(a[24] & b[121])^(a[23] & b[122])^(a[22] & b[123])^(a[21] & b[124])^(a[20] & b[125])^(a[19] & b[126])^(a[18] & b[127])^(a[17] & b[128])^(a[16] & b[129])^(a[15] & b[130])^(a[14] & b[131])^(a[13] & b[132])^(a[12] & b[133])^(a[11] & b[134])^(a[10] & b[135])^(a[9] & b[136])^(a[8] & b[137])^(a[7] & b[138])^(a[6] & b[139])^(a[5] & b[140])^(a[4] & b[141])^(a[3] & b[142])^(a[2] & b[143])^(a[1] & b[144])^(a[0] & b[145]);
assign y[146] = (a[146] & b[0])^(a[145] & b[1])^(a[144] & b[2])^(a[143] & b[3])^(a[142] & b[4])^(a[141] & b[5])^(a[140] & b[6])^(a[139] & b[7])^(a[138] & b[8])^(a[137] & b[9])^(a[136] & b[10])^(a[135] & b[11])^(a[134] & b[12])^(a[133] & b[13])^(a[132] & b[14])^(a[131] & b[15])^(a[130] & b[16])^(a[129] & b[17])^(a[128] & b[18])^(a[127] & b[19])^(a[126] & b[20])^(a[125] & b[21])^(a[124] & b[22])^(a[123] & b[23])^(a[122] & b[24])^(a[121] & b[25])^(a[120] & b[26])^(a[119] & b[27])^(a[118] & b[28])^(a[117] & b[29])^(a[116] & b[30])^(a[115] & b[31])^(a[114] & b[32])^(a[113] & b[33])^(a[112] & b[34])^(a[111] & b[35])^(a[110] & b[36])^(a[109] & b[37])^(a[108] & b[38])^(a[107] & b[39])^(a[106] & b[40])^(a[105] & b[41])^(a[104] & b[42])^(a[103] & b[43])^(a[102] & b[44])^(a[101] & b[45])^(a[100] & b[46])^(a[99] & b[47])^(a[98] & b[48])^(a[97] & b[49])^(a[96] & b[50])^(a[95] & b[51])^(a[94] & b[52])^(a[93] & b[53])^(a[92] & b[54])^(a[91] & b[55])^(a[90] & b[56])^(a[89] & b[57])^(a[88] & b[58])^(a[87] & b[59])^(a[86] & b[60])^(a[85] & b[61])^(a[84] & b[62])^(a[83] & b[63])^(a[82] & b[64])^(a[81] & b[65])^(a[80] & b[66])^(a[79] & b[67])^(a[78] & b[68])^(a[77] & b[69])^(a[76] & b[70])^(a[75] & b[71])^(a[74] & b[72])^(a[73] & b[73])^(a[72] & b[74])^(a[71] & b[75])^(a[70] & b[76])^(a[69] & b[77])^(a[68] & b[78])^(a[67] & b[79])^(a[66] & b[80])^(a[65] & b[81])^(a[64] & b[82])^(a[63] & b[83])^(a[62] & b[84])^(a[61] & b[85])^(a[60] & b[86])^(a[59] & b[87])^(a[58] & b[88])^(a[57] & b[89])^(a[56] & b[90])^(a[55] & b[91])^(a[54] & b[92])^(a[53] & b[93])^(a[52] & b[94])^(a[51] & b[95])^(a[50] & b[96])^(a[49] & b[97])^(a[48] & b[98])^(a[47] & b[99])^(a[46] & b[100])^(a[45] & b[101])^(a[44] & b[102])^(a[43] & b[103])^(a[42] & b[104])^(a[41] & b[105])^(a[40] & b[106])^(a[39] & b[107])^(a[38] & b[108])^(a[37] & b[109])^(a[36] & b[110])^(a[35] & b[111])^(a[34] & b[112])^(a[33] & b[113])^(a[32] & b[114])^(a[31] & b[115])^(a[30] & b[116])^(a[29] & b[117])^(a[28] & b[118])^(a[27] & b[119])^(a[26] & b[120])^(a[25] & b[121])^(a[24] & b[122])^(a[23] & b[123])^(a[22] & b[124])^(a[21] & b[125])^(a[20] & b[126])^(a[19] & b[127])^(a[18] & b[128])^(a[17] & b[129])^(a[16] & b[130])^(a[15] & b[131])^(a[14] & b[132])^(a[13] & b[133])^(a[12] & b[134])^(a[11] & b[135])^(a[10] & b[136])^(a[9] & b[137])^(a[8] & b[138])^(a[7] & b[139])^(a[6] & b[140])^(a[5] & b[141])^(a[4] & b[142])^(a[3] & b[143])^(a[2] & b[144])^(a[1] & b[145])^(a[0] & b[146]);
assign y[147] = (a[147] & b[0])^(a[146] & b[1])^(a[145] & b[2])^(a[144] & b[3])^(a[143] & b[4])^(a[142] & b[5])^(a[141] & b[6])^(a[140] & b[7])^(a[139] & b[8])^(a[138] & b[9])^(a[137] & b[10])^(a[136] & b[11])^(a[135] & b[12])^(a[134] & b[13])^(a[133] & b[14])^(a[132] & b[15])^(a[131] & b[16])^(a[130] & b[17])^(a[129] & b[18])^(a[128] & b[19])^(a[127] & b[20])^(a[126] & b[21])^(a[125] & b[22])^(a[124] & b[23])^(a[123] & b[24])^(a[122] & b[25])^(a[121] & b[26])^(a[120] & b[27])^(a[119] & b[28])^(a[118] & b[29])^(a[117] & b[30])^(a[116] & b[31])^(a[115] & b[32])^(a[114] & b[33])^(a[113] & b[34])^(a[112] & b[35])^(a[111] & b[36])^(a[110] & b[37])^(a[109] & b[38])^(a[108] & b[39])^(a[107] & b[40])^(a[106] & b[41])^(a[105] & b[42])^(a[104] & b[43])^(a[103] & b[44])^(a[102] & b[45])^(a[101] & b[46])^(a[100] & b[47])^(a[99] & b[48])^(a[98] & b[49])^(a[97] & b[50])^(a[96] & b[51])^(a[95] & b[52])^(a[94] & b[53])^(a[93] & b[54])^(a[92] & b[55])^(a[91] & b[56])^(a[90] & b[57])^(a[89] & b[58])^(a[88] & b[59])^(a[87] & b[60])^(a[86] & b[61])^(a[85] & b[62])^(a[84] & b[63])^(a[83] & b[64])^(a[82] & b[65])^(a[81] & b[66])^(a[80] & b[67])^(a[79] & b[68])^(a[78] & b[69])^(a[77] & b[70])^(a[76] & b[71])^(a[75] & b[72])^(a[74] & b[73])^(a[73] & b[74])^(a[72] & b[75])^(a[71] & b[76])^(a[70] & b[77])^(a[69] & b[78])^(a[68] & b[79])^(a[67] & b[80])^(a[66] & b[81])^(a[65] & b[82])^(a[64] & b[83])^(a[63] & b[84])^(a[62] & b[85])^(a[61] & b[86])^(a[60] & b[87])^(a[59] & b[88])^(a[58] & b[89])^(a[57] & b[90])^(a[56] & b[91])^(a[55] & b[92])^(a[54] & b[93])^(a[53] & b[94])^(a[52] & b[95])^(a[51] & b[96])^(a[50] & b[97])^(a[49] & b[98])^(a[48] & b[99])^(a[47] & b[100])^(a[46] & b[101])^(a[45] & b[102])^(a[44] & b[103])^(a[43] & b[104])^(a[42] & b[105])^(a[41] & b[106])^(a[40] & b[107])^(a[39] & b[108])^(a[38] & b[109])^(a[37] & b[110])^(a[36] & b[111])^(a[35] & b[112])^(a[34] & b[113])^(a[33] & b[114])^(a[32] & b[115])^(a[31] & b[116])^(a[30] & b[117])^(a[29] & b[118])^(a[28] & b[119])^(a[27] & b[120])^(a[26] & b[121])^(a[25] & b[122])^(a[24] & b[123])^(a[23] & b[124])^(a[22] & b[125])^(a[21] & b[126])^(a[20] & b[127])^(a[19] & b[128])^(a[18] & b[129])^(a[17] & b[130])^(a[16] & b[131])^(a[15] & b[132])^(a[14] & b[133])^(a[13] & b[134])^(a[12] & b[135])^(a[11] & b[136])^(a[10] & b[137])^(a[9] & b[138])^(a[8] & b[139])^(a[7] & b[140])^(a[6] & b[141])^(a[5] & b[142])^(a[4] & b[143])^(a[3] & b[144])^(a[2] & b[145])^(a[1] & b[146])^(a[0] & b[147]);
assign y[148] = (a[148] & b[0])^(a[147] & b[1])^(a[146] & b[2])^(a[145] & b[3])^(a[144] & b[4])^(a[143] & b[5])^(a[142] & b[6])^(a[141] & b[7])^(a[140] & b[8])^(a[139] & b[9])^(a[138] & b[10])^(a[137] & b[11])^(a[136] & b[12])^(a[135] & b[13])^(a[134] & b[14])^(a[133] & b[15])^(a[132] & b[16])^(a[131] & b[17])^(a[130] & b[18])^(a[129] & b[19])^(a[128] & b[20])^(a[127] & b[21])^(a[126] & b[22])^(a[125] & b[23])^(a[124] & b[24])^(a[123] & b[25])^(a[122] & b[26])^(a[121] & b[27])^(a[120] & b[28])^(a[119] & b[29])^(a[118] & b[30])^(a[117] & b[31])^(a[116] & b[32])^(a[115] & b[33])^(a[114] & b[34])^(a[113] & b[35])^(a[112] & b[36])^(a[111] & b[37])^(a[110] & b[38])^(a[109] & b[39])^(a[108] & b[40])^(a[107] & b[41])^(a[106] & b[42])^(a[105] & b[43])^(a[104] & b[44])^(a[103] & b[45])^(a[102] & b[46])^(a[101] & b[47])^(a[100] & b[48])^(a[99] & b[49])^(a[98] & b[50])^(a[97] & b[51])^(a[96] & b[52])^(a[95] & b[53])^(a[94] & b[54])^(a[93] & b[55])^(a[92] & b[56])^(a[91] & b[57])^(a[90] & b[58])^(a[89] & b[59])^(a[88] & b[60])^(a[87] & b[61])^(a[86] & b[62])^(a[85] & b[63])^(a[84] & b[64])^(a[83] & b[65])^(a[82] & b[66])^(a[81] & b[67])^(a[80] & b[68])^(a[79] & b[69])^(a[78] & b[70])^(a[77] & b[71])^(a[76] & b[72])^(a[75] & b[73])^(a[74] & b[74])^(a[73] & b[75])^(a[72] & b[76])^(a[71] & b[77])^(a[70] & b[78])^(a[69] & b[79])^(a[68] & b[80])^(a[67] & b[81])^(a[66] & b[82])^(a[65] & b[83])^(a[64] & b[84])^(a[63] & b[85])^(a[62] & b[86])^(a[61] & b[87])^(a[60] & b[88])^(a[59] & b[89])^(a[58] & b[90])^(a[57] & b[91])^(a[56] & b[92])^(a[55] & b[93])^(a[54] & b[94])^(a[53] & b[95])^(a[52] & b[96])^(a[51] & b[97])^(a[50] & b[98])^(a[49] & b[99])^(a[48] & b[100])^(a[47] & b[101])^(a[46] & b[102])^(a[45] & b[103])^(a[44] & b[104])^(a[43] & b[105])^(a[42] & b[106])^(a[41] & b[107])^(a[40] & b[108])^(a[39] & b[109])^(a[38] & b[110])^(a[37] & b[111])^(a[36] & b[112])^(a[35] & b[113])^(a[34] & b[114])^(a[33] & b[115])^(a[32] & b[116])^(a[31] & b[117])^(a[30] & b[118])^(a[29] & b[119])^(a[28] & b[120])^(a[27] & b[121])^(a[26] & b[122])^(a[25] & b[123])^(a[24] & b[124])^(a[23] & b[125])^(a[22] & b[126])^(a[21] & b[127])^(a[20] & b[128])^(a[19] & b[129])^(a[18] & b[130])^(a[17] & b[131])^(a[16] & b[132])^(a[15] & b[133])^(a[14] & b[134])^(a[13] & b[135])^(a[12] & b[136])^(a[11] & b[137])^(a[10] & b[138])^(a[9] & b[139])^(a[8] & b[140])^(a[7] & b[141])^(a[6] & b[142])^(a[5] & b[143])^(a[4] & b[144])^(a[3] & b[145])^(a[2] & b[146])^(a[1] & b[147])^(a[0] & b[148]);
assign y[149] = (a[149] & b[0])^(a[148] & b[1])^(a[147] & b[2])^(a[146] & b[3])^(a[145] & b[4])^(a[144] & b[5])^(a[143] & b[6])^(a[142] & b[7])^(a[141] & b[8])^(a[140] & b[9])^(a[139] & b[10])^(a[138] & b[11])^(a[137] & b[12])^(a[136] & b[13])^(a[135] & b[14])^(a[134] & b[15])^(a[133] & b[16])^(a[132] & b[17])^(a[131] & b[18])^(a[130] & b[19])^(a[129] & b[20])^(a[128] & b[21])^(a[127] & b[22])^(a[126] & b[23])^(a[125] & b[24])^(a[124] & b[25])^(a[123] & b[26])^(a[122] & b[27])^(a[121] & b[28])^(a[120] & b[29])^(a[119] & b[30])^(a[118] & b[31])^(a[117] & b[32])^(a[116] & b[33])^(a[115] & b[34])^(a[114] & b[35])^(a[113] & b[36])^(a[112] & b[37])^(a[111] & b[38])^(a[110] & b[39])^(a[109] & b[40])^(a[108] & b[41])^(a[107] & b[42])^(a[106] & b[43])^(a[105] & b[44])^(a[104] & b[45])^(a[103] & b[46])^(a[102] & b[47])^(a[101] & b[48])^(a[100] & b[49])^(a[99] & b[50])^(a[98] & b[51])^(a[97] & b[52])^(a[96] & b[53])^(a[95] & b[54])^(a[94] & b[55])^(a[93] & b[56])^(a[92] & b[57])^(a[91] & b[58])^(a[90] & b[59])^(a[89] & b[60])^(a[88] & b[61])^(a[87] & b[62])^(a[86] & b[63])^(a[85] & b[64])^(a[84] & b[65])^(a[83] & b[66])^(a[82] & b[67])^(a[81] & b[68])^(a[80] & b[69])^(a[79] & b[70])^(a[78] & b[71])^(a[77] & b[72])^(a[76] & b[73])^(a[75] & b[74])^(a[74] & b[75])^(a[73] & b[76])^(a[72] & b[77])^(a[71] & b[78])^(a[70] & b[79])^(a[69] & b[80])^(a[68] & b[81])^(a[67] & b[82])^(a[66] & b[83])^(a[65] & b[84])^(a[64] & b[85])^(a[63] & b[86])^(a[62] & b[87])^(a[61] & b[88])^(a[60] & b[89])^(a[59] & b[90])^(a[58] & b[91])^(a[57] & b[92])^(a[56] & b[93])^(a[55] & b[94])^(a[54] & b[95])^(a[53] & b[96])^(a[52] & b[97])^(a[51] & b[98])^(a[50] & b[99])^(a[49] & b[100])^(a[48] & b[101])^(a[47] & b[102])^(a[46] & b[103])^(a[45] & b[104])^(a[44] & b[105])^(a[43] & b[106])^(a[42] & b[107])^(a[41] & b[108])^(a[40] & b[109])^(a[39] & b[110])^(a[38] & b[111])^(a[37] & b[112])^(a[36] & b[113])^(a[35] & b[114])^(a[34] & b[115])^(a[33] & b[116])^(a[32] & b[117])^(a[31] & b[118])^(a[30] & b[119])^(a[29] & b[120])^(a[28] & b[121])^(a[27] & b[122])^(a[26] & b[123])^(a[25] & b[124])^(a[24] & b[125])^(a[23] & b[126])^(a[22] & b[127])^(a[21] & b[128])^(a[20] & b[129])^(a[19] & b[130])^(a[18] & b[131])^(a[17] & b[132])^(a[16] & b[133])^(a[15] & b[134])^(a[14] & b[135])^(a[13] & b[136])^(a[12] & b[137])^(a[11] & b[138])^(a[10] & b[139])^(a[9] & b[140])^(a[8] & b[141])^(a[7] & b[142])^(a[6] & b[143])^(a[5] & b[144])^(a[4] & b[145])^(a[3] & b[146])^(a[2] & b[147])^(a[1] & b[148])^(a[0] & b[149]);
assign y[150] = (a[150] & b[0])^(a[149] & b[1])^(a[148] & b[2])^(a[147] & b[3])^(a[146] & b[4])^(a[145] & b[5])^(a[144] & b[6])^(a[143] & b[7])^(a[142] & b[8])^(a[141] & b[9])^(a[140] & b[10])^(a[139] & b[11])^(a[138] & b[12])^(a[137] & b[13])^(a[136] & b[14])^(a[135] & b[15])^(a[134] & b[16])^(a[133] & b[17])^(a[132] & b[18])^(a[131] & b[19])^(a[130] & b[20])^(a[129] & b[21])^(a[128] & b[22])^(a[127] & b[23])^(a[126] & b[24])^(a[125] & b[25])^(a[124] & b[26])^(a[123] & b[27])^(a[122] & b[28])^(a[121] & b[29])^(a[120] & b[30])^(a[119] & b[31])^(a[118] & b[32])^(a[117] & b[33])^(a[116] & b[34])^(a[115] & b[35])^(a[114] & b[36])^(a[113] & b[37])^(a[112] & b[38])^(a[111] & b[39])^(a[110] & b[40])^(a[109] & b[41])^(a[108] & b[42])^(a[107] & b[43])^(a[106] & b[44])^(a[105] & b[45])^(a[104] & b[46])^(a[103] & b[47])^(a[102] & b[48])^(a[101] & b[49])^(a[100] & b[50])^(a[99] & b[51])^(a[98] & b[52])^(a[97] & b[53])^(a[96] & b[54])^(a[95] & b[55])^(a[94] & b[56])^(a[93] & b[57])^(a[92] & b[58])^(a[91] & b[59])^(a[90] & b[60])^(a[89] & b[61])^(a[88] & b[62])^(a[87] & b[63])^(a[86] & b[64])^(a[85] & b[65])^(a[84] & b[66])^(a[83] & b[67])^(a[82] & b[68])^(a[81] & b[69])^(a[80] & b[70])^(a[79] & b[71])^(a[78] & b[72])^(a[77] & b[73])^(a[76] & b[74])^(a[75] & b[75])^(a[74] & b[76])^(a[73] & b[77])^(a[72] & b[78])^(a[71] & b[79])^(a[70] & b[80])^(a[69] & b[81])^(a[68] & b[82])^(a[67] & b[83])^(a[66] & b[84])^(a[65] & b[85])^(a[64] & b[86])^(a[63] & b[87])^(a[62] & b[88])^(a[61] & b[89])^(a[60] & b[90])^(a[59] & b[91])^(a[58] & b[92])^(a[57] & b[93])^(a[56] & b[94])^(a[55] & b[95])^(a[54] & b[96])^(a[53] & b[97])^(a[52] & b[98])^(a[51] & b[99])^(a[50] & b[100])^(a[49] & b[101])^(a[48] & b[102])^(a[47] & b[103])^(a[46] & b[104])^(a[45] & b[105])^(a[44] & b[106])^(a[43] & b[107])^(a[42] & b[108])^(a[41] & b[109])^(a[40] & b[110])^(a[39] & b[111])^(a[38] & b[112])^(a[37] & b[113])^(a[36] & b[114])^(a[35] & b[115])^(a[34] & b[116])^(a[33] & b[117])^(a[32] & b[118])^(a[31] & b[119])^(a[30] & b[120])^(a[29] & b[121])^(a[28] & b[122])^(a[27] & b[123])^(a[26] & b[124])^(a[25] & b[125])^(a[24] & b[126])^(a[23] & b[127])^(a[22] & b[128])^(a[21] & b[129])^(a[20] & b[130])^(a[19] & b[131])^(a[18] & b[132])^(a[17] & b[133])^(a[16] & b[134])^(a[15] & b[135])^(a[14] & b[136])^(a[13] & b[137])^(a[12] & b[138])^(a[11] & b[139])^(a[10] & b[140])^(a[9] & b[141])^(a[8] & b[142])^(a[7] & b[143])^(a[6] & b[144])^(a[5] & b[145])^(a[4] & b[146])^(a[3] & b[147])^(a[2] & b[148])^(a[1] & b[149])^(a[0] & b[150]);
assign y[151] = (a[151] & b[0])^(a[150] & b[1])^(a[149] & b[2])^(a[148] & b[3])^(a[147] & b[4])^(a[146] & b[5])^(a[145] & b[6])^(a[144] & b[7])^(a[143] & b[8])^(a[142] & b[9])^(a[141] & b[10])^(a[140] & b[11])^(a[139] & b[12])^(a[138] & b[13])^(a[137] & b[14])^(a[136] & b[15])^(a[135] & b[16])^(a[134] & b[17])^(a[133] & b[18])^(a[132] & b[19])^(a[131] & b[20])^(a[130] & b[21])^(a[129] & b[22])^(a[128] & b[23])^(a[127] & b[24])^(a[126] & b[25])^(a[125] & b[26])^(a[124] & b[27])^(a[123] & b[28])^(a[122] & b[29])^(a[121] & b[30])^(a[120] & b[31])^(a[119] & b[32])^(a[118] & b[33])^(a[117] & b[34])^(a[116] & b[35])^(a[115] & b[36])^(a[114] & b[37])^(a[113] & b[38])^(a[112] & b[39])^(a[111] & b[40])^(a[110] & b[41])^(a[109] & b[42])^(a[108] & b[43])^(a[107] & b[44])^(a[106] & b[45])^(a[105] & b[46])^(a[104] & b[47])^(a[103] & b[48])^(a[102] & b[49])^(a[101] & b[50])^(a[100] & b[51])^(a[99] & b[52])^(a[98] & b[53])^(a[97] & b[54])^(a[96] & b[55])^(a[95] & b[56])^(a[94] & b[57])^(a[93] & b[58])^(a[92] & b[59])^(a[91] & b[60])^(a[90] & b[61])^(a[89] & b[62])^(a[88] & b[63])^(a[87] & b[64])^(a[86] & b[65])^(a[85] & b[66])^(a[84] & b[67])^(a[83] & b[68])^(a[82] & b[69])^(a[81] & b[70])^(a[80] & b[71])^(a[79] & b[72])^(a[78] & b[73])^(a[77] & b[74])^(a[76] & b[75])^(a[75] & b[76])^(a[74] & b[77])^(a[73] & b[78])^(a[72] & b[79])^(a[71] & b[80])^(a[70] & b[81])^(a[69] & b[82])^(a[68] & b[83])^(a[67] & b[84])^(a[66] & b[85])^(a[65] & b[86])^(a[64] & b[87])^(a[63] & b[88])^(a[62] & b[89])^(a[61] & b[90])^(a[60] & b[91])^(a[59] & b[92])^(a[58] & b[93])^(a[57] & b[94])^(a[56] & b[95])^(a[55] & b[96])^(a[54] & b[97])^(a[53] & b[98])^(a[52] & b[99])^(a[51] & b[100])^(a[50] & b[101])^(a[49] & b[102])^(a[48] & b[103])^(a[47] & b[104])^(a[46] & b[105])^(a[45] & b[106])^(a[44] & b[107])^(a[43] & b[108])^(a[42] & b[109])^(a[41] & b[110])^(a[40] & b[111])^(a[39] & b[112])^(a[38] & b[113])^(a[37] & b[114])^(a[36] & b[115])^(a[35] & b[116])^(a[34] & b[117])^(a[33] & b[118])^(a[32] & b[119])^(a[31] & b[120])^(a[30] & b[121])^(a[29] & b[122])^(a[28] & b[123])^(a[27] & b[124])^(a[26] & b[125])^(a[25] & b[126])^(a[24] & b[127])^(a[23] & b[128])^(a[22] & b[129])^(a[21] & b[130])^(a[20] & b[131])^(a[19] & b[132])^(a[18] & b[133])^(a[17] & b[134])^(a[16] & b[135])^(a[15] & b[136])^(a[14] & b[137])^(a[13] & b[138])^(a[12] & b[139])^(a[11] & b[140])^(a[10] & b[141])^(a[9] & b[142])^(a[8] & b[143])^(a[7] & b[144])^(a[6] & b[145])^(a[5] & b[146])^(a[4] & b[147])^(a[3] & b[148])^(a[2] & b[149])^(a[1] & b[150])^(a[0] & b[151]);
assign y[152] = (a[152] & b[0])^(a[151] & b[1])^(a[150] & b[2])^(a[149] & b[3])^(a[148] & b[4])^(a[147] & b[5])^(a[146] & b[6])^(a[145] & b[7])^(a[144] & b[8])^(a[143] & b[9])^(a[142] & b[10])^(a[141] & b[11])^(a[140] & b[12])^(a[139] & b[13])^(a[138] & b[14])^(a[137] & b[15])^(a[136] & b[16])^(a[135] & b[17])^(a[134] & b[18])^(a[133] & b[19])^(a[132] & b[20])^(a[131] & b[21])^(a[130] & b[22])^(a[129] & b[23])^(a[128] & b[24])^(a[127] & b[25])^(a[126] & b[26])^(a[125] & b[27])^(a[124] & b[28])^(a[123] & b[29])^(a[122] & b[30])^(a[121] & b[31])^(a[120] & b[32])^(a[119] & b[33])^(a[118] & b[34])^(a[117] & b[35])^(a[116] & b[36])^(a[115] & b[37])^(a[114] & b[38])^(a[113] & b[39])^(a[112] & b[40])^(a[111] & b[41])^(a[110] & b[42])^(a[109] & b[43])^(a[108] & b[44])^(a[107] & b[45])^(a[106] & b[46])^(a[105] & b[47])^(a[104] & b[48])^(a[103] & b[49])^(a[102] & b[50])^(a[101] & b[51])^(a[100] & b[52])^(a[99] & b[53])^(a[98] & b[54])^(a[97] & b[55])^(a[96] & b[56])^(a[95] & b[57])^(a[94] & b[58])^(a[93] & b[59])^(a[92] & b[60])^(a[91] & b[61])^(a[90] & b[62])^(a[89] & b[63])^(a[88] & b[64])^(a[87] & b[65])^(a[86] & b[66])^(a[85] & b[67])^(a[84] & b[68])^(a[83] & b[69])^(a[82] & b[70])^(a[81] & b[71])^(a[80] & b[72])^(a[79] & b[73])^(a[78] & b[74])^(a[77] & b[75])^(a[76] & b[76])^(a[75] & b[77])^(a[74] & b[78])^(a[73] & b[79])^(a[72] & b[80])^(a[71] & b[81])^(a[70] & b[82])^(a[69] & b[83])^(a[68] & b[84])^(a[67] & b[85])^(a[66] & b[86])^(a[65] & b[87])^(a[64] & b[88])^(a[63] & b[89])^(a[62] & b[90])^(a[61] & b[91])^(a[60] & b[92])^(a[59] & b[93])^(a[58] & b[94])^(a[57] & b[95])^(a[56] & b[96])^(a[55] & b[97])^(a[54] & b[98])^(a[53] & b[99])^(a[52] & b[100])^(a[51] & b[101])^(a[50] & b[102])^(a[49] & b[103])^(a[48] & b[104])^(a[47] & b[105])^(a[46] & b[106])^(a[45] & b[107])^(a[44] & b[108])^(a[43] & b[109])^(a[42] & b[110])^(a[41] & b[111])^(a[40] & b[112])^(a[39] & b[113])^(a[38] & b[114])^(a[37] & b[115])^(a[36] & b[116])^(a[35] & b[117])^(a[34] & b[118])^(a[33] & b[119])^(a[32] & b[120])^(a[31] & b[121])^(a[30] & b[122])^(a[29] & b[123])^(a[28] & b[124])^(a[27] & b[125])^(a[26] & b[126])^(a[25] & b[127])^(a[24] & b[128])^(a[23] & b[129])^(a[22] & b[130])^(a[21] & b[131])^(a[20] & b[132])^(a[19] & b[133])^(a[18] & b[134])^(a[17] & b[135])^(a[16] & b[136])^(a[15] & b[137])^(a[14] & b[138])^(a[13] & b[139])^(a[12] & b[140])^(a[11] & b[141])^(a[10] & b[142])^(a[9] & b[143])^(a[8] & b[144])^(a[7] & b[145])^(a[6] & b[146])^(a[5] & b[147])^(a[4] & b[148])^(a[3] & b[149])^(a[2] & b[150])^(a[1] & b[151])^(a[0] & b[152]);
assign y[153] = (a[153] & b[0])^(a[152] & b[1])^(a[151] & b[2])^(a[150] & b[3])^(a[149] & b[4])^(a[148] & b[5])^(a[147] & b[6])^(a[146] & b[7])^(a[145] & b[8])^(a[144] & b[9])^(a[143] & b[10])^(a[142] & b[11])^(a[141] & b[12])^(a[140] & b[13])^(a[139] & b[14])^(a[138] & b[15])^(a[137] & b[16])^(a[136] & b[17])^(a[135] & b[18])^(a[134] & b[19])^(a[133] & b[20])^(a[132] & b[21])^(a[131] & b[22])^(a[130] & b[23])^(a[129] & b[24])^(a[128] & b[25])^(a[127] & b[26])^(a[126] & b[27])^(a[125] & b[28])^(a[124] & b[29])^(a[123] & b[30])^(a[122] & b[31])^(a[121] & b[32])^(a[120] & b[33])^(a[119] & b[34])^(a[118] & b[35])^(a[117] & b[36])^(a[116] & b[37])^(a[115] & b[38])^(a[114] & b[39])^(a[113] & b[40])^(a[112] & b[41])^(a[111] & b[42])^(a[110] & b[43])^(a[109] & b[44])^(a[108] & b[45])^(a[107] & b[46])^(a[106] & b[47])^(a[105] & b[48])^(a[104] & b[49])^(a[103] & b[50])^(a[102] & b[51])^(a[101] & b[52])^(a[100] & b[53])^(a[99] & b[54])^(a[98] & b[55])^(a[97] & b[56])^(a[96] & b[57])^(a[95] & b[58])^(a[94] & b[59])^(a[93] & b[60])^(a[92] & b[61])^(a[91] & b[62])^(a[90] & b[63])^(a[89] & b[64])^(a[88] & b[65])^(a[87] & b[66])^(a[86] & b[67])^(a[85] & b[68])^(a[84] & b[69])^(a[83] & b[70])^(a[82] & b[71])^(a[81] & b[72])^(a[80] & b[73])^(a[79] & b[74])^(a[78] & b[75])^(a[77] & b[76])^(a[76] & b[77])^(a[75] & b[78])^(a[74] & b[79])^(a[73] & b[80])^(a[72] & b[81])^(a[71] & b[82])^(a[70] & b[83])^(a[69] & b[84])^(a[68] & b[85])^(a[67] & b[86])^(a[66] & b[87])^(a[65] & b[88])^(a[64] & b[89])^(a[63] & b[90])^(a[62] & b[91])^(a[61] & b[92])^(a[60] & b[93])^(a[59] & b[94])^(a[58] & b[95])^(a[57] & b[96])^(a[56] & b[97])^(a[55] & b[98])^(a[54] & b[99])^(a[53] & b[100])^(a[52] & b[101])^(a[51] & b[102])^(a[50] & b[103])^(a[49] & b[104])^(a[48] & b[105])^(a[47] & b[106])^(a[46] & b[107])^(a[45] & b[108])^(a[44] & b[109])^(a[43] & b[110])^(a[42] & b[111])^(a[41] & b[112])^(a[40] & b[113])^(a[39] & b[114])^(a[38] & b[115])^(a[37] & b[116])^(a[36] & b[117])^(a[35] & b[118])^(a[34] & b[119])^(a[33] & b[120])^(a[32] & b[121])^(a[31] & b[122])^(a[30] & b[123])^(a[29] & b[124])^(a[28] & b[125])^(a[27] & b[126])^(a[26] & b[127])^(a[25] & b[128])^(a[24] & b[129])^(a[23] & b[130])^(a[22] & b[131])^(a[21] & b[132])^(a[20] & b[133])^(a[19] & b[134])^(a[18] & b[135])^(a[17] & b[136])^(a[16] & b[137])^(a[15] & b[138])^(a[14] & b[139])^(a[13] & b[140])^(a[12] & b[141])^(a[11] & b[142])^(a[10] & b[143])^(a[9] & b[144])^(a[8] & b[145])^(a[7] & b[146])^(a[6] & b[147])^(a[5] & b[148])^(a[4] & b[149])^(a[3] & b[150])^(a[2] & b[151])^(a[1] & b[152])^(a[0] & b[153]);
assign y[154] = (a[154] & b[0])^(a[153] & b[1])^(a[152] & b[2])^(a[151] & b[3])^(a[150] & b[4])^(a[149] & b[5])^(a[148] & b[6])^(a[147] & b[7])^(a[146] & b[8])^(a[145] & b[9])^(a[144] & b[10])^(a[143] & b[11])^(a[142] & b[12])^(a[141] & b[13])^(a[140] & b[14])^(a[139] & b[15])^(a[138] & b[16])^(a[137] & b[17])^(a[136] & b[18])^(a[135] & b[19])^(a[134] & b[20])^(a[133] & b[21])^(a[132] & b[22])^(a[131] & b[23])^(a[130] & b[24])^(a[129] & b[25])^(a[128] & b[26])^(a[127] & b[27])^(a[126] & b[28])^(a[125] & b[29])^(a[124] & b[30])^(a[123] & b[31])^(a[122] & b[32])^(a[121] & b[33])^(a[120] & b[34])^(a[119] & b[35])^(a[118] & b[36])^(a[117] & b[37])^(a[116] & b[38])^(a[115] & b[39])^(a[114] & b[40])^(a[113] & b[41])^(a[112] & b[42])^(a[111] & b[43])^(a[110] & b[44])^(a[109] & b[45])^(a[108] & b[46])^(a[107] & b[47])^(a[106] & b[48])^(a[105] & b[49])^(a[104] & b[50])^(a[103] & b[51])^(a[102] & b[52])^(a[101] & b[53])^(a[100] & b[54])^(a[99] & b[55])^(a[98] & b[56])^(a[97] & b[57])^(a[96] & b[58])^(a[95] & b[59])^(a[94] & b[60])^(a[93] & b[61])^(a[92] & b[62])^(a[91] & b[63])^(a[90] & b[64])^(a[89] & b[65])^(a[88] & b[66])^(a[87] & b[67])^(a[86] & b[68])^(a[85] & b[69])^(a[84] & b[70])^(a[83] & b[71])^(a[82] & b[72])^(a[81] & b[73])^(a[80] & b[74])^(a[79] & b[75])^(a[78] & b[76])^(a[77] & b[77])^(a[76] & b[78])^(a[75] & b[79])^(a[74] & b[80])^(a[73] & b[81])^(a[72] & b[82])^(a[71] & b[83])^(a[70] & b[84])^(a[69] & b[85])^(a[68] & b[86])^(a[67] & b[87])^(a[66] & b[88])^(a[65] & b[89])^(a[64] & b[90])^(a[63] & b[91])^(a[62] & b[92])^(a[61] & b[93])^(a[60] & b[94])^(a[59] & b[95])^(a[58] & b[96])^(a[57] & b[97])^(a[56] & b[98])^(a[55] & b[99])^(a[54] & b[100])^(a[53] & b[101])^(a[52] & b[102])^(a[51] & b[103])^(a[50] & b[104])^(a[49] & b[105])^(a[48] & b[106])^(a[47] & b[107])^(a[46] & b[108])^(a[45] & b[109])^(a[44] & b[110])^(a[43] & b[111])^(a[42] & b[112])^(a[41] & b[113])^(a[40] & b[114])^(a[39] & b[115])^(a[38] & b[116])^(a[37] & b[117])^(a[36] & b[118])^(a[35] & b[119])^(a[34] & b[120])^(a[33] & b[121])^(a[32] & b[122])^(a[31] & b[123])^(a[30] & b[124])^(a[29] & b[125])^(a[28] & b[126])^(a[27] & b[127])^(a[26] & b[128])^(a[25] & b[129])^(a[24] & b[130])^(a[23] & b[131])^(a[22] & b[132])^(a[21] & b[133])^(a[20] & b[134])^(a[19] & b[135])^(a[18] & b[136])^(a[17] & b[137])^(a[16] & b[138])^(a[15] & b[139])^(a[14] & b[140])^(a[13] & b[141])^(a[12] & b[142])^(a[11] & b[143])^(a[10] & b[144])^(a[9] & b[145])^(a[8] & b[146])^(a[7] & b[147])^(a[6] & b[148])^(a[5] & b[149])^(a[4] & b[150])^(a[3] & b[151])^(a[2] & b[152])^(a[1] & b[153])^(a[0] & b[154]);
assign y[155] = (a[155] & b[0])^(a[154] & b[1])^(a[153] & b[2])^(a[152] & b[3])^(a[151] & b[4])^(a[150] & b[5])^(a[149] & b[6])^(a[148] & b[7])^(a[147] & b[8])^(a[146] & b[9])^(a[145] & b[10])^(a[144] & b[11])^(a[143] & b[12])^(a[142] & b[13])^(a[141] & b[14])^(a[140] & b[15])^(a[139] & b[16])^(a[138] & b[17])^(a[137] & b[18])^(a[136] & b[19])^(a[135] & b[20])^(a[134] & b[21])^(a[133] & b[22])^(a[132] & b[23])^(a[131] & b[24])^(a[130] & b[25])^(a[129] & b[26])^(a[128] & b[27])^(a[127] & b[28])^(a[126] & b[29])^(a[125] & b[30])^(a[124] & b[31])^(a[123] & b[32])^(a[122] & b[33])^(a[121] & b[34])^(a[120] & b[35])^(a[119] & b[36])^(a[118] & b[37])^(a[117] & b[38])^(a[116] & b[39])^(a[115] & b[40])^(a[114] & b[41])^(a[113] & b[42])^(a[112] & b[43])^(a[111] & b[44])^(a[110] & b[45])^(a[109] & b[46])^(a[108] & b[47])^(a[107] & b[48])^(a[106] & b[49])^(a[105] & b[50])^(a[104] & b[51])^(a[103] & b[52])^(a[102] & b[53])^(a[101] & b[54])^(a[100] & b[55])^(a[99] & b[56])^(a[98] & b[57])^(a[97] & b[58])^(a[96] & b[59])^(a[95] & b[60])^(a[94] & b[61])^(a[93] & b[62])^(a[92] & b[63])^(a[91] & b[64])^(a[90] & b[65])^(a[89] & b[66])^(a[88] & b[67])^(a[87] & b[68])^(a[86] & b[69])^(a[85] & b[70])^(a[84] & b[71])^(a[83] & b[72])^(a[82] & b[73])^(a[81] & b[74])^(a[80] & b[75])^(a[79] & b[76])^(a[78] & b[77])^(a[77] & b[78])^(a[76] & b[79])^(a[75] & b[80])^(a[74] & b[81])^(a[73] & b[82])^(a[72] & b[83])^(a[71] & b[84])^(a[70] & b[85])^(a[69] & b[86])^(a[68] & b[87])^(a[67] & b[88])^(a[66] & b[89])^(a[65] & b[90])^(a[64] & b[91])^(a[63] & b[92])^(a[62] & b[93])^(a[61] & b[94])^(a[60] & b[95])^(a[59] & b[96])^(a[58] & b[97])^(a[57] & b[98])^(a[56] & b[99])^(a[55] & b[100])^(a[54] & b[101])^(a[53] & b[102])^(a[52] & b[103])^(a[51] & b[104])^(a[50] & b[105])^(a[49] & b[106])^(a[48] & b[107])^(a[47] & b[108])^(a[46] & b[109])^(a[45] & b[110])^(a[44] & b[111])^(a[43] & b[112])^(a[42] & b[113])^(a[41] & b[114])^(a[40] & b[115])^(a[39] & b[116])^(a[38] & b[117])^(a[37] & b[118])^(a[36] & b[119])^(a[35] & b[120])^(a[34] & b[121])^(a[33] & b[122])^(a[32] & b[123])^(a[31] & b[124])^(a[30] & b[125])^(a[29] & b[126])^(a[28] & b[127])^(a[27] & b[128])^(a[26] & b[129])^(a[25] & b[130])^(a[24] & b[131])^(a[23] & b[132])^(a[22] & b[133])^(a[21] & b[134])^(a[20] & b[135])^(a[19] & b[136])^(a[18] & b[137])^(a[17] & b[138])^(a[16] & b[139])^(a[15] & b[140])^(a[14] & b[141])^(a[13] & b[142])^(a[12] & b[143])^(a[11] & b[144])^(a[10] & b[145])^(a[9] & b[146])^(a[8] & b[147])^(a[7] & b[148])^(a[6] & b[149])^(a[5] & b[150])^(a[4] & b[151])^(a[3] & b[152])^(a[2] & b[153])^(a[1] & b[154])^(a[0] & b[155]);
assign y[156] = (a[156] & b[0])^(a[155] & b[1])^(a[154] & b[2])^(a[153] & b[3])^(a[152] & b[4])^(a[151] & b[5])^(a[150] & b[6])^(a[149] & b[7])^(a[148] & b[8])^(a[147] & b[9])^(a[146] & b[10])^(a[145] & b[11])^(a[144] & b[12])^(a[143] & b[13])^(a[142] & b[14])^(a[141] & b[15])^(a[140] & b[16])^(a[139] & b[17])^(a[138] & b[18])^(a[137] & b[19])^(a[136] & b[20])^(a[135] & b[21])^(a[134] & b[22])^(a[133] & b[23])^(a[132] & b[24])^(a[131] & b[25])^(a[130] & b[26])^(a[129] & b[27])^(a[128] & b[28])^(a[127] & b[29])^(a[126] & b[30])^(a[125] & b[31])^(a[124] & b[32])^(a[123] & b[33])^(a[122] & b[34])^(a[121] & b[35])^(a[120] & b[36])^(a[119] & b[37])^(a[118] & b[38])^(a[117] & b[39])^(a[116] & b[40])^(a[115] & b[41])^(a[114] & b[42])^(a[113] & b[43])^(a[112] & b[44])^(a[111] & b[45])^(a[110] & b[46])^(a[109] & b[47])^(a[108] & b[48])^(a[107] & b[49])^(a[106] & b[50])^(a[105] & b[51])^(a[104] & b[52])^(a[103] & b[53])^(a[102] & b[54])^(a[101] & b[55])^(a[100] & b[56])^(a[99] & b[57])^(a[98] & b[58])^(a[97] & b[59])^(a[96] & b[60])^(a[95] & b[61])^(a[94] & b[62])^(a[93] & b[63])^(a[92] & b[64])^(a[91] & b[65])^(a[90] & b[66])^(a[89] & b[67])^(a[88] & b[68])^(a[87] & b[69])^(a[86] & b[70])^(a[85] & b[71])^(a[84] & b[72])^(a[83] & b[73])^(a[82] & b[74])^(a[81] & b[75])^(a[80] & b[76])^(a[79] & b[77])^(a[78] & b[78])^(a[77] & b[79])^(a[76] & b[80])^(a[75] & b[81])^(a[74] & b[82])^(a[73] & b[83])^(a[72] & b[84])^(a[71] & b[85])^(a[70] & b[86])^(a[69] & b[87])^(a[68] & b[88])^(a[67] & b[89])^(a[66] & b[90])^(a[65] & b[91])^(a[64] & b[92])^(a[63] & b[93])^(a[62] & b[94])^(a[61] & b[95])^(a[60] & b[96])^(a[59] & b[97])^(a[58] & b[98])^(a[57] & b[99])^(a[56] & b[100])^(a[55] & b[101])^(a[54] & b[102])^(a[53] & b[103])^(a[52] & b[104])^(a[51] & b[105])^(a[50] & b[106])^(a[49] & b[107])^(a[48] & b[108])^(a[47] & b[109])^(a[46] & b[110])^(a[45] & b[111])^(a[44] & b[112])^(a[43] & b[113])^(a[42] & b[114])^(a[41] & b[115])^(a[40] & b[116])^(a[39] & b[117])^(a[38] & b[118])^(a[37] & b[119])^(a[36] & b[120])^(a[35] & b[121])^(a[34] & b[122])^(a[33] & b[123])^(a[32] & b[124])^(a[31] & b[125])^(a[30] & b[126])^(a[29] & b[127])^(a[28] & b[128])^(a[27] & b[129])^(a[26] & b[130])^(a[25] & b[131])^(a[24] & b[132])^(a[23] & b[133])^(a[22] & b[134])^(a[21] & b[135])^(a[20] & b[136])^(a[19] & b[137])^(a[18] & b[138])^(a[17] & b[139])^(a[16] & b[140])^(a[15] & b[141])^(a[14] & b[142])^(a[13] & b[143])^(a[12] & b[144])^(a[11] & b[145])^(a[10] & b[146])^(a[9] & b[147])^(a[8] & b[148])^(a[7] & b[149])^(a[6] & b[150])^(a[5] & b[151])^(a[4] & b[152])^(a[3] & b[153])^(a[2] & b[154])^(a[1] & b[155])^(a[0] & b[156]);
assign y[157] = (a[157] & b[0])^(a[156] & b[1])^(a[155] & b[2])^(a[154] & b[3])^(a[153] & b[4])^(a[152] & b[5])^(a[151] & b[6])^(a[150] & b[7])^(a[149] & b[8])^(a[148] & b[9])^(a[147] & b[10])^(a[146] & b[11])^(a[145] & b[12])^(a[144] & b[13])^(a[143] & b[14])^(a[142] & b[15])^(a[141] & b[16])^(a[140] & b[17])^(a[139] & b[18])^(a[138] & b[19])^(a[137] & b[20])^(a[136] & b[21])^(a[135] & b[22])^(a[134] & b[23])^(a[133] & b[24])^(a[132] & b[25])^(a[131] & b[26])^(a[130] & b[27])^(a[129] & b[28])^(a[128] & b[29])^(a[127] & b[30])^(a[126] & b[31])^(a[125] & b[32])^(a[124] & b[33])^(a[123] & b[34])^(a[122] & b[35])^(a[121] & b[36])^(a[120] & b[37])^(a[119] & b[38])^(a[118] & b[39])^(a[117] & b[40])^(a[116] & b[41])^(a[115] & b[42])^(a[114] & b[43])^(a[113] & b[44])^(a[112] & b[45])^(a[111] & b[46])^(a[110] & b[47])^(a[109] & b[48])^(a[108] & b[49])^(a[107] & b[50])^(a[106] & b[51])^(a[105] & b[52])^(a[104] & b[53])^(a[103] & b[54])^(a[102] & b[55])^(a[101] & b[56])^(a[100] & b[57])^(a[99] & b[58])^(a[98] & b[59])^(a[97] & b[60])^(a[96] & b[61])^(a[95] & b[62])^(a[94] & b[63])^(a[93] & b[64])^(a[92] & b[65])^(a[91] & b[66])^(a[90] & b[67])^(a[89] & b[68])^(a[88] & b[69])^(a[87] & b[70])^(a[86] & b[71])^(a[85] & b[72])^(a[84] & b[73])^(a[83] & b[74])^(a[82] & b[75])^(a[81] & b[76])^(a[80] & b[77])^(a[79] & b[78])^(a[78] & b[79])^(a[77] & b[80])^(a[76] & b[81])^(a[75] & b[82])^(a[74] & b[83])^(a[73] & b[84])^(a[72] & b[85])^(a[71] & b[86])^(a[70] & b[87])^(a[69] & b[88])^(a[68] & b[89])^(a[67] & b[90])^(a[66] & b[91])^(a[65] & b[92])^(a[64] & b[93])^(a[63] & b[94])^(a[62] & b[95])^(a[61] & b[96])^(a[60] & b[97])^(a[59] & b[98])^(a[58] & b[99])^(a[57] & b[100])^(a[56] & b[101])^(a[55] & b[102])^(a[54] & b[103])^(a[53] & b[104])^(a[52] & b[105])^(a[51] & b[106])^(a[50] & b[107])^(a[49] & b[108])^(a[48] & b[109])^(a[47] & b[110])^(a[46] & b[111])^(a[45] & b[112])^(a[44] & b[113])^(a[43] & b[114])^(a[42] & b[115])^(a[41] & b[116])^(a[40] & b[117])^(a[39] & b[118])^(a[38] & b[119])^(a[37] & b[120])^(a[36] & b[121])^(a[35] & b[122])^(a[34] & b[123])^(a[33] & b[124])^(a[32] & b[125])^(a[31] & b[126])^(a[30] & b[127])^(a[29] & b[128])^(a[28] & b[129])^(a[27] & b[130])^(a[26] & b[131])^(a[25] & b[132])^(a[24] & b[133])^(a[23] & b[134])^(a[22] & b[135])^(a[21] & b[136])^(a[20] & b[137])^(a[19] & b[138])^(a[18] & b[139])^(a[17] & b[140])^(a[16] & b[141])^(a[15] & b[142])^(a[14] & b[143])^(a[13] & b[144])^(a[12] & b[145])^(a[11] & b[146])^(a[10] & b[147])^(a[9] & b[148])^(a[8] & b[149])^(a[7] & b[150])^(a[6] & b[151])^(a[5] & b[152])^(a[4] & b[153])^(a[3] & b[154])^(a[2] & b[155])^(a[1] & b[156])^(a[0] & b[157]);
assign y[158] = (a[158] & b[0])^(a[157] & b[1])^(a[156] & b[2])^(a[155] & b[3])^(a[154] & b[4])^(a[153] & b[5])^(a[152] & b[6])^(a[151] & b[7])^(a[150] & b[8])^(a[149] & b[9])^(a[148] & b[10])^(a[147] & b[11])^(a[146] & b[12])^(a[145] & b[13])^(a[144] & b[14])^(a[143] & b[15])^(a[142] & b[16])^(a[141] & b[17])^(a[140] & b[18])^(a[139] & b[19])^(a[138] & b[20])^(a[137] & b[21])^(a[136] & b[22])^(a[135] & b[23])^(a[134] & b[24])^(a[133] & b[25])^(a[132] & b[26])^(a[131] & b[27])^(a[130] & b[28])^(a[129] & b[29])^(a[128] & b[30])^(a[127] & b[31])^(a[126] & b[32])^(a[125] & b[33])^(a[124] & b[34])^(a[123] & b[35])^(a[122] & b[36])^(a[121] & b[37])^(a[120] & b[38])^(a[119] & b[39])^(a[118] & b[40])^(a[117] & b[41])^(a[116] & b[42])^(a[115] & b[43])^(a[114] & b[44])^(a[113] & b[45])^(a[112] & b[46])^(a[111] & b[47])^(a[110] & b[48])^(a[109] & b[49])^(a[108] & b[50])^(a[107] & b[51])^(a[106] & b[52])^(a[105] & b[53])^(a[104] & b[54])^(a[103] & b[55])^(a[102] & b[56])^(a[101] & b[57])^(a[100] & b[58])^(a[99] & b[59])^(a[98] & b[60])^(a[97] & b[61])^(a[96] & b[62])^(a[95] & b[63])^(a[94] & b[64])^(a[93] & b[65])^(a[92] & b[66])^(a[91] & b[67])^(a[90] & b[68])^(a[89] & b[69])^(a[88] & b[70])^(a[87] & b[71])^(a[86] & b[72])^(a[85] & b[73])^(a[84] & b[74])^(a[83] & b[75])^(a[82] & b[76])^(a[81] & b[77])^(a[80] & b[78])^(a[79] & b[79])^(a[78] & b[80])^(a[77] & b[81])^(a[76] & b[82])^(a[75] & b[83])^(a[74] & b[84])^(a[73] & b[85])^(a[72] & b[86])^(a[71] & b[87])^(a[70] & b[88])^(a[69] & b[89])^(a[68] & b[90])^(a[67] & b[91])^(a[66] & b[92])^(a[65] & b[93])^(a[64] & b[94])^(a[63] & b[95])^(a[62] & b[96])^(a[61] & b[97])^(a[60] & b[98])^(a[59] & b[99])^(a[58] & b[100])^(a[57] & b[101])^(a[56] & b[102])^(a[55] & b[103])^(a[54] & b[104])^(a[53] & b[105])^(a[52] & b[106])^(a[51] & b[107])^(a[50] & b[108])^(a[49] & b[109])^(a[48] & b[110])^(a[47] & b[111])^(a[46] & b[112])^(a[45] & b[113])^(a[44] & b[114])^(a[43] & b[115])^(a[42] & b[116])^(a[41] & b[117])^(a[40] & b[118])^(a[39] & b[119])^(a[38] & b[120])^(a[37] & b[121])^(a[36] & b[122])^(a[35] & b[123])^(a[34] & b[124])^(a[33] & b[125])^(a[32] & b[126])^(a[31] & b[127])^(a[30] & b[128])^(a[29] & b[129])^(a[28] & b[130])^(a[27] & b[131])^(a[26] & b[132])^(a[25] & b[133])^(a[24] & b[134])^(a[23] & b[135])^(a[22] & b[136])^(a[21] & b[137])^(a[20] & b[138])^(a[19] & b[139])^(a[18] & b[140])^(a[17] & b[141])^(a[16] & b[142])^(a[15] & b[143])^(a[14] & b[144])^(a[13] & b[145])^(a[12] & b[146])^(a[11] & b[147])^(a[10] & b[148])^(a[9] & b[149])^(a[8] & b[150])^(a[7] & b[151])^(a[6] & b[152])^(a[5] & b[153])^(a[4] & b[154])^(a[3] & b[155])^(a[2] & b[156])^(a[1] & b[157])^(a[0] & b[158]);
assign y[159] = (a[159] & b[0])^(a[158] & b[1])^(a[157] & b[2])^(a[156] & b[3])^(a[155] & b[4])^(a[154] & b[5])^(a[153] & b[6])^(a[152] & b[7])^(a[151] & b[8])^(a[150] & b[9])^(a[149] & b[10])^(a[148] & b[11])^(a[147] & b[12])^(a[146] & b[13])^(a[145] & b[14])^(a[144] & b[15])^(a[143] & b[16])^(a[142] & b[17])^(a[141] & b[18])^(a[140] & b[19])^(a[139] & b[20])^(a[138] & b[21])^(a[137] & b[22])^(a[136] & b[23])^(a[135] & b[24])^(a[134] & b[25])^(a[133] & b[26])^(a[132] & b[27])^(a[131] & b[28])^(a[130] & b[29])^(a[129] & b[30])^(a[128] & b[31])^(a[127] & b[32])^(a[126] & b[33])^(a[125] & b[34])^(a[124] & b[35])^(a[123] & b[36])^(a[122] & b[37])^(a[121] & b[38])^(a[120] & b[39])^(a[119] & b[40])^(a[118] & b[41])^(a[117] & b[42])^(a[116] & b[43])^(a[115] & b[44])^(a[114] & b[45])^(a[113] & b[46])^(a[112] & b[47])^(a[111] & b[48])^(a[110] & b[49])^(a[109] & b[50])^(a[108] & b[51])^(a[107] & b[52])^(a[106] & b[53])^(a[105] & b[54])^(a[104] & b[55])^(a[103] & b[56])^(a[102] & b[57])^(a[101] & b[58])^(a[100] & b[59])^(a[99] & b[60])^(a[98] & b[61])^(a[97] & b[62])^(a[96] & b[63])^(a[95] & b[64])^(a[94] & b[65])^(a[93] & b[66])^(a[92] & b[67])^(a[91] & b[68])^(a[90] & b[69])^(a[89] & b[70])^(a[88] & b[71])^(a[87] & b[72])^(a[86] & b[73])^(a[85] & b[74])^(a[84] & b[75])^(a[83] & b[76])^(a[82] & b[77])^(a[81] & b[78])^(a[80] & b[79])^(a[79] & b[80])^(a[78] & b[81])^(a[77] & b[82])^(a[76] & b[83])^(a[75] & b[84])^(a[74] & b[85])^(a[73] & b[86])^(a[72] & b[87])^(a[71] & b[88])^(a[70] & b[89])^(a[69] & b[90])^(a[68] & b[91])^(a[67] & b[92])^(a[66] & b[93])^(a[65] & b[94])^(a[64] & b[95])^(a[63] & b[96])^(a[62] & b[97])^(a[61] & b[98])^(a[60] & b[99])^(a[59] & b[100])^(a[58] & b[101])^(a[57] & b[102])^(a[56] & b[103])^(a[55] & b[104])^(a[54] & b[105])^(a[53] & b[106])^(a[52] & b[107])^(a[51] & b[108])^(a[50] & b[109])^(a[49] & b[110])^(a[48] & b[111])^(a[47] & b[112])^(a[46] & b[113])^(a[45] & b[114])^(a[44] & b[115])^(a[43] & b[116])^(a[42] & b[117])^(a[41] & b[118])^(a[40] & b[119])^(a[39] & b[120])^(a[38] & b[121])^(a[37] & b[122])^(a[36] & b[123])^(a[35] & b[124])^(a[34] & b[125])^(a[33] & b[126])^(a[32] & b[127])^(a[31] & b[128])^(a[30] & b[129])^(a[29] & b[130])^(a[28] & b[131])^(a[27] & b[132])^(a[26] & b[133])^(a[25] & b[134])^(a[24] & b[135])^(a[23] & b[136])^(a[22] & b[137])^(a[21] & b[138])^(a[20] & b[139])^(a[19] & b[140])^(a[18] & b[141])^(a[17] & b[142])^(a[16] & b[143])^(a[15] & b[144])^(a[14] & b[145])^(a[13] & b[146])^(a[12] & b[147])^(a[11] & b[148])^(a[10] & b[149])^(a[9] & b[150])^(a[8] & b[151])^(a[7] & b[152])^(a[6] & b[153])^(a[5] & b[154])^(a[4] & b[155])^(a[3] & b[156])^(a[2] & b[157])^(a[1] & b[158])^(a[0] & b[159]);
assign y[160] = (a[160] & b[0])^(a[159] & b[1])^(a[158] & b[2])^(a[157] & b[3])^(a[156] & b[4])^(a[155] & b[5])^(a[154] & b[6])^(a[153] & b[7])^(a[152] & b[8])^(a[151] & b[9])^(a[150] & b[10])^(a[149] & b[11])^(a[148] & b[12])^(a[147] & b[13])^(a[146] & b[14])^(a[145] & b[15])^(a[144] & b[16])^(a[143] & b[17])^(a[142] & b[18])^(a[141] & b[19])^(a[140] & b[20])^(a[139] & b[21])^(a[138] & b[22])^(a[137] & b[23])^(a[136] & b[24])^(a[135] & b[25])^(a[134] & b[26])^(a[133] & b[27])^(a[132] & b[28])^(a[131] & b[29])^(a[130] & b[30])^(a[129] & b[31])^(a[128] & b[32])^(a[127] & b[33])^(a[126] & b[34])^(a[125] & b[35])^(a[124] & b[36])^(a[123] & b[37])^(a[122] & b[38])^(a[121] & b[39])^(a[120] & b[40])^(a[119] & b[41])^(a[118] & b[42])^(a[117] & b[43])^(a[116] & b[44])^(a[115] & b[45])^(a[114] & b[46])^(a[113] & b[47])^(a[112] & b[48])^(a[111] & b[49])^(a[110] & b[50])^(a[109] & b[51])^(a[108] & b[52])^(a[107] & b[53])^(a[106] & b[54])^(a[105] & b[55])^(a[104] & b[56])^(a[103] & b[57])^(a[102] & b[58])^(a[101] & b[59])^(a[100] & b[60])^(a[99] & b[61])^(a[98] & b[62])^(a[97] & b[63])^(a[96] & b[64])^(a[95] & b[65])^(a[94] & b[66])^(a[93] & b[67])^(a[92] & b[68])^(a[91] & b[69])^(a[90] & b[70])^(a[89] & b[71])^(a[88] & b[72])^(a[87] & b[73])^(a[86] & b[74])^(a[85] & b[75])^(a[84] & b[76])^(a[83] & b[77])^(a[82] & b[78])^(a[81] & b[79])^(a[80] & b[80])^(a[79] & b[81])^(a[78] & b[82])^(a[77] & b[83])^(a[76] & b[84])^(a[75] & b[85])^(a[74] & b[86])^(a[73] & b[87])^(a[72] & b[88])^(a[71] & b[89])^(a[70] & b[90])^(a[69] & b[91])^(a[68] & b[92])^(a[67] & b[93])^(a[66] & b[94])^(a[65] & b[95])^(a[64] & b[96])^(a[63] & b[97])^(a[62] & b[98])^(a[61] & b[99])^(a[60] & b[100])^(a[59] & b[101])^(a[58] & b[102])^(a[57] & b[103])^(a[56] & b[104])^(a[55] & b[105])^(a[54] & b[106])^(a[53] & b[107])^(a[52] & b[108])^(a[51] & b[109])^(a[50] & b[110])^(a[49] & b[111])^(a[48] & b[112])^(a[47] & b[113])^(a[46] & b[114])^(a[45] & b[115])^(a[44] & b[116])^(a[43] & b[117])^(a[42] & b[118])^(a[41] & b[119])^(a[40] & b[120])^(a[39] & b[121])^(a[38] & b[122])^(a[37] & b[123])^(a[36] & b[124])^(a[35] & b[125])^(a[34] & b[126])^(a[33] & b[127])^(a[32] & b[128])^(a[31] & b[129])^(a[30] & b[130])^(a[29] & b[131])^(a[28] & b[132])^(a[27] & b[133])^(a[26] & b[134])^(a[25] & b[135])^(a[24] & b[136])^(a[23] & b[137])^(a[22] & b[138])^(a[21] & b[139])^(a[20] & b[140])^(a[19] & b[141])^(a[18] & b[142])^(a[17] & b[143])^(a[16] & b[144])^(a[15] & b[145])^(a[14] & b[146])^(a[13] & b[147])^(a[12] & b[148])^(a[11] & b[149])^(a[10] & b[150])^(a[9] & b[151])^(a[8] & b[152])^(a[7] & b[153])^(a[6] & b[154])^(a[5] & b[155])^(a[4] & b[156])^(a[3] & b[157])^(a[2] & b[158])^(a[1] & b[159])^(a[0] & b[160]);
assign y[161] = (a[161] & b[0])^(a[160] & b[1])^(a[159] & b[2])^(a[158] & b[3])^(a[157] & b[4])^(a[156] & b[5])^(a[155] & b[6])^(a[154] & b[7])^(a[153] & b[8])^(a[152] & b[9])^(a[151] & b[10])^(a[150] & b[11])^(a[149] & b[12])^(a[148] & b[13])^(a[147] & b[14])^(a[146] & b[15])^(a[145] & b[16])^(a[144] & b[17])^(a[143] & b[18])^(a[142] & b[19])^(a[141] & b[20])^(a[140] & b[21])^(a[139] & b[22])^(a[138] & b[23])^(a[137] & b[24])^(a[136] & b[25])^(a[135] & b[26])^(a[134] & b[27])^(a[133] & b[28])^(a[132] & b[29])^(a[131] & b[30])^(a[130] & b[31])^(a[129] & b[32])^(a[128] & b[33])^(a[127] & b[34])^(a[126] & b[35])^(a[125] & b[36])^(a[124] & b[37])^(a[123] & b[38])^(a[122] & b[39])^(a[121] & b[40])^(a[120] & b[41])^(a[119] & b[42])^(a[118] & b[43])^(a[117] & b[44])^(a[116] & b[45])^(a[115] & b[46])^(a[114] & b[47])^(a[113] & b[48])^(a[112] & b[49])^(a[111] & b[50])^(a[110] & b[51])^(a[109] & b[52])^(a[108] & b[53])^(a[107] & b[54])^(a[106] & b[55])^(a[105] & b[56])^(a[104] & b[57])^(a[103] & b[58])^(a[102] & b[59])^(a[101] & b[60])^(a[100] & b[61])^(a[99] & b[62])^(a[98] & b[63])^(a[97] & b[64])^(a[96] & b[65])^(a[95] & b[66])^(a[94] & b[67])^(a[93] & b[68])^(a[92] & b[69])^(a[91] & b[70])^(a[90] & b[71])^(a[89] & b[72])^(a[88] & b[73])^(a[87] & b[74])^(a[86] & b[75])^(a[85] & b[76])^(a[84] & b[77])^(a[83] & b[78])^(a[82] & b[79])^(a[81] & b[80])^(a[80] & b[81])^(a[79] & b[82])^(a[78] & b[83])^(a[77] & b[84])^(a[76] & b[85])^(a[75] & b[86])^(a[74] & b[87])^(a[73] & b[88])^(a[72] & b[89])^(a[71] & b[90])^(a[70] & b[91])^(a[69] & b[92])^(a[68] & b[93])^(a[67] & b[94])^(a[66] & b[95])^(a[65] & b[96])^(a[64] & b[97])^(a[63] & b[98])^(a[62] & b[99])^(a[61] & b[100])^(a[60] & b[101])^(a[59] & b[102])^(a[58] & b[103])^(a[57] & b[104])^(a[56] & b[105])^(a[55] & b[106])^(a[54] & b[107])^(a[53] & b[108])^(a[52] & b[109])^(a[51] & b[110])^(a[50] & b[111])^(a[49] & b[112])^(a[48] & b[113])^(a[47] & b[114])^(a[46] & b[115])^(a[45] & b[116])^(a[44] & b[117])^(a[43] & b[118])^(a[42] & b[119])^(a[41] & b[120])^(a[40] & b[121])^(a[39] & b[122])^(a[38] & b[123])^(a[37] & b[124])^(a[36] & b[125])^(a[35] & b[126])^(a[34] & b[127])^(a[33] & b[128])^(a[32] & b[129])^(a[31] & b[130])^(a[30] & b[131])^(a[29] & b[132])^(a[28] & b[133])^(a[27] & b[134])^(a[26] & b[135])^(a[25] & b[136])^(a[24] & b[137])^(a[23] & b[138])^(a[22] & b[139])^(a[21] & b[140])^(a[20] & b[141])^(a[19] & b[142])^(a[18] & b[143])^(a[17] & b[144])^(a[16] & b[145])^(a[15] & b[146])^(a[14] & b[147])^(a[13] & b[148])^(a[12] & b[149])^(a[11] & b[150])^(a[10] & b[151])^(a[9] & b[152])^(a[8] & b[153])^(a[7] & b[154])^(a[6] & b[155])^(a[5] & b[156])^(a[4] & b[157])^(a[3] & b[158])^(a[2] & b[159])^(a[1] & b[160])^(a[0] & b[161]);
assign y[162] = (a[162] & b[0])^(a[161] & b[1])^(a[160] & b[2])^(a[159] & b[3])^(a[158] & b[4])^(a[157] & b[5])^(a[156] & b[6])^(a[155] & b[7])^(a[154] & b[8])^(a[153] & b[9])^(a[152] & b[10])^(a[151] & b[11])^(a[150] & b[12])^(a[149] & b[13])^(a[148] & b[14])^(a[147] & b[15])^(a[146] & b[16])^(a[145] & b[17])^(a[144] & b[18])^(a[143] & b[19])^(a[142] & b[20])^(a[141] & b[21])^(a[140] & b[22])^(a[139] & b[23])^(a[138] & b[24])^(a[137] & b[25])^(a[136] & b[26])^(a[135] & b[27])^(a[134] & b[28])^(a[133] & b[29])^(a[132] & b[30])^(a[131] & b[31])^(a[130] & b[32])^(a[129] & b[33])^(a[128] & b[34])^(a[127] & b[35])^(a[126] & b[36])^(a[125] & b[37])^(a[124] & b[38])^(a[123] & b[39])^(a[122] & b[40])^(a[121] & b[41])^(a[120] & b[42])^(a[119] & b[43])^(a[118] & b[44])^(a[117] & b[45])^(a[116] & b[46])^(a[115] & b[47])^(a[114] & b[48])^(a[113] & b[49])^(a[112] & b[50])^(a[111] & b[51])^(a[110] & b[52])^(a[109] & b[53])^(a[108] & b[54])^(a[107] & b[55])^(a[106] & b[56])^(a[105] & b[57])^(a[104] & b[58])^(a[103] & b[59])^(a[102] & b[60])^(a[101] & b[61])^(a[100] & b[62])^(a[99] & b[63])^(a[98] & b[64])^(a[97] & b[65])^(a[96] & b[66])^(a[95] & b[67])^(a[94] & b[68])^(a[93] & b[69])^(a[92] & b[70])^(a[91] & b[71])^(a[90] & b[72])^(a[89] & b[73])^(a[88] & b[74])^(a[87] & b[75])^(a[86] & b[76])^(a[85] & b[77])^(a[84] & b[78])^(a[83] & b[79])^(a[82] & b[80])^(a[81] & b[81])^(a[80] & b[82])^(a[79] & b[83])^(a[78] & b[84])^(a[77] & b[85])^(a[76] & b[86])^(a[75] & b[87])^(a[74] & b[88])^(a[73] & b[89])^(a[72] & b[90])^(a[71] & b[91])^(a[70] & b[92])^(a[69] & b[93])^(a[68] & b[94])^(a[67] & b[95])^(a[66] & b[96])^(a[65] & b[97])^(a[64] & b[98])^(a[63] & b[99])^(a[62] & b[100])^(a[61] & b[101])^(a[60] & b[102])^(a[59] & b[103])^(a[58] & b[104])^(a[57] & b[105])^(a[56] & b[106])^(a[55] & b[107])^(a[54] & b[108])^(a[53] & b[109])^(a[52] & b[110])^(a[51] & b[111])^(a[50] & b[112])^(a[49] & b[113])^(a[48] & b[114])^(a[47] & b[115])^(a[46] & b[116])^(a[45] & b[117])^(a[44] & b[118])^(a[43] & b[119])^(a[42] & b[120])^(a[41] & b[121])^(a[40] & b[122])^(a[39] & b[123])^(a[38] & b[124])^(a[37] & b[125])^(a[36] & b[126])^(a[35] & b[127])^(a[34] & b[128])^(a[33] & b[129])^(a[32] & b[130])^(a[31] & b[131])^(a[30] & b[132])^(a[29] & b[133])^(a[28] & b[134])^(a[27] & b[135])^(a[26] & b[136])^(a[25] & b[137])^(a[24] & b[138])^(a[23] & b[139])^(a[22] & b[140])^(a[21] & b[141])^(a[20] & b[142])^(a[19] & b[143])^(a[18] & b[144])^(a[17] & b[145])^(a[16] & b[146])^(a[15] & b[147])^(a[14] & b[148])^(a[13] & b[149])^(a[12] & b[150])^(a[11] & b[151])^(a[10] & b[152])^(a[9] & b[153])^(a[8] & b[154])^(a[7] & b[155])^(a[6] & b[156])^(a[5] & b[157])^(a[4] & b[158])^(a[3] & b[159])^(a[2] & b[160])^(a[1] & b[161])^(a[0] & b[162]);
assign y[163] = (a[163] & b[0])^(a[162] & b[1])^(a[161] & b[2])^(a[160] & b[3])^(a[159] & b[4])^(a[158] & b[5])^(a[157] & b[6])^(a[156] & b[7])^(a[155] & b[8])^(a[154] & b[9])^(a[153] & b[10])^(a[152] & b[11])^(a[151] & b[12])^(a[150] & b[13])^(a[149] & b[14])^(a[148] & b[15])^(a[147] & b[16])^(a[146] & b[17])^(a[145] & b[18])^(a[144] & b[19])^(a[143] & b[20])^(a[142] & b[21])^(a[141] & b[22])^(a[140] & b[23])^(a[139] & b[24])^(a[138] & b[25])^(a[137] & b[26])^(a[136] & b[27])^(a[135] & b[28])^(a[134] & b[29])^(a[133] & b[30])^(a[132] & b[31])^(a[131] & b[32])^(a[130] & b[33])^(a[129] & b[34])^(a[128] & b[35])^(a[127] & b[36])^(a[126] & b[37])^(a[125] & b[38])^(a[124] & b[39])^(a[123] & b[40])^(a[122] & b[41])^(a[121] & b[42])^(a[120] & b[43])^(a[119] & b[44])^(a[118] & b[45])^(a[117] & b[46])^(a[116] & b[47])^(a[115] & b[48])^(a[114] & b[49])^(a[113] & b[50])^(a[112] & b[51])^(a[111] & b[52])^(a[110] & b[53])^(a[109] & b[54])^(a[108] & b[55])^(a[107] & b[56])^(a[106] & b[57])^(a[105] & b[58])^(a[104] & b[59])^(a[103] & b[60])^(a[102] & b[61])^(a[101] & b[62])^(a[100] & b[63])^(a[99] & b[64])^(a[98] & b[65])^(a[97] & b[66])^(a[96] & b[67])^(a[95] & b[68])^(a[94] & b[69])^(a[93] & b[70])^(a[92] & b[71])^(a[91] & b[72])^(a[90] & b[73])^(a[89] & b[74])^(a[88] & b[75])^(a[87] & b[76])^(a[86] & b[77])^(a[85] & b[78])^(a[84] & b[79])^(a[83] & b[80])^(a[82] & b[81])^(a[81] & b[82])^(a[80] & b[83])^(a[79] & b[84])^(a[78] & b[85])^(a[77] & b[86])^(a[76] & b[87])^(a[75] & b[88])^(a[74] & b[89])^(a[73] & b[90])^(a[72] & b[91])^(a[71] & b[92])^(a[70] & b[93])^(a[69] & b[94])^(a[68] & b[95])^(a[67] & b[96])^(a[66] & b[97])^(a[65] & b[98])^(a[64] & b[99])^(a[63] & b[100])^(a[62] & b[101])^(a[61] & b[102])^(a[60] & b[103])^(a[59] & b[104])^(a[58] & b[105])^(a[57] & b[106])^(a[56] & b[107])^(a[55] & b[108])^(a[54] & b[109])^(a[53] & b[110])^(a[52] & b[111])^(a[51] & b[112])^(a[50] & b[113])^(a[49] & b[114])^(a[48] & b[115])^(a[47] & b[116])^(a[46] & b[117])^(a[45] & b[118])^(a[44] & b[119])^(a[43] & b[120])^(a[42] & b[121])^(a[41] & b[122])^(a[40] & b[123])^(a[39] & b[124])^(a[38] & b[125])^(a[37] & b[126])^(a[36] & b[127])^(a[35] & b[128])^(a[34] & b[129])^(a[33] & b[130])^(a[32] & b[131])^(a[31] & b[132])^(a[30] & b[133])^(a[29] & b[134])^(a[28] & b[135])^(a[27] & b[136])^(a[26] & b[137])^(a[25] & b[138])^(a[24] & b[139])^(a[23] & b[140])^(a[22] & b[141])^(a[21] & b[142])^(a[20] & b[143])^(a[19] & b[144])^(a[18] & b[145])^(a[17] & b[146])^(a[16] & b[147])^(a[15] & b[148])^(a[14] & b[149])^(a[13] & b[150])^(a[12] & b[151])^(a[11] & b[152])^(a[10] & b[153])^(a[9] & b[154])^(a[8] & b[155])^(a[7] & b[156])^(a[6] & b[157])^(a[5] & b[158])^(a[4] & b[159])^(a[3] & b[160])^(a[2] & b[161])^(a[1] & b[162])^(a[0] & b[163]);
assign y[164] = (a[164] & b[0])^(a[163] & b[1])^(a[162] & b[2])^(a[161] & b[3])^(a[160] & b[4])^(a[159] & b[5])^(a[158] & b[6])^(a[157] & b[7])^(a[156] & b[8])^(a[155] & b[9])^(a[154] & b[10])^(a[153] & b[11])^(a[152] & b[12])^(a[151] & b[13])^(a[150] & b[14])^(a[149] & b[15])^(a[148] & b[16])^(a[147] & b[17])^(a[146] & b[18])^(a[145] & b[19])^(a[144] & b[20])^(a[143] & b[21])^(a[142] & b[22])^(a[141] & b[23])^(a[140] & b[24])^(a[139] & b[25])^(a[138] & b[26])^(a[137] & b[27])^(a[136] & b[28])^(a[135] & b[29])^(a[134] & b[30])^(a[133] & b[31])^(a[132] & b[32])^(a[131] & b[33])^(a[130] & b[34])^(a[129] & b[35])^(a[128] & b[36])^(a[127] & b[37])^(a[126] & b[38])^(a[125] & b[39])^(a[124] & b[40])^(a[123] & b[41])^(a[122] & b[42])^(a[121] & b[43])^(a[120] & b[44])^(a[119] & b[45])^(a[118] & b[46])^(a[117] & b[47])^(a[116] & b[48])^(a[115] & b[49])^(a[114] & b[50])^(a[113] & b[51])^(a[112] & b[52])^(a[111] & b[53])^(a[110] & b[54])^(a[109] & b[55])^(a[108] & b[56])^(a[107] & b[57])^(a[106] & b[58])^(a[105] & b[59])^(a[104] & b[60])^(a[103] & b[61])^(a[102] & b[62])^(a[101] & b[63])^(a[100] & b[64])^(a[99] & b[65])^(a[98] & b[66])^(a[97] & b[67])^(a[96] & b[68])^(a[95] & b[69])^(a[94] & b[70])^(a[93] & b[71])^(a[92] & b[72])^(a[91] & b[73])^(a[90] & b[74])^(a[89] & b[75])^(a[88] & b[76])^(a[87] & b[77])^(a[86] & b[78])^(a[85] & b[79])^(a[84] & b[80])^(a[83] & b[81])^(a[82] & b[82])^(a[81] & b[83])^(a[80] & b[84])^(a[79] & b[85])^(a[78] & b[86])^(a[77] & b[87])^(a[76] & b[88])^(a[75] & b[89])^(a[74] & b[90])^(a[73] & b[91])^(a[72] & b[92])^(a[71] & b[93])^(a[70] & b[94])^(a[69] & b[95])^(a[68] & b[96])^(a[67] & b[97])^(a[66] & b[98])^(a[65] & b[99])^(a[64] & b[100])^(a[63] & b[101])^(a[62] & b[102])^(a[61] & b[103])^(a[60] & b[104])^(a[59] & b[105])^(a[58] & b[106])^(a[57] & b[107])^(a[56] & b[108])^(a[55] & b[109])^(a[54] & b[110])^(a[53] & b[111])^(a[52] & b[112])^(a[51] & b[113])^(a[50] & b[114])^(a[49] & b[115])^(a[48] & b[116])^(a[47] & b[117])^(a[46] & b[118])^(a[45] & b[119])^(a[44] & b[120])^(a[43] & b[121])^(a[42] & b[122])^(a[41] & b[123])^(a[40] & b[124])^(a[39] & b[125])^(a[38] & b[126])^(a[37] & b[127])^(a[36] & b[128])^(a[35] & b[129])^(a[34] & b[130])^(a[33] & b[131])^(a[32] & b[132])^(a[31] & b[133])^(a[30] & b[134])^(a[29] & b[135])^(a[28] & b[136])^(a[27] & b[137])^(a[26] & b[138])^(a[25] & b[139])^(a[24] & b[140])^(a[23] & b[141])^(a[22] & b[142])^(a[21] & b[143])^(a[20] & b[144])^(a[19] & b[145])^(a[18] & b[146])^(a[17] & b[147])^(a[16] & b[148])^(a[15] & b[149])^(a[14] & b[150])^(a[13] & b[151])^(a[12] & b[152])^(a[11] & b[153])^(a[10] & b[154])^(a[9] & b[155])^(a[8] & b[156])^(a[7] & b[157])^(a[6] & b[158])^(a[5] & b[159])^(a[4] & b[160])^(a[3] & b[161])^(a[2] & b[162])^(a[1] & b[163])^(a[0] & b[164]);
assign y[165] = (a[165] & b[0])^(a[164] & b[1])^(a[163] & b[2])^(a[162] & b[3])^(a[161] & b[4])^(a[160] & b[5])^(a[159] & b[6])^(a[158] & b[7])^(a[157] & b[8])^(a[156] & b[9])^(a[155] & b[10])^(a[154] & b[11])^(a[153] & b[12])^(a[152] & b[13])^(a[151] & b[14])^(a[150] & b[15])^(a[149] & b[16])^(a[148] & b[17])^(a[147] & b[18])^(a[146] & b[19])^(a[145] & b[20])^(a[144] & b[21])^(a[143] & b[22])^(a[142] & b[23])^(a[141] & b[24])^(a[140] & b[25])^(a[139] & b[26])^(a[138] & b[27])^(a[137] & b[28])^(a[136] & b[29])^(a[135] & b[30])^(a[134] & b[31])^(a[133] & b[32])^(a[132] & b[33])^(a[131] & b[34])^(a[130] & b[35])^(a[129] & b[36])^(a[128] & b[37])^(a[127] & b[38])^(a[126] & b[39])^(a[125] & b[40])^(a[124] & b[41])^(a[123] & b[42])^(a[122] & b[43])^(a[121] & b[44])^(a[120] & b[45])^(a[119] & b[46])^(a[118] & b[47])^(a[117] & b[48])^(a[116] & b[49])^(a[115] & b[50])^(a[114] & b[51])^(a[113] & b[52])^(a[112] & b[53])^(a[111] & b[54])^(a[110] & b[55])^(a[109] & b[56])^(a[108] & b[57])^(a[107] & b[58])^(a[106] & b[59])^(a[105] & b[60])^(a[104] & b[61])^(a[103] & b[62])^(a[102] & b[63])^(a[101] & b[64])^(a[100] & b[65])^(a[99] & b[66])^(a[98] & b[67])^(a[97] & b[68])^(a[96] & b[69])^(a[95] & b[70])^(a[94] & b[71])^(a[93] & b[72])^(a[92] & b[73])^(a[91] & b[74])^(a[90] & b[75])^(a[89] & b[76])^(a[88] & b[77])^(a[87] & b[78])^(a[86] & b[79])^(a[85] & b[80])^(a[84] & b[81])^(a[83] & b[82])^(a[82] & b[83])^(a[81] & b[84])^(a[80] & b[85])^(a[79] & b[86])^(a[78] & b[87])^(a[77] & b[88])^(a[76] & b[89])^(a[75] & b[90])^(a[74] & b[91])^(a[73] & b[92])^(a[72] & b[93])^(a[71] & b[94])^(a[70] & b[95])^(a[69] & b[96])^(a[68] & b[97])^(a[67] & b[98])^(a[66] & b[99])^(a[65] & b[100])^(a[64] & b[101])^(a[63] & b[102])^(a[62] & b[103])^(a[61] & b[104])^(a[60] & b[105])^(a[59] & b[106])^(a[58] & b[107])^(a[57] & b[108])^(a[56] & b[109])^(a[55] & b[110])^(a[54] & b[111])^(a[53] & b[112])^(a[52] & b[113])^(a[51] & b[114])^(a[50] & b[115])^(a[49] & b[116])^(a[48] & b[117])^(a[47] & b[118])^(a[46] & b[119])^(a[45] & b[120])^(a[44] & b[121])^(a[43] & b[122])^(a[42] & b[123])^(a[41] & b[124])^(a[40] & b[125])^(a[39] & b[126])^(a[38] & b[127])^(a[37] & b[128])^(a[36] & b[129])^(a[35] & b[130])^(a[34] & b[131])^(a[33] & b[132])^(a[32] & b[133])^(a[31] & b[134])^(a[30] & b[135])^(a[29] & b[136])^(a[28] & b[137])^(a[27] & b[138])^(a[26] & b[139])^(a[25] & b[140])^(a[24] & b[141])^(a[23] & b[142])^(a[22] & b[143])^(a[21] & b[144])^(a[20] & b[145])^(a[19] & b[146])^(a[18] & b[147])^(a[17] & b[148])^(a[16] & b[149])^(a[15] & b[150])^(a[14] & b[151])^(a[13] & b[152])^(a[12] & b[153])^(a[11] & b[154])^(a[10] & b[155])^(a[9] & b[156])^(a[8] & b[157])^(a[7] & b[158])^(a[6] & b[159])^(a[5] & b[160])^(a[4] & b[161])^(a[3] & b[162])^(a[2] & b[163])^(a[1] & b[164])^(a[0] & b[165]);
assign y[166] = (a[166] & b[0])^(a[165] & b[1])^(a[164] & b[2])^(a[163] & b[3])^(a[162] & b[4])^(a[161] & b[5])^(a[160] & b[6])^(a[159] & b[7])^(a[158] & b[8])^(a[157] & b[9])^(a[156] & b[10])^(a[155] & b[11])^(a[154] & b[12])^(a[153] & b[13])^(a[152] & b[14])^(a[151] & b[15])^(a[150] & b[16])^(a[149] & b[17])^(a[148] & b[18])^(a[147] & b[19])^(a[146] & b[20])^(a[145] & b[21])^(a[144] & b[22])^(a[143] & b[23])^(a[142] & b[24])^(a[141] & b[25])^(a[140] & b[26])^(a[139] & b[27])^(a[138] & b[28])^(a[137] & b[29])^(a[136] & b[30])^(a[135] & b[31])^(a[134] & b[32])^(a[133] & b[33])^(a[132] & b[34])^(a[131] & b[35])^(a[130] & b[36])^(a[129] & b[37])^(a[128] & b[38])^(a[127] & b[39])^(a[126] & b[40])^(a[125] & b[41])^(a[124] & b[42])^(a[123] & b[43])^(a[122] & b[44])^(a[121] & b[45])^(a[120] & b[46])^(a[119] & b[47])^(a[118] & b[48])^(a[117] & b[49])^(a[116] & b[50])^(a[115] & b[51])^(a[114] & b[52])^(a[113] & b[53])^(a[112] & b[54])^(a[111] & b[55])^(a[110] & b[56])^(a[109] & b[57])^(a[108] & b[58])^(a[107] & b[59])^(a[106] & b[60])^(a[105] & b[61])^(a[104] & b[62])^(a[103] & b[63])^(a[102] & b[64])^(a[101] & b[65])^(a[100] & b[66])^(a[99] & b[67])^(a[98] & b[68])^(a[97] & b[69])^(a[96] & b[70])^(a[95] & b[71])^(a[94] & b[72])^(a[93] & b[73])^(a[92] & b[74])^(a[91] & b[75])^(a[90] & b[76])^(a[89] & b[77])^(a[88] & b[78])^(a[87] & b[79])^(a[86] & b[80])^(a[85] & b[81])^(a[84] & b[82])^(a[83] & b[83])^(a[82] & b[84])^(a[81] & b[85])^(a[80] & b[86])^(a[79] & b[87])^(a[78] & b[88])^(a[77] & b[89])^(a[76] & b[90])^(a[75] & b[91])^(a[74] & b[92])^(a[73] & b[93])^(a[72] & b[94])^(a[71] & b[95])^(a[70] & b[96])^(a[69] & b[97])^(a[68] & b[98])^(a[67] & b[99])^(a[66] & b[100])^(a[65] & b[101])^(a[64] & b[102])^(a[63] & b[103])^(a[62] & b[104])^(a[61] & b[105])^(a[60] & b[106])^(a[59] & b[107])^(a[58] & b[108])^(a[57] & b[109])^(a[56] & b[110])^(a[55] & b[111])^(a[54] & b[112])^(a[53] & b[113])^(a[52] & b[114])^(a[51] & b[115])^(a[50] & b[116])^(a[49] & b[117])^(a[48] & b[118])^(a[47] & b[119])^(a[46] & b[120])^(a[45] & b[121])^(a[44] & b[122])^(a[43] & b[123])^(a[42] & b[124])^(a[41] & b[125])^(a[40] & b[126])^(a[39] & b[127])^(a[38] & b[128])^(a[37] & b[129])^(a[36] & b[130])^(a[35] & b[131])^(a[34] & b[132])^(a[33] & b[133])^(a[32] & b[134])^(a[31] & b[135])^(a[30] & b[136])^(a[29] & b[137])^(a[28] & b[138])^(a[27] & b[139])^(a[26] & b[140])^(a[25] & b[141])^(a[24] & b[142])^(a[23] & b[143])^(a[22] & b[144])^(a[21] & b[145])^(a[20] & b[146])^(a[19] & b[147])^(a[18] & b[148])^(a[17] & b[149])^(a[16] & b[150])^(a[15] & b[151])^(a[14] & b[152])^(a[13] & b[153])^(a[12] & b[154])^(a[11] & b[155])^(a[10] & b[156])^(a[9] & b[157])^(a[8] & b[158])^(a[7] & b[159])^(a[6] & b[160])^(a[5] & b[161])^(a[4] & b[162])^(a[3] & b[163])^(a[2] & b[164])^(a[1] & b[165])^(a[0] & b[166]);
assign y[167] = (a[167] & b[0])^(a[166] & b[1])^(a[165] & b[2])^(a[164] & b[3])^(a[163] & b[4])^(a[162] & b[5])^(a[161] & b[6])^(a[160] & b[7])^(a[159] & b[8])^(a[158] & b[9])^(a[157] & b[10])^(a[156] & b[11])^(a[155] & b[12])^(a[154] & b[13])^(a[153] & b[14])^(a[152] & b[15])^(a[151] & b[16])^(a[150] & b[17])^(a[149] & b[18])^(a[148] & b[19])^(a[147] & b[20])^(a[146] & b[21])^(a[145] & b[22])^(a[144] & b[23])^(a[143] & b[24])^(a[142] & b[25])^(a[141] & b[26])^(a[140] & b[27])^(a[139] & b[28])^(a[138] & b[29])^(a[137] & b[30])^(a[136] & b[31])^(a[135] & b[32])^(a[134] & b[33])^(a[133] & b[34])^(a[132] & b[35])^(a[131] & b[36])^(a[130] & b[37])^(a[129] & b[38])^(a[128] & b[39])^(a[127] & b[40])^(a[126] & b[41])^(a[125] & b[42])^(a[124] & b[43])^(a[123] & b[44])^(a[122] & b[45])^(a[121] & b[46])^(a[120] & b[47])^(a[119] & b[48])^(a[118] & b[49])^(a[117] & b[50])^(a[116] & b[51])^(a[115] & b[52])^(a[114] & b[53])^(a[113] & b[54])^(a[112] & b[55])^(a[111] & b[56])^(a[110] & b[57])^(a[109] & b[58])^(a[108] & b[59])^(a[107] & b[60])^(a[106] & b[61])^(a[105] & b[62])^(a[104] & b[63])^(a[103] & b[64])^(a[102] & b[65])^(a[101] & b[66])^(a[100] & b[67])^(a[99] & b[68])^(a[98] & b[69])^(a[97] & b[70])^(a[96] & b[71])^(a[95] & b[72])^(a[94] & b[73])^(a[93] & b[74])^(a[92] & b[75])^(a[91] & b[76])^(a[90] & b[77])^(a[89] & b[78])^(a[88] & b[79])^(a[87] & b[80])^(a[86] & b[81])^(a[85] & b[82])^(a[84] & b[83])^(a[83] & b[84])^(a[82] & b[85])^(a[81] & b[86])^(a[80] & b[87])^(a[79] & b[88])^(a[78] & b[89])^(a[77] & b[90])^(a[76] & b[91])^(a[75] & b[92])^(a[74] & b[93])^(a[73] & b[94])^(a[72] & b[95])^(a[71] & b[96])^(a[70] & b[97])^(a[69] & b[98])^(a[68] & b[99])^(a[67] & b[100])^(a[66] & b[101])^(a[65] & b[102])^(a[64] & b[103])^(a[63] & b[104])^(a[62] & b[105])^(a[61] & b[106])^(a[60] & b[107])^(a[59] & b[108])^(a[58] & b[109])^(a[57] & b[110])^(a[56] & b[111])^(a[55] & b[112])^(a[54] & b[113])^(a[53] & b[114])^(a[52] & b[115])^(a[51] & b[116])^(a[50] & b[117])^(a[49] & b[118])^(a[48] & b[119])^(a[47] & b[120])^(a[46] & b[121])^(a[45] & b[122])^(a[44] & b[123])^(a[43] & b[124])^(a[42] & b[125])^(a[41] & b[126])^(a[40] & b[127])^(a[39] & b[128])^(a[38] & b[129])^(a[37] & b[130])^(a[36] & b[131])^(a[35] & b[132])^(a[34] & b[133])^(a[33] & b[134])^(a[32] & b[135])^(a[31] & b[136])^(a[30] & b[137])^(a[29] & b[138])^(a[28] & b[139])^(a[27] & b[140])^(a[26] & b[141])^(a[25] & b[142])^(a[24] & b[143])^(a[23] & b[144])^(a[22] & b[145])^(a[21] & b[146])^(a[20] & b[147])^(a[19] & b[148])^(a[18] & b[149])^(a[17] & b[150])^(a[16] & b[151])^(a[15] & b[152])^(a[14] & b[153])^(a[13] & b[154])^(a[12] & b[155])^(a[11] & b[156])^(a[10] & b[157])^(a[9] & b[158])^(a[8] & b[159])^(a[7] & b[160])^(a[6] & b[161])^(a[5] & b[162])^(a[4] & b[163])^(a[3] & b[164])^(a[2] & b[165])^(a[1] & b[166])^(a[0] & b[167]);
assign y[168] = (a[168] & b[0])^(a[167] & b[1])^(a[166] & b[2])^(a[165] & b[3])^(a[164] & b[4])^(a[163] & b[5])^(a[162] & b[6])^(a[161] & b[7])^(a[160] & b[8])^(a[159] & b[9])^(a[158] & b[10])^(a[157] & b[11])^(a[156] & b[12])^(a[155] & b[13])^(a[154] & b[14])^(a[153] & b[15])^(a[152] & b[16])^(a[151] & b[17])^(a[150] & b[18])^(a[149] & b[19])^(a[148] & b[20])^(a[147] & b[21])^(a[146] & b[22])^(a[145] & b[23])^(a[144] & b[24])^(a[143] & b[25])^(a[142] & b[26])^(a[141] & b[27])^(a[140] & b[28])^(a[139] & b[29])^(a[138] & b[30])^(a[137] & b[31])^(a[136] & b[32])^(a[135] & b[33])^(a[134] & b[34])^(a[133] & b[35])^(a[132] & b[36])^(a[131] & b[37])^(a[130] & b[38])^(a[129] & b[39])^(a[128] & b[40])^(a[127] & b[41])^(a[126] & b[42])^(a[125] & b[43])^(a[124] & b[44])^(a[123] & b[45])^(a[122] & b[46])^(a[121] & b[47])^(a[120] & b[48])^(a[119] & b[49])^(a[118] & b[50])^(a[117] & b[51])^(a[116] & b[52])^(a[115] & b[53])^(a[114] & b[54])^(a[113] & b[55])^(a[112] & b[56])^(a[111] & b[57])^(a[110] & b[58])^(a[109] & b[59])^(a[108] & b[60])^(a[107] & b[61])^(a[106] & b[62])^(a[105] & b[63])^(a[104] & b[64])^(a[103] & b[65])^(a[102] & b[66])^(a[101] & b[67])^(a[100] & b[68])^(a[99] & b[69])^(a[98] & b[70])^(a[97] & b[71])^(a[96] & b[72])^(a[95] & b[73])^(a[94] & b[74])^(a[93] & b[75])^(a[92] & b[76])^(a[91] & b[77])^(a[90] & b[78])^(a[89] & b[79])^(a[88] & b[80])^(a[87] & b[81])^(a[86] & b[82])^(a[85] & b[83])^(a[84] & b[84])^(a[83] & b[85])^(a[82] & b[86])^(a[81] & b[87])^(a[80] & b[88])^(a[79] & b[89])^(a[78] & b[90])^(a[77] & b[91])^(a[76] & b[92])^(a[75] & b[93])^(a[74] & b[94])^(a[73] & b[95])^(a[72] & b[96])^(a[71] & b[97])^(a[70] & b[98])^(a[69] & b[99])^(a[68] & b[100])^(a[67] & b[101])^(a[66] & b[102])^(a[65] & b[103])^(a[64] & b[104])^(a[63] & b[105])^(a[62] & b[106])^(a[61] & b[107])^(a[60] & b[108])^(a[59] & b[109])^(a[58] & b[110])^(a[57] & b[111])^(a[56] & b[112])^(a[55] & b[113])^(a[54] & b[114])^(a[53] & b[115])^(a[52] & b[116])^(a[51] & b[117])^(a[50] & b[118])^(a[49] & b[119])^(a[48] & b[120])^(a[47] & b[121])^(a[46] & b[122])^(a[45] & b[123])^(a[44] & b[124])^(a[43] & b[125])^(a[42] & b[126])^(a[41] & b[127])^(a[40] & b[128])^(a[39] & b[129])^(a[38] & b[130])^(a[37] & b[131])^(a[36] & b[132])^(a[35] & b[133])^(a[34] & b[134])^(a[33] & b[135])^(a[32] & b[136])^(a[31] & b[137])^(a[30] & b[138])^(a[29] & b[139])^(a[28] & b[140])^(a[27] & b[141])^(a[26] & b[142])^(a[25] & b[143])^(a[24] & b[144])^(a[23] & b[145])^(a[22] & b[146])^(a[21] & b[147])^(a[20] & b[148])^(a[19] & b[149])^(a[18] & b[150])^(a[17] & b[151])^(a[16] & b[152])^(a[15] & b[153])^(a[14] & b[154])^(a[13] & b[155])^(a[12] & b[156])^(a[11] & b[157])^(a[10] & b[158])^(a[9] & b[159])^(a[8] & b[160])^(a[7] & b[161])^(a[6] & b[162])^(a[5] & b[163])^(a[4] & b[164])^(a[3] & b[165])^(a[2] & b[166])^(a[1] & b[167])^(a[0] & b[168]);
assign y[169] = (a[169] & b[0])^(a[168] & b[1])^(a[167] & b[2])^(a[166] & b[3])^(a[165] & b[4])^(a[164] & b[5])^(a[163] & b[6])^(a[162] & b[7])^(a[161] & b[8])^(a[160] & b[9])^(a[159] & b[10])^(a[158] & b[11])^(a[157] & b[12])^(a[156] & b[13])^(a[155] & b[14])^(a[154] & b[15])^(a[153] & b[16])^(a[152] & b[17])^(a[151] & b[18])^(a[150] & b[19])^(a[149] & b[20])^(a[148] & b[21])^(a[147] & b[22])^(a[146] & b[23])^(a[145] & b[24])^(a[144] & b[25])^(a[143] & b[26])^(a[142] & b[27])^(a[141] & b[28])^(a[140] & b[29])^(a[139] & b[30])^(a[138] & b[31])^(a[137] & b[32])^(a[136] & b[33])^(a[135] & b[34])^(a[134] & b[35])^(a[133] & b[36])^(a[132] & b[37])^(a[131] & b[38])^(a[130] & b[39])^(a[129] & b[40])^(a[128] & b[41])^(a[127] & b[42])^(a[126] & b[43])^(a[125] & b[44])^(a[124] & b[45])^(a[123] & b[46])^(a[122] & b[47])^(a[121] & b[48])^(a[120] & b[49])^(a[119] & b[50])^(a[118] & b[51])^(a[117] & b[52])^(a[116] & b[53])^(a[115] & b[54])^(a[114] & b[55])^(a[113] & b[56])^(a[112] & b[57])^(a[111] & b[58])^(a[110] & b[59])^(a[109] & b[60])^(a[108] & b[61])^(a[107] & b[62])^(a[106] & b[63])^(a[105] & b[64])^(a[104] & b[65])^(a[103] & b[66])^(a[102] & b[67])^(a[101] & b[68])^(a[100] & b[69])^(a[99] & b[70])^(a[98] & b[71])^(a[97] & b[72])^(a[96] & b[73])^(a[95] & b[74])^(a[94] & b[75])^(a[93] & b[76])^(a[92] & b[77])^(a[91] & b[78])^(a[90] & b[79])^(a[89] & b[80])^(a[88] & b[81])^(a[87] & b[82])^(a[86] & b[83])^(a[85] & b[84])^(a[84] & b[85])^(a[83] & b[86])^(a[82] & b[87])^(a[81] & b[88])^(a[80] & b[89])^(a[79] & b[90])^(a[78] & b[91])^(a[77] & b[92])^(a[76] & b[93])^(a[75] & b[94])^(a[74] & b[95])^(a[73] & b[96])^(a[72] & b[97])^(a[71] & b[98])^(a[70] & b[99])^(a[69] & b[100])^(a[68] & b[101])^(a[67] & b[102])^(a[66] & b[103])^(a[65] & b[104])^(a[64] & b[105])^(a[63] & b[106])^(a[62] & b[107])^(a[61] & b[108])^(a[60] & b[109])^(a[59] & b[110])^(a[58] & b[111])^(a[57] & b[112])^(a[56] & b[113])^(a[55] & b[114])^(a[54] & b[115])^(a[53] & b[116])^(a[52] & b[117])^(a[51] & b[118])^(a[50] & b[119])^(a[49] & b[120])^(a[48] & b[121])^(a[47] & b[122])^(a[46] & b[123])^(a[45] & b[124])^(a[44] & b[125])^(a[43] & b[126])^(a[42] & b[127])^(a[41] & b[128])^(a[40] & b[129])^(a[39] & b[130])^(a[38] & b[131])^(a[37] & b[132])^(a[36] & b[133])^(a[35] & b[134])^(a[34] & b[135])^(a[33] & b[136])^(a[32] & b[137])^(a[31] & b[138])^(a[30] & b[139])^(a[29] & b[140])^(a[28] & b[141])^(a[27] & b[142])^(a[26] & b[143])^(a[25] & b[144])^(a[24] & b[145])^(a[23] & b[146])^(a[22] & b[147])^(a[21] & b[148])^(a[20] & b[149])^(a[19] & b[150])^(a[18] & b[151])^(a[17] & b[152])^(a[16] & b[153])^(a[15] & b[154])^(a[14] & b[155])^(a[13] & b[156])^(a[12] & b[157])^(a[11] & b[158])^(a[10] & b[159])^(a[9] & b[160])^(a[8] & b[161])^(a[7] & b[162])^(a[6] & b[163])^(a[5] & b[164])^(a[4] & b[165])^(a[3] & b[166])^(a[2] & b[167])^(a[1] & b[168])^(a[0] & b[169]);
assign y[170] = (a[170] & b[0])^(a[169] & b[1])^(a[168] & b[2])^(a[167] & b[3])^(a[166] & b[4])^(a[165] & b[5])^(a[164] & b[6])^(a[163] & b[7])^(a[162] & b[8])^(a[161] & b[9])^(a[160] & b[10])^(a[159] & b[11])^(a[158] & b[12])^(a[157] & b[13])^(a[156] & b[14])^(a[155] & b[15])^(a[154] & b[16])^(a[153] & b[17])^(a[152] & b[18])^(a[151] & b[19])^(a[150] & b[20])^(a[149] & b[21])^(a[148] & b[22])^(a[147] & b[23])^(a[146] & b[24])^(a[145] & b[25])^(a[144] & b[26])^(a[143] & b[27])^(a[142] & b[28])^(a[141] & b[29])^(a[140] & b[30])^(a[139] & b[31])^(a[138] & b[32])^(a[137] & b[33])^(a[136] & b[34])^(a[135] & b[35])^(a[134] & b[36])^(a[133] & b[37])^(a[132] & b[38])^(a[131] & b[39])^(a[130] & b[40])^(a[129] & b[41])^(a[128] & b[42])^(a[127] & b[43])^(a[126] & b[44])^(a[125] & b[45])^(a[124] & b[46])^(a[123] & b[47])^(a[122] & b[48])^(a[121] & b[49])^(a[120] & b[50])^(a[119] & b[51])^(a[118] & b[52])^(a[117] & b[53])^(a[116] & b[54])^(a[115] & b[55])^(a[114] & b[56])^(a[113] & b[57])^(a[112] & b[58])^(a[111] & b[59])^(a[110] & b[60])^(a[109] & b[61])^(a[108] & b[62])^(a[107] & b[63])^(a[106] & b[64])^(a[105] & b[65])^(a[104] & b[66])^(a[103] & b[67])^(a[102] & b[68])^(a[101] & b[69])^(a[100] & b[70])^(a[99] & b[71])^(a[98] & b[72])^(a[97] & b[73])^(a[96] & b[74])^(a[95] & b[75])^(a[94] & b[76])^(a[93] & b[77])^(a[92] & b[78])^(a[91] & b[79])^(a[90] & b[80])^(a[89] & b[81])^(a[88] & b[82])^(a[87] & b[83])^(a[86] & b[84])^(a[85] & b[85])^(a[84] & b[86])^(a[83] & b[87])^(a[82] & b[88])^(a[81] & b[89])^(a[80] & b[90])^(a[79] & b[91])^(a[78] & b[92])^(a[77] & b[93])^(a[76] & b[94])^(a[75] & b[95])^(a[74] & b[96])^(a[73] & b[97])^(a[72] & b[98])^(a[71] & b[99])^(a[70] & b[100])^(a[69] & b[101])^(a[68] & b[102])^(a[67] & b[103])^(a[66] & b[104])^(a[65] & b[105])^(a[64] & b[106])^(a[63] & b[107])^(a[62] & b[108])^(a[61] & b[109])^(a[60] & b[110])^(a[59] & b[111])^(a[58] & b[112])^(a[57] & b[113])^(a[56] & b[114])^(a[55] & b[115])^(a[54] & b[116])^(a[53] & b[117])^(a[52] & b[118])^(a[51] & b[119])^(a[50] & b[120])^(a[49] & b[121])^(a[48] & b[122])^(a[47] & b[123])^(a[46] & b[124])^(a[45] & b[125])^(a[44] & b[126])^(a[43] & b[127])^(a[42] & b[128])^(a[41] & b[129])^(a[40] & b[130])^(a[39] & b[131])^(a[38] & b[132])^(a[37] & b[133])^(a[36] & b[134])^(a[35] & b[135])^(a[34] & b[136])^(a[33] & b[137])^(a[32] & b[138])^(a[31] & b[139])^(a[30] & b[140])^(a[29] & b[141])^(a[28] & b[142])^(a[27] & b[143])^(a[26] & b[144])^(a[25] & b[145])^(a[24] & b[146])^(a[23] & b[147])^(a[22] & b[148])^(a[21] & b[149])^(a[20] & b[150])^(a[19] & b[151])^(a[18] & b[152])^(a[17] & b[153])^(a[16] & b[154])^(a[15] & b[155])^(a[14] & b[156])^(a[13] & b[157])^(a[12] & b[158])^(a[11] & b[159])^(a[10] & b[160])^(a[9] & b[161])^(a[8] & b[162])^(a[7] & b[163])^(a[6] & b[164])^(a[5] & b[165])^(a[4] & b[166])^(a[3] & b[167])^(a[2] & b[168])^(a[1] & b[169])^(a[0] & b[170]);
assign y[171] = (a[171] & b[0])^(a[170] & b[1])^(a[169] & b[2])^(a[168] & b[3])^(a[167] & b[4])^(a[166] & b[5])^(a[165] & b[6])^(a[164] & b[7])^(a[163] & b[8])^(a[162] & b[9])^(a[161] & b[10])^(a[160] & b[11])^(a[159] & b[12])^(a[158] & b[13])^(a[157] & b[14])^(a[156] & b[15])^(a[155] & b[16])^(a[154] & b[17])^(a[153] & b[18])^(a[152] & b[19])^(a[151] & b[20])^(a[150] & b[21])^(a[149] & b[22])^(a[148] & b[23])^(a[147] & b[24])^(a[146] & b[25])^(a[145] & b[26])^(a[144] & b[27])^(a[143] & b[28])^(a[142] & b[29])^(a[141] & b[30])^(a[140] & b[31])^(a[139] & b[32])^(a[138] & b[33])^(a[137] & b[34])^(a[136] & b[35])^(a[135] & b[36])^(a[134] & b[37])^(a[133] & b[38])^(a[132] & b[39])^(a[131] & b[40])^(a[130] & b[41])^(a[129] & b[42])^(a[128] & b[43])^(a[127] & b[44])^(a[126] & b[45])^(a[125] & b[46])^(a[124] & b[47])^(a[123] & b[48])^(a[122] & b[49])^(a[121] & b[50])^(a[120] & b[51])^(a[119] & b[52])^(a[118] & b[53])^(a[117] & b[54])^(a[116] & b[55])^(a[115] & b[56])^(a[114] & b[57])^(a[113] & b[58])^(a[112] & b[59])^(a[111] & b[60])^(a[110] & b[61])^(a[109] & b[62])^(a[108] & b[63])^(a[107] & b[64])^(a[106] & b[65])^(a[105] & b[66])^(a[104] & b[67])^(a[103] & b[68])^(a[102] & b[69])^(a[101] & b[70])^(a[100] & b[71])^(a[99] & b[72])^(a[98] & b[73])^(a[97] & b[74])^(a[96] & b[75])^(a[95] & b[76])^(a[94] & b[77])^(a[93] & b[78])^(a[92] & b[79])^(a[91] & b[80])^(a[90] & b[81])^(a[89] & b[82])^(a[88] & b[83])^(a[87] & b[84])^(a[86] & b[85])^(a[85] & b[86])^(a[84] & b[87])^(a[83] & b[88])^(a[82] & b[89])^(a[81] & b[90])^(a[80] & b[91])^(a[79] & b[92])^(a[78] & b[93])^(a[77] & b[94])^(a[76] & b[95])^(a[75] & b[96])^(a[74] & b[97])^(a[73] & b[98])^(a[72] & b[99])^(a[71] & b[100])^(a[70] & b[101])^(a[69] & b[102])^(a[68] & b[103])^(a[67] & b[104])^(a[66] & b[105])^(a[65] & b[106])^(a[64] & b[107])^(a[63] & b[108])^(a[62] & b[109])^(a[61] & b[110])^(a[60] & b[111])^(a[59] & b[112])^(a[58] & b[113])^(a[57] & b[114])^(a[56] & b[115])^(a[55] & b[116])^(a[54] & b[117])^(a[53] & b[118])^(a[52] & b[119])^(a[51] & b[120])^(a[50] & b[121])^(a[49] & b[122])^(a[48] & b[123])^(a[47] & b[124])^(a[46] & b[125])^(a[45] & b[126])^(a[44] & b[127])^(a[43] & b[128])^(a[42] & b[129])^(a[41] & b[130])^(a[40] & b[131])^(a[39] & b[132])^(a[38] & b[133])^(a[37] & b[134])^(a[36] & b[135])^(a[35] & b[136])^(a[34] & b[137])^(a[33] & b[138])^(a[32] & b[139])^(a[31] & b[140])^(a[30] & b[141])^(a[29] & b[142])^(a[28] & b[143])^(a[27] & b[144])^(a[26] & b[145])^(a[25] & b[146])^(a[24] & b[147])^(a[23] & b[148])^(a[22] & b[149])^(a[21] & b[150])^(a[20] & b[151])^(a[19] & b[152])^(a[18] & b[153])^(a[17] & b[154])^(a[16] & b[155])^(a[15] & b[156])^(a[14] & b[157])^(a[13] & b[158])^(a[12] & b[159])^(a[11] & b[160])^(a[10] & b[161])^(a[9] & b[162])^(a[8] & b[163])^(a[7] & b[164])^(a[6] & b[165])^(a[5] & b[166])^(a[4] & b[167])^(a[3] & b[168])^(a[2] & b[169])^(a[1] & b[170])^(a[0] & b[171]);
assign y[172] = (a[172] & b[0])^(a[171] & b[1])^(a[170] & b[2])^(a[169] & b[3])^(a[168] & b[4])^(a[167] & b[5])^(a[166] & b[6])^(a[165] & b[7])^(a[164] & b[8])^(a[163] & b[9])^(a[162] & b[10])^(a[161] & b[11])^(a[160] & b[12])^(a[159] & b[13])^(a[158] & b[14])^(a[157] & b[15])^(a[156] & b[16])^(a[155] & b[17])^(a[154] & b[18])^(a[153] & b[19])^(a[152] & b[20])^(a[151] & b[21])^(a[150] & b[22])^(a[149] & b[23])^(a[148] & b[24])^(a[147] & b[25])^(a[146] & b[26])^(a[145] & b[27])^(a[144] & b[28])^(a[143] & b[29])^(a[142] & b[30])^(a[141] & b[31])^(a[140] & b[32])^(a[139] & b[33])^(a[138] & b[34])^(a[137] & b[35])^(a[136] & b[36])^(a[135] & b[37])^(a[134] & b[38])^(a[133] & b[39])^(a[132] & b[40])^(a[131] & b[41])^(a[130] & b[42])^(a[129] & b[43])^(a[128] & b[44])^(a[127] & b[45])^(a[126] & b[46])^(a[125] & b[47])^(a[124] & b[48])^(a[123] & b[49])^(a[122] & b[50])^(a[121] & b[51])^(a[120] & b[52])^(a[119] & b[53])^(a[118] & b[54])^(a[117] & b[55])^(a[116] & b[56])^(a[115] & b[57])^(a[114] & b[58])^(a[113] & b[59])^(a[112] & b[60])^(a[111] & b[61])^(a[110] & b[62])^(a[109] & b[63])^(a[108] & b[64])^(a[107] & b[65])^(a[106] & b[66])^(a[105] & b[67])^(a[104] & b[68])^(a[103] & b[69])^(a[102] & b[70])^(a[101] & b[71])^(a[100] & b[72])^(a[99] & b[73])^(a[98] & b[74])^(a[97] & b[75])^(a[96] & b[76])^(a[95] & b[77])^(a[94] & b[78])^(a[93] & b[79])^(a[92] & b[80])^(a[91] & b[81])^(a[90] & b[82])^(a[89] & b[83])^(a[88] & b[84])^(a[87] & b[85])^(a[86] & b[86])^(a[85] & b[87])^(a[84] & b[88])^(a[83] & b[89])^(a[82] & b[90])^(a[81] & b[91])^(a[80] & b[92])^(a[79] & b[93])^(a[78] & b[94])^(a[77] & b[95])^(a[76] & b[96])^(a[75] & b[97])^(a[74] & b[98])^(a[73] & b[99])^(a[72] & b[100])^(a[71] & b[101])^(a[70] & b[102])^(a[69] & b[103])^(a[68] & b[104])^(a[67] & b[105])^(a[66] & b[106])^(a[65] & b[107])^(a[64] & b[108])^(a[63] & b[109])^(a[62] & b[110])^(a[61] & b[111])^(a[60] & b[112])^(a[59] & b[113])^(a[58] & b[114])^(a[57] & b[115])^(a[56] & b[116])^(a[55] & b[117])^(a[54] & b[118])^(a[53] & b[119])^(a[52] & b[120])^(a[51] & b[121])^(a[50] & b[122])^(a[49] & b[123])^(a[48] & b[124])^(a[47] & b[125])^(a[46] & b[126])^(a[45] & b[127])^(a[44] & b[128])^(a[43] & b[129])^(a[42] & b[130])^(a[41] & b[131])^(a[40] & b[132])^(a[39] & b[133])^(a[38] & b[134])^(a[37] & b[135])^(a[36] & b[136])^(a[35] & b[137])^(a[34] & b[138])^(a[33] & b[139])^(a[32] & b[140])^(a[31] & b[141])^(a[30] & b[142])^(a[29] & b[143])^(a[28] & b[144])^(a[27] & b[145])^(a[26] & b[146])^(a[25] & b[147])^(a[24] & b[148])^(a[23] & b[149])^(a[22] & b[150])^(a[21] & b[151])^(a[20] & b[152])^(a[19] & b[153])^(a[18] & b[154])^(a[17] & b[155])^(a[16] & b[156])^(a[15] & b[157])^(a[14] & b[158])^(a[13] & b[159])^(a[12] & b[160])^(a[11] & b[161])^(a[10] & b[162])^(a[9] & b[163])^(a[8] & b[164])^(a[7] & b[165])^(a[6] & b[166])^(a[5] & b[167])^(a[4] & b[168])^(a[3] & b[169])^(a[2] & b[170])^(a[1] & b[171])^(a[0] & b[172]);
assign y[173] = (a[173] & b[0])^(a[172] & b[1])^(a[171] & b[2])^(a[170] & b[3])^(a[169] & b[4])^(a[168] & b[5])^(a[167] & b[6])^(a[166] & b[7])^(a[165] & b[8])^(a[164] & b[9])^(a[163] & b[10])^(a[162] & b[11])^(a[161] & b[12])^(a[160] & b[13])^(a[159] & b[14])^(a[158] & b[15])^(a[157] & b[16])^(a[156] & b[17])^(a[155] & b[18])^(a[154] & b[19])^(a[153] & b[20])^(a[152] & b[21])^(a[151] & b[22])^(a[150] & b[23])^(a[149] & b[24])^(a[148] & b[25])^(a[147] & b[26])^(a[146] & b[27])^(a[145] & b[28])^(a[144] & b[29])^(a[143] & b[30])^(a[142] & b[31])^(a[141] & b[32])^(a[140] & b[33])^(a[139] & b[34])^(a[138] & b[35])^(a[137] & b[36])^(a[136] & b[37])^(a[135] & b[38])^(a[134] & b[39])^(a[133] & b[40])^(a[132] & b[41])^(a[131] & b[42])^(a[130] & b[43])^(a[129] & b[44])^(a[128] & b[45])^(a[127] & b[46])^(a[126] & b[47])^(a[125] & b[48])^(a[124] & b[49])^(a[123] & b[50])^(a[122] & b[51])^(a[121] & b[52])^(a[120] & b[53])^(a[119] & b[54])^(a[118] & b[55])^(a[117] & b[56])^(a[116] & b[57])^(a[115] & b[58])^(a[114] & b[59])^(a[113] & b[60])^(a[112] & b[61])^(a[111] & b[62])^(a[110] & b[63])^(a[109] & b[64])^(a[108] & b[65])^(a[107] & b[66])^(a[106] & b[67])^(a[105] & b[68])^(a[104] & b[69])^(a[103] & b[70])^(a[102] & b[71])^(a[101] & b[72])^(a[100] & b[73])^(a[99] & b[74])^(a[98] & b[75])^(a[97] & b[76])^(a[96] & b[77])^(a[95] & b[78])^(a[94] & b[79])^(a[93] & b[80])^(a[92] & b[81])^(a[91] & b[82])^(a[90] & b[83])^(a[89] & b[84])^(a[88] & b[85])^(a[87] & b[86])^(a[86] & b[87])^(a[85] & b[88])^(a[84] & b[89])^(a[83] & b[90])^(a[82] & b[91])^(a[81] & b[92])^(a[80] & b[93])^(a[79] & b[94])^(a[78] & b[95])^(a[77] & b[96])^(a[76] & b[97])^(a[75] & b[98])^(a[74] & b[99])^(a[73] & b[100])^(a[72] & b[101])^(a[71] & b[102])^(a[70] & b[103])^(a[69] & b[104])^(a[68] & b[105])^(a[67] & b[106])^(a[66] & b[107])^(a[65] & b[108])^(a[64] & b[109])^(a[63] & b[110])^(a[62] & b[111])^(a[61] & b[112])^(a[60] & b[113])^(a[59] & b[114])^(a[58] & b[115])^(a[57] & b[116])^(a[56] & b[117])^(a[55] & b[118])^(a[54] & b[119])^(a[53] & b[120])^(a[52] & b[121])^(a[51] & b[122])^(a[50] & b[123])^(a[49] & b[124])^(a[48] & b[125])^(a[47] & b[126])^(a[46] & b[127])^(a[45] & b[128])^(a[44] & b[129])^(a[43] & b[130])^(a[42] & b[131])^(a[41] & b[132])^(a[40] & b[133])^(a[39] & b[134])^(a[38] & b[135])^(a[37] & b[136])^(a[36] & b[137])^(a[35] & b[138])^(a[34] & b[139])^(a[33] & b[140])^(a[32] & b[141])^(a[31] & b[142])^(a[30] & b[143])^(a[29] & b[144])^(a[28] & b[145])^(a[27] & b[146])^(a[26] & b[147])^(a[25] & b[148])^(a[24] & b[149])^(a[23] & b[150])^(a[22] & b[151])^(a[21] & b[152])^(a[20] & b[153])^(a[19] & b[154])^(a[18] & b[155])^(a[17] & b[156])^(a[16] & b[157])^(a[15] & b[158])^(a[14] & b[159])^(a[13] & b[160])^(a[12] & b[161])^(a[11] & b[162])^(a[10] & b[163])^(a[9] & b[164])^(a[8] & b[165])^(a[7] & b[166])^(a[6] & b[167])^(a[5] & b[168])^(a[4] & b[169])^(a[3] & b[170])^(a[2] & b[171])^(a[1] & b[172])^(a[0] & b[173]);
assign y[174] = (a[174] & b[0])^(a[173] & b[1])^(a[172] & b[2])^(a[171] & b[3])^(a[170] & b[4])^(a[169] & b[5])^(a[168] & b[6])^(a[167] & b[7])^(a[166] & b[8])^(a[165] & b[9])^(a[164] & b[10])^(a[163] & b[11])^(a[162] & b[12])^(a[161] & b[13])^(a[160] & b[14])^(a[159] & b[15])^(a[158] & b[16])^(a[157] & b[17])^(a[156] & b[18])^(a[155] & b[19])^(a[154] & b[20])^(a[153] & b[21])^(a[152] & b[22])^(a[151] & b[23])^(a[150] & b[24])^(a[149] & b[25])^(a[148] & b[26])^(a[147] & b[27])^(a[146] & b[28])^(a[145] & b[29])^(a[144] & b[30])^(a[143] & b[31])^(a[142] & b[32])^(a[141] & b[33])^(a[140] & b[34])^(a[139] & b[35])^(a[138] & b[36])^(a[137] & b[37])^(a[136] & b[38])^(a[135] & b[39])^(a[134] & b[40])^(a[133] & b[41])^(a[132] & b[42])^(a[131] & b[43])^(a[130] & b[44])^(a[129] & b[45])^(a[128] & b[46])^(a[127] & b[47])^(a[126] & b[48])^(a[125] & b[49])^(a[124] & b[50])^(a[123] & b[51])^(a[122] & b[52])^(a[121] & b[53])^(a[120] & b[54])^(a[119] & b[55])^(a[118] & b[56])^(a[117] & b[57])^(a[116] & b[58])^(a[115] & b[59])^(a[114] & b[60])^(a[113] & b[61])^(a[112] & b[62])^(a[111] & b[63])^(a[110] & b[64])^(a[109] & b[65])^(a[108] & b[66])^(a[107] & b[67])^(a[106] & b[68])^(a[105] & b[69])^(a[104] & b[70])^(a[103] & b[71])^(a[102] & b[72])^(a[101] & b[73])^(a[100] & b[74])^(a[99] & b[75])^(a[98] & b[76])^(a[97] & b[77])^(a[96] & b[78])^(a[95] & b[79])^(a[94] & b[80])^(a[93] & b[81])^(a[92] & b[82])^(a[91] & b[83])^(a[90] & b[84])^(a[89] & b[85])^(a[88] & b[86])^(a[87] & b[87])^(a[86] & b[88])^(a[85] & b[89])^(a[84] & b[90])^(a[83] & b[91])^(a[82] & b[92])^(a[81] & b[93])^(a[80] & b[94])^(a[79] & b[95])^(a[78] & b[96])^(a[77] & b[97])^(a[76] & b[98])^(a[75] & b[99])^(a[74] & b[100])^(a[73] & b[101])^(a[72] & b[102])^(a[71] & b[103])^(a[70] & b[104])^(a[69] & b[105])^(a[68] & b[106])^(a[67] & b[107])^(a[66] & b[108])^(a[65] & b[109])^(a[64] & b[110])^(a[63] & b[111])^(a[62] & b[112])^(a[61] & b[113])^(a[60] & b[114])^(a[59] & b[115])^(a[58] & b[116])^(a[57] & b[117])^(a[56] & b[118])^(a[55] & b[119])^(a[54] & b[120])^(a[53] & b[121])^(a[52] & b[122])^(a[51] & b[123])^(a[50] & b[124])^(a[49] & b[125])^(a[48] & b[126])^(a[47] & b[127])^(a[46] & b[128])^(a[45] & b[129])^(a[44] & b[130])^(a[43] & b[131])^(a[42] & b[132])^(a[41] & b[133])^(a[40] & b[134])^(a[39] & b[135])^(a[38] & b[136])^(a[37] & b[137])^(a[36] & b[138])^(a[35] & b[139])^(a[34] & b[140])^(a[33] & b[141])^(a[32] & b[142])^(a[31] & b[143])^(a[30] & b[144])^(a[29] & b[145])^(a[28] & b[146])^(a[27] & b[147])^(a[26] & b[148])^(a[25] & b[149])^(a[24] & b[150])^(a[23] & b[151])^(a[22] & b[152])^(a[21] & b[153])^(a[20] & b[154])^(a[19] & b[155])^(a[18] & b[156])^(a[17] & b[157])^(a[16] & b[158])^(a[15] & b[159])^(a[14] & b[160])^(a[13] & b[161])^(a[12] & b[162])^(a[11] & b[163])^(a[10] & b[164])^(a[9] & b[165])^(a[8] & b[166])^(a[7] & b[167])^(a[6] & b[168])^(a[5] & b[169])^(a[4] & b[170])^(a[3] & b[171])^(a[2] & b[172])^(a[1] & b[173])^(a[0] & b[174]);
assign y[175] = (a[175] & b[0])^(a[174] & b[1])^(a[173] & b[2])^(a[172] & b[3])^(a[171] & b[4])^(a[170] & b[5])^(a[169] & b[6])^(a[168] & b[7])^(a[167] & b[8])^(a[166] & b[9])^(a[165] & b[10])^(a[164] & b[11])^(a[163] & b[12])^(a[162] & b[13])^(a[161] & b[14])^(a[160] & b[15])^(a[159] & b[16])^(a[158] & b[17])^(a[157] & b[18])^(a[156] & b[19])^(a[155] & b[20])^(a[154] & b[21])^(a[153] & b[22])^(a[152] & b[23])^(a[151] & b[24])^(a[150] & b[25])^(a[149] & b[26])^(a[148] & b[27])^(a[147] & b[28])^(a[146] & b[29])^(a[145] & b[30])^(a[144] & b[31])^(a[143] & b[32])^(a[142] & b[33])^(a[141] & b[34])^(a[140] & b[35])^(a[139] & b[36])^(a[138] & b[37])^(a[137] & b[38])^(a[136] & b[39])^(a[135] & b[40])^(a[134] & b[41])^(a[133] & b[42])^(a[132] & b[43])^(a[131] & b[44])^(a[130] & b[45])^(a[129] & b[46])^(a[128] & b[47])^(a[127] & b[48])^(a[126] & b[49])^(a[125] & b[50])^(a[124] & b[51])^(a[123] & b[52])^(a[122] & b[53])^(a[121] & b[54])^(a[120] & b[55])^(a[119] & b[56])^(a[118] & b[57])^(a[117] & b[58])^(a[116] & b[59])^(a[115] & b[60])^(a[114] & b[61])^(a[113] & b[62])^(a[112] & b[63])^(a[111] & b[64])^(a[110] & b[65])^(a[109] & b[66])^(a[108] & b[67])^(a[107] & b[68])^(a[106] & b[69])^(a[105] & b[70])^(a[104] & b[71])^(a[103] & b[72])^(a[102] & b[73])^(a[101] & b[74])^(a[100] & b[75])^(a[99] & b[76])^(a[98] & b[77])^(a[97] & b[78])^(a[96] & b[79])^(a[95] & b[80])^(a[94] & b[81])^(a[93] & b[82])^(a[92] & b[83])^(a[91] & b[84])^(a[90] & b[85])^(a[89] & b[86])^(a[88] & b[87])^(a[87] & b[88])^(a[86] & b[89])^(a[85] & b[90])^(a[84] & b[91])^(a[83] & b[92])^(a[82] & b[93])^(a[81] & b[94])^(a[80] & b[95])^(a[79] & b[96])^(a[78] & b[97])^(a[77] & b[98])^(a[76] & b[99])^(a[75] & b[100])^(a[74] & b[101])^(a[73] & b[102])^(a[72] & b[103])^(a[71] & b[104])^(a[70] & b[105])^(a[69] & b[106])^(a[68] & b[107])^(a[67] & b[108])^(a[66] & b[109])^(a[65] & b[110])^(a[64] & b[111])^(a[63] & b[112])^(a[62] & b[113])^(a[61] & b[114])^(a[60] & b[115])^(a[59] & b[116])^(a[58] & b[117])^(a[57] & b[118])^(a[56] & b[119])^(a[55] & b[120])^(a[54] & b[121])^(a[53] & b[122])^(a[52] & b[123])^(a[51] & b[124])^(a[50] & b[125])^(a[49] & b[126])^(a[48] & b[127])^(a[47] & b[128])^(a[46] & b[129])^(a[45] & b[130])^(a[44] & b[131])^(a[43] & b[132])^(a[42] & b[133])^(a[41] & b[134])^(a[40] & b[135])^(a[39] & b[136])^(a[38] & b[137])^(a[37] & b[138])^(a[36] & b[139])^(a[35] & b[140])^(a[34] & b[141])^(a[33] & b[142])^(a[32] & b[143])^(a[31] & b[144])^(a[30] & b[145])^(a[29] & b[146])^(a[28] & b[147])^(a[27] & b[148])^(a[26] & b[149])^(a[25] & b[150])^(a[24] & b[151])^(a[23] & b[152])^(a[22] & b[153])^(a[21] & b[154])^(a[20] & b[155])^(a[19] & b[156])^(a[18] & b[157])^(a[17] & b[158])^(a[16] & b[159])^(a[15] & b[160])^(a[14] & b[161])^(a[13] & b[162])^(a[12] & b[163])^(a[11] & b[164])^(a[10] & b[165])^(a[9] & b[166])^(a[8] & b[167])^(a[7] & b[168])^(a[6] & b[169])^(a[5] & b[170])^(a[4] & b[171])^(a[3] & b[172])^(a[2] & b[173])^(a[1] & b[174])^(a[0] & b[175]);
assign y[176] = (a[176] & b[0])^(a[175] & b[1])^(a[174] & b[2])^(a[173] & b[3])^(a[172] & b[4])^(a[171] & b[5])^(a[170] & b[6])^(a[169] & b[7])^(a[168] & b[8])^(a[167] & b[9])^(a[166] & b[10])^(a[165] & b[11])^(a[164] & b[12])^(a[163] & b[13])^(a[162] & b[14])^(a[161] & b[15])^(a[160] & b[16])^(a[159] & b[17])^(a[158] & b[18])^(a[157] & b[19])^(a[156] & b[20])^(a[155] & b[21])^(a[154] & b[22])^(a[153] & b[23])^(a[152] & b[24])^(a[151] & b[25])^(a[150] & b[26])^(a[149] & b[27])^(a[148] & b[28])^(a[147] & b[29])^(a[146] & b[30])^(a[145] & b[31])^(a[144] & b[32])^(a[143] & b[33])^(a[142] & b[34])^(a[141] & b[35])^(a[140] & b[36])^(a[139] & b[37])^(a[138] & b[38])^(a[137] & b[39])^(a[136] & b[40])^(a[135] & b[41])^(a[134] & b[42])^(a[133] & b[43])^(a[132] & b[44])^(a[131] & b[45])^(a[130] & b[46])^(a[129] & b[47])^(a[128] & b[48])^(a[127] & b[49])^(a[126] & b[50])^(a[125] & b[51])^(a[124] & b[52])^(a[123] & b[53])^(a[122] & b[54])^(a[121] & b[55])^(a[120] & b[56])^(a[119] & b[57])^(a[118] & b[58])^(a[117] & b[59])^(a[116] & b[60])^(a[115] & b[61])^(a[114] & b[62])^(a[113] & b[63])^(a[112] & b[64])^(a[111] & b[65])^(a[110] & b[66])^(a[109] & b[67])^(a[108] & b[68])^(a[107] & b[69])^(a[106] & b[70])^(a[105] & b[71])^(a[104] & b[72])^(a[103] & b[73])^(a[102] & b[74])^(a[101] & b[75])^(a[100] & b[76])^(a[99] & b[77])^(a[98] & b[78])^(a[97] & b[79])^(a[96] & b[80])^(a[95] & b[81])^(a[94] & b[82])^(a[93] & b[83])^(a[92] & b[84])^(a[91] & b[85])^(a[90] & b[86])^(a[89] & b[87])^(a[88] & b[88])^(a[87] & b[89])^(a[86] & b[90])^(a[85] & b[91])^(a[84] & b[92])^(a[83] & b[93])^(a[82] & b[94])^(a[81] & b[95])^(a[80] & b[96])^(a[79] & b[97])^(a[78] & b[98])^(a[77] & b[99])^(a[76] & b[100])^(a[75] & b[101])^(a[74] & b[102])^(a[73] & b[103])^(a[72] & b[104])^(a[71] & b[105])^(a[70] & b[106])^(a[69] & b[107])^(a[68] & b[108])^(a[67] & b[109])^(a[66] & b[110])^(a[65] & b[111])^(a[64] & b[112])^(a[63] & b[113])^(a[62] & b[114])^(a[61] & b[115])^(a[60] & b[116])^(a[59] & b[117])^(a[58] & b[118])^(a[57] & b[119])^(a[56] & b[120])^(a[55] & b[121])^(a[54] & b[122])^(a[53] & b[123])^(a[52] & b[124])^(a[51] & b[125])^(a[50] & b[126])^(a[49] & b[127])^(a[48] & b[128])^(a[47] & b[129])^(a[46] & b[130])^(a[45] & b[131])^(a[44] & b[132])^(a[43] & b[133])^(a[42] & b[134])^(a[41] & b[135])^(a[40] & b[136])^(a[39] & b[137])^(a[38] & b[138])^(a[37] & b[139])^(a[36] & b[140])^(a[35] & b[141])^(a[34] & b[142])^(a[33] & b[143])^(a[32] & b[144])^(a[31] & b[145])^(a[30] & b[146])^(a[29] & b[147])^(a[28] & b[148])^(a[27] & b[149])^(a[26] & b[150])^(a[25] & b[151])^(a[24] & b[152])^(a[23] & b[153])^(a[22] & b[154])^(a[21] & b[155])^(a[20] & b[156])^(a[19] & b[157])^(a[18] & b[158])^(a[17] & b[159])^(a[16] & b[160])^(a[15] & b[161])^(a[14] & b[162])^(a[13] & b[163])^(a[12] & b[164])^(a[11] & b[165])^(a[10] & b[166])^(a[9] & b[167])^(a[8] & b[168])^(a[7] & b[169])^(a[6] & b[170])^(a[5] & b[171])^(a[4] & b[172])^(a[3] & b[173])^(a[2] & b[174])^(a[1] & b[175])^(a[0] & b[176]);
assign y[177] = (a[177] & b[0])^(a[176] & b[1])^(a[175] & b[2])^(a[174] & b[3])^(a[173] & b[4])^(a[172] & b[5])^(a[171] & b[6])^(a[170] & b[7])^(a[169] & b[8])^(a[168] & b[9])^(a[167] & b[10])^(a[166] & b[11])^(a[165] & b[12])^(a[164] & b[13])^(a[163] & b[14])^(a[162] & b[15])^(a[161] & b[16])^(a[160] & b[17])^(a[159] & b[18])^(a[158] & b[19])^(a[157] & b[20])^(a[156] & b[21])^(a[155] & b[22])^(a[154] & b[23])^(a[153] & b[24])^(a[152] & b[25])^(a[151] & b[26])^(a[150] & b[27])^(a[149] & b[28])^(a[148] & b[29])^(a[147] & b[30])^(a[146] & b[31])^(a[145] & b[32])^(a[144] & b[33])^(a[143] & b[34])^(a[142] & b[35])^(a[141] & b[36])^(a[140] & b[37])^(a[139] & b[38])^(a[138] & b[39])^(a[137] & b[40])^(a[136] & b[41])^(a[135] & b[42])^(a[134] & b[43])^(a[133] & b[44])^(a[132] & b[45])^(a[131] & b[46])^(a[130] & b[47])^(a[129] & b[48])^(a[128] & b[49])^(a[127] & b[50])^(a[126] & b[51])^(a[125] & b[52])^(a[124] & b[53])^(a[123] & b[54])^(a[122] & b[55])^(a[121] & b[56])^(a[120] & b[57])^(a[119] & b[58])^(a[118] & b[59])^(a[117] & b[60])^(a[116] & b[61])^(a[115] & b[62])^(a[114] & b[63])^(a[113] & b[64])^(a[112] & b[65])^(a[111] & b[66])^(a[110] & b[67])^(a[109] & b[68])^(a[108] & b[69])^(a[107] & b[70])^(a[106] & b[71])^(a[105] & b[72])^(a[104] & b[73])^(a[103] & b[74])^(a[102] & b[75])^(a[101] & b[76])^(a[100] & b[77])^(a[99] & b[78])^(a[98] & b[79])^(a[97] & b[80])^(a[96] & b[81])^(a[95] & b[82])^(a[94] & b[83])^(a[93] & b[84])^(a[92] & b[85])^(a[91] & b[86])^(a[90] & b[87])^(a[89] & b[88])^(a[88] & b[89])^(a[87] & b[90])^(a[86] & b[91])^(a[85] & b[92])^(a[84] & b[93])^(a[83] & b[94])^(a[82] & b[95])^(a[81] & b[96])^(a[80] & b[97])^(a[79] & b[98])^(a[78] & b[99])^(a[77] & b[100])^(a[76] & b[101])^(a[75] & b[102])^(a[74] & b[103])^(a[73] & b[104])^(a[72] & b[105])^(a[71] & b[106])^(a[70] & b[107])^(a[69] & b[108])^(a[68] & b[109])^(a[67] & b[110])^(a[66] & b[111])^(a[65] & b[112])^(a[64] & b[113])^(a[63] & b[114])^(a[62] & b[115])^(a[61] & b[116])^(a[60] & b[117])^(a[59] & b[118])^(a[58] & b[119])^(a[57] & b[120])^(a[56] & b[121])^(a[55] & b[122])^(a[54] & b[123])^(a[53] & b[124])^(a[52] & b[125])^(a[51] & b[126])^(a[50] & b[127])^(a[49] & b[128])^(a[48] & b[129])^(a[47] & b[130])^(a[46] & b[131])^(a[45] & b[132])^(a[44] & b[133])^(a[43] & b[134])^(a[42] & b[135])^(a[41] & b[136])^(a[40] & b[137])^(a[39] & b[138])^(a[38] & b[139])^(a[37] & b[140])^(a[36] & b[141])^(a[35] & b[142])^(a[34] & b[143])^(a[33] & b[144])^(a[32] & b[145])^(a[31] & b[146])^(a[30] & b[147])^(a[29] & b[148])^(a[28] & b[149])^(a[27] & b[150])^(a[26] & b[151])^(a[25] & b[152])^(a[24] & b[153])^(a[23] & b[154])^(a[22] & b[155])^(a[21] & b[156])^(a[20] & b[157])^(a[19] & b[158])^(a[18] & b[159])^(a[17] & b[160])^(a[16] & b[161])^(a[15] & b[162])^(a[14] & b[163])^(a[13] & b[164])^(a[12] & b[165])^(a[11] & b[166])^(a[10] & b[167])^(a[9] & b[168])^(a[8] & b[169])^(a[7] & b[170])^(a[6] & b[171])^(a[5] & b[172])^(a[4] & b[173])^(a[3] & b[174])^(a[2] & b[175])^(a[1] & b[176])^(a[0] & b[177]);
assign y[178] = (a[178] & b[0])^(a[177] & b[1])^(a[176] & b[2])^(a[175] & b[3])^(a[174] & b[4])^(a[173] & b[5])^(a[172] & b[6])^(a[171] & b[7])^(a[170] & b[8])^(a[169] & b[9])^(a[168] & b[10])^(a[167] & b[11])^(a[166] & b[12])^(a[165] & b[13])^(a[164] & b[14])^(a[163] & b[15])^(a[162] & b[16])^(a[161] & b[17])^(a[160] & b[18])^(a[159] & b[19])^(a[158] & b[20])^(a[157] & b[21])^(a[156] & b[22])^(a[155] & b[23])^(a[154] & b[24])^(a[153] & b[25])^(a[152] & b[26])^(a[151] & b[27])^(a[150] & b[28])^(a[149] & b[29])^(a[148] & b[30])^(a[147] & b[31])^(a[146] & b[32])^(a[145] & b[33])^(a[144] & b[34])^(a[143] & b[35])^(a[142] & b[36])^(a[141] & b[37])^(a[140] & b[38])^(a[139] & b[39])^(a[138] & b[40])^(a[137] & b[41])^(a[136] & b[42])^(a[135] & b[43])^(a[134] & b[44])^(a[133] & b[45])^(a[132] & b[46])^(a[131] & b[47])^(a[130] & b[48])^(a[129] & b[49])^(a[128] & b[50])^(a[127] & b[51])^(a[126] & b[52])^(a[125] & b[53])^(a[124] & b[54])^(a[123] & b[55])^(a[122] & b[56])^(a[121] & b[57])^(a[120] & b[58])^(a[119] & b[59])^(a[118] & b[60])^(a[117] & b[61])^(a[116] & b[62])^(a[115] & b[63])^(a[114] & b[64])^(a[113] & b[65])^(a[112] & b[66])^(a[111] & b[67])^(a[110] & b[68])^(a[109] & b[69])^(a[108] & b[70])^(a[107] & b[71])^(a[106] & b[72])^(a[105] & b[73])^(a[104] & b[74])^(a[103] & b[75])^(a[102] & b[76])^(a[101] & b[77])^(a[100] & b[78])^(a[99] & b[79])^(a[98] & b[80])^(a[97] & b[81])^(a[96] & b[82])^(a[95] & b[83])^(a[94] & b[84])^(a[93] & b[85])^(a[92] & b[86])^(a[91] & b[87])^(a[90] & b[88])^(a[89] & b[89])^(a[88] & b[90])^(a[87] & b[91])^(a[86] & b[92])^(a[85] & b[93])^(a[84] & b[94])^(a[83] & b[95])^(a[82] & b[96])^(a[81] & b[97])^(a[80] & b[98])^(a[79] & b[99])^(a[78] & b[100])^(a[77] & b[101])^(a[76] & b[102])^(a[75] & b[103])^(a[74] & b[104])^(a[73] & b[105])^(a[72] & b[106])^(a[71] & b[107])^(a[70] & b[108])^(a[69] & b[109])^(a[68] & b[110])^(a[67] & b[111])^(a[66] & b[112])^(a[65] & b[113])^(a[64] & b[114])^(a[63] & b[115])^(a[62] & b[116])^(a[61] & b[117])^(a[60] & b[118])^(a[59] & b[119])^(a[58] & b[120])^(a[57] & b[121])^(a[56] & b[122])^(a[55] & b[123])^(a[54] & b[124])^(a[53] & b[125])^(a[52] & b[126])^(a[51] & b[127])^(a[50] & b[128])^(a[49] & b[129])^(a[48] & b[130])^(a[47] & b[131])^(a[46] & b[132])^(a[45] & b[133])^(a[44] & b[134])^(a[43] & b[135])^(a[42] & b[136])^(a[41] & b[137])^(a[40] & b[138])^(a[39] & b[139])^(a[38] & b[140])^(a[37] & b[141])^(a[36] & b[142])^(a[35] & b[143])^(a[34] & b[144])^(a[33] & b[145])^(a[32] & b[146])^(a[31] & b[147])^(a[30] & b[148])^(a[29] & b[149])^(a[28] & b[150])^(a[27] & b[151])^(a[26] & b[152])^(a[25] & b[153])^(a[24] & b[154])^(a[23] & b[155])^(a[22] & b[156])^(a[21] & b[157])^(a[20] & b[158])^(a[19] & b[159])^(a[18] & b[160])^(a[17] & b[161])^(a[16] & b[162])^(a[15] & b[163])^(a[14] & b[164])^(a[13] & b[165])^(a[12] & b[166])^(a[11] & b[167])^(a[10] & b[168])^(a[9] & b[169])^(a[8] & b[170])^(a[7] & b[171])^(a[6] & b[172])^(a[5] & b[173])^(a[4] & b[174])^(a[3] & b[175])^(a[2] & b[176])^(a[1] & b[177])^(a[0] & b[178]);
assign y[179] = (a[179] & b[0])^(a[178] & b[1])^(a[177] & b[2])^(a[176] & b[3])^(a[175] & b[4])^(a[174] & b[5])^(a[173] & b[6])^(a[172] & b[7])^(a[171] & b[8])^(a[170] & b[9])^(a[169] & b[10])^(a[168] & b[11])^(a[167] & b[12])^(a[166] & b[13])^(a[165] & b[14])^(a[164] & b[15])^(a[163] & b[16])^(a[162] & b[17])^(a[161] & b[18])^(a[160] & b[19])^(a[159] & b[20])^(a[158] & b[21])^(a[157] & b[22])^(a[156] & b[23])^(a[155] & b[24])^(a[154] & b[25])^(a[153] & b[26])^(a[152] & b[27])^(a[151] & b[28])^(a[150] & b[29])^(a[149] & b[30])^(a[148] & b[31])^(a[147] & b[32])^(a[146] & b[33])^(a[145] & b[34])^(a[144] & b[35])^(a[143] & b[36])^(a[142] & b[37])^(a[141] & b[38])^(a[140] & b[39])^(a[139] & b[40])^(a[138] & b[41])^(a[137] & b[42])^(a[136] & b[43])^(a[135] & b[44])^(a[134] & b[45])^(a[133] & b[46])^(a[132] & b[47])^(a[131] & b[48])^(a[130] & b[49])^(a[129] & b[50])^(a[128] & b[51])^(a[127] & b[52])^(a[126] & b[53])^(a[125] & b[54])^(a[124] & b[55])^(a[123] & b[56])^(a[122] & b[57])^(a[121] & b[58])^(a[120] & b[59])^(a[119] & b[60])^(a[118] & b[61])^(a[117] & b[62])^(a[116] & b[63])^(a[115] & b[64])^(a[114] & b[65])^(a[113] & b[66])^(a[112] & b[67])^(a[111] & b[68])^(a[110] & b[69])^(a[109] & b[70])^(a[108] & b[71])^(a[107] & b[72])^(a[106] & b[73])^(a[105] & b[74])^(a[104] & b[75])^(a[103] & b[76])^(a[102] & b[77])^(a[101] & b[78])^(a[100] & b[79])^(a[99] & b[80])^(a[98] & b[81])^(a[97] & b[82])^(a[96] & b[83])^(a[95] & b[84])^(a[94] & b[85])^(a[93] & b[86])^(a[92] & b[87])^(a[91] & b[88])^(a[90] & b[89])^(a[89] & b[90])^(a[88] & b[91])^(a[87] & b[92])^(a[86] & b[93])^(a[85] & b[94])^(a[84] & b[95])^(a[83] & b[96])^(a[82] & b[97])^(a[81] & b[98])^(a[80] & b[99])^(a[79] & b[100])^(a[78] & b[101])^(a[77] & b[102])^(a[76] & b[103])^(a[75] & b[104])^(a[74] & b[105])^(a[73] & b[106])^(a[72] & b[107])^(a[71] & b[108])^(a[70] & b[109])^(a[69] & b[110])^(a[68] & b[111])^(a[67] & b[112])^(a[66] & b[113])^(a[65] & b[114])^(a[64] & b[115])^(a[63] & b[116])^(a[62] & b[117])^(a[61] & b[118])^(a[60] & b[119])^(a[59] & b[120])^(a[58] & b[121])^(a[57] & b[122])^(a[56] & b[123])^(a[55] & b[124])^(a[54] & b[125])^(a[53] & b[126])^(a[52] & b[127])^(a[51] & b[128])^(a[50] & b[129])^(a[49] & b[130])^(a[48] & b[131])^(a[47] & b[132])^(a[46] & b[133])^(a[45] & b[134])^(a[44] & b[135])^(a[43] & b[136])^(a[42] & b[137])^(a[41] & b[138])^(a[40] & b[139])^(a[39] & b[140])^(a[38] & b[141])^(a[37] & b[142])^(a[36] & b[143])^(a[35] & b[144])^(a[34] & b[145])^(a[33] & b[146])^(a[32] & b[147])^(a[31] & b[148])^(a[30] & b[149])^(a[29] & b[150])^(a[28] & b[151])^(a[27] & b[152])^(a[26] & b[153])^(a[25] & b[154])^(a[24] & b[155])^(a[23] & b[156])^(a[22] & b[157])^(a[21] & b[158])^(a[20] & b[159])^(a[19] & b[160])^(a[18] & b[161])^(a[17] & b[162])^(a[16] & b[163])^(a[15] & b[164])^(a[14] & b[165])^(a[13] & b[166])^(a[12] & b[167])^(a[11] & b[168])^(a[10] & b[169])^(a[9] & b[170])^(a[8] & b[171])^(a[7] & b[172])^(a[6] & b[173])^(a[5] & b[174])^(a[4] & b[175])^(a[3] & b[176])^(a[2] & b[177])^(a[1] & b[178])^(a[0] & b[179]);
assign y[180] = (a[180] & b[0])^(a[179] & b[1])^(a[178] & b[2])^(a[177] & b[3])^(a[176] & b[4])^(a[175] & b[5])^(a[174] & b[6])^(a[173] & b[7])^(a[172] & b[8])^(a[171] & b[9])^(a[170] & b[10])^(a[169] & b[11])^(a[168] & b[12])^(a[167] & b[13])^(a[166] & b[14])^(a[165] & b[15])^(a[164] & b[16])^(a[163] & b[17])^(a[162] & b[18])^(a[161] & b[19])^(a[160] & b[20])^(a[159] & b[21])^(a[158] & b[22])^(a[157] & b[23])^(a[156] & b[24])^(a[155] & b[25])^(a[154] & b[26])^(a[153] & b[27])^(a[152] & b[28])^(a[151] & b[29])^(a[150] & b[30])^(a[149] & b[31])^(a[148] & b[32])^(a[147] & b[33])^(a[146] & b[34])^(a[145] & b[35])^(a[144] & b[36])^(a[143] & b[37])^(a[142] & b[38])^(a[141] & b[39])^(a[140] & b[40])^(a[139] & b[41])^(a[138] & b[42])^(a[137] & b[43])^(a[136] & b[44])^(a[135] & b[45])^(a[134] & b[46])^(a[133] & b[47])^(a[132] & b[48])^(a[131] & b[49])^(a[130] & b[50])^(a[129] & b[51])^(a[128] & b[52])^(a[127] & b[53])^(a[126] & b[54])^(a[125] & b[55])^(a[124] & b[56])^(a[123] & b[57])^(a[122] & b[58])^(a[121] & b[59])^(a[120] & b[60])^(a[119] & b[61])^(a[118] & b[62])^(a[117] & b[63])^(a[116] & b[64])^(a[115] & b[65])^(a[114] & b[66])^(a[113] & b[67])^(a[112] & b[68])^(a[111] & b[69])^(a[110] & b[70])^(a[109] & b[71])^(a[108] & b[72])^(a[107] & b[73])^(a[106] & b[74])^(a[105] & b[75])^(a[104] & b[76])^(a[103] & b[77])^(a[102] & b[78])^(a[101] & b[79])^(a[100] & b[80])^(a[99] & b[81])^(a[98] & b[82])^(a[97] & b[83])^(a[96] & b[84])^(a[95] & b[85])^(a[94] & b[86])^(a[93] & b[87])^(a[92] & b[88])^(a[91] & b[89])^(a[90] & b[90])^(a[89] & b[91])^(a[88] & b[92])^(a[87] & b[93])^(a[86] & b[94])^(a[85] & b[95])^(a[84] & b[96])^(a[83] & b[97])^(a[82] & b[98])^(a[81] & b[99])^(a[80] & b[100])^(a[79] & b[101])^(a[78] & b[102])^(a[77] & b[103])^(a[76] & b[104])^(a[75] & b[105])^(a[74] & b[106])^(a[73] & b[107])^(a[72] & b[108])^(a[71] & b[109])^(a[70] & b[110])^(a[69] & b[111])^(a[68] & b[112])^(a[67] & b[113])^(a[66] & b[114])^(a[65] & b[115])^(a[64] & b[116])^(a[63] & b[117])^(a[62] & b[118])^(a[61] & b[119])^(a[60] & b[120])^(a[59] & b[121])^(a[58] & b[122])^(a[57] & b[123])^(a[56] & b[124])^(a[55] & b[125])^(a[54] & b[126])^(a[53] & b[127])^(a[52] & b[128])^(a[51] & b[129])^(a[50] & b[130])^(a[49] & b[131])^(a[48] & b[132])^(a[47] & b[133])^(a[46] & b[134])^(a[45] & b[135])^(a[44] & b[136])^(a[43] & b[137])^(a[42] & b[138])^(a[41] & b[139])^(a[40] & b[140])^(a[39] & b[141])^(a[38] & b[142])^(a[37] & b[143])^(a[36] & b[144])^(a[35] & b[145])^(a[34] & b[146])^(a[33] & b[147])^(a[32] & b[148])^(a[31] & b[149])^(a[30] & b[150])^(a[29] & b[151])^(a[28] & b[152])^(a[27] & b[153])^(a[26] & b[154])^(a[25] & b[155])^(a[24] & b[156])^(a[23] & b[157])^(a[22] & b[158])^(a[21] & b[159])^(a[20] & b[160])^(a[19] & b[161])^(a[18] & b[162])^(a[17] & b[163])^(a[16] & b[164])^(a[15] & b[165])^(a[14] & b[166])^(a[13] & b[167])^(a[12] & b[168])^(a[11] & b[169])^(a[10] & b[170])^(a[9] & b[171])^(a[8] & b[172])^(a[7] & b[173])^(a[6] & b[174])^(a[5] & b[175])^(a[4] & b[176])^(a[3] & b[177])^(a[2] & b[178])^(a[1] & b[179])^(a[0] & b[180]);
assign y[181] = (a[181] & b[0])^(a[180] & b[1])^(a[179] & b[2])^(a[178] & b[3])^(a[177] & b[4])^(a[176] & b[5])^(a[175] & b[6])^(a[174] & b[7])^(a[173] & b[8])^(a[172] & b[9])^(a[171] & b[10])^(a[170] & b[11])^(a[169] & b[12])^(a[168] & b[13])^(a[167] & b[14])^(a[166] & b[15])^(a[165] & b[16])^(a[164] & b[17])^(a[163] & b[18])^(a[162] & b[19])^(a[161] & b[20])^(a[160] & b[21])^(a[159] & b[22])^(a[158] & b[23])^(a[157] & b[24])^(a[156] & b[25])^(a[155] & b[26])^(a[154] & b[27])^(a[153] & b[28])^(a[152] & b[29])^(a[151] & b[30])^(a[150] & b[31])^(a[149] & b[32])^(a[148] & b[33])^(a[147] & b[34])^(a[146] & b[35])^(a[145] & b[36])^(a[144] & b[37])^(a[143] & b[38])^(a[142] & b[39])^(a[141] & b[40])^(a[140] & b[41])^(a[139] & b[42])^(a[138] & b[43])^(a[137] & b[44])^(a[136] & b[45])^(a[135] & b[46])^(a[134] & b[47])^(a[133] & b[48])^(a[132] & b[49])^(a[131] & b[50])^(a[130] & b[51])^(a[129] & b[52])^(a[128] & b[53])^(a[127] & b[54])^(a[126] & b[55])^(a[125] & b[56])^(a[124] & b[57])^(a[123] & b[58])^(a[122] & b[59])^(a[121] & b[60])^(a[120] & b[61])^(a[119] & b[62])^(a[118] & b[63])^(a[117] & b[64])^(a[116] & b[65])^(a[115] & b[66])^(a[114] & b[67])^(a[113] & b[68])^(a[112] & b[69])^(a[111] & b[70])^(a[110] & b[71])^(a[109] & b[72])^(a[108] & b[73])^(a[107] & b[74])^(a[106] & b[75])^(a[105] & b[76])^(a[104] & b[77])^(a[103] & b[78])^(a[102] & b[79])^(a[101] & b[80])^(a[100] & b[81])^(a[99] & b[82])^(a[98] & b[83])^(a[97] & b[84])^(a[96] & b[85])^(a[95] & b[86])^(a[94] & b[87])^(a[93] & b[88])^(a[92] & b[89])^(a[91] & b[90])^(a[90] & b[91])^(a[89] & b[92])^(a[88] & b[93])^(a[87] & b[94])^(a[86] & b[95])^(a[85] & b[96])^(a[84] & b[97])^(a[83] & b[98])^(a[82] & b[99])^(a[81] & b[100])^(a[80] & b[101])^(a[79] & b[102])^(a[78] & b[103])^(a[77] & b[104])^(a[76] & b[105])^(a[75] & b[106])^(a[74] & b[107])^(a[73] & b[108])^(a[72] & b[109])^(a[71] & b[110])^(a[70] & b[111])^(a[69] & b[112])^(a[68] & b[113])^(a[67] & b[114])^(a[66] & b[115])^(a[65] & b[116])^(a[64] & b[117])^(a[63] & b[118])^(a[62] & b[119])^(a[61] & b[120])^(a[60] & b[121])^(a[59] & b[122])^(a[58] & b[123])^(a[57] & b[124])^(a[56] & b[125])^(a[55] & b[126])^(a[54] & b[127])^(a[53] & b[128])^(a[52] & b[129])^(a[51] & b[130])^(a[50] & b[131])^(a[49] & b[132])^(a[48] & b[133])^(a[47] & b[134])^(a[46] & b[135])^(a[45] & b[136])^(a[44] & b[137])^(a[43] & b[138])^(a[42] & b[139])^(a[41] & b[140])^(a[40] & b[141])^(a[39] & b[142])^(a[38] & b[143])^(a[37] & b[144])^(a[36] & b[145])^(a[35] & b[146])^(a[34] & b[147])^(a[33] & b[148])^(a[32] & b[149])^(a[31] & b[150])^(a[30] & b[151])^(a[29] & b[152])^(a[28] & b[153])^(a[27] & b[154])^(a[26] & b[155])^(a[25] & b[156])^(a[24] & b[157])^(a[23] & b[158])^(a[22] & b[159])^(a[21] & b[160])^(a[20] & b[161])^(a[19] & b[162])^(a[18] & b[163])^(a[17] & b[164])^(a[16] & b[165])^(a[15] & b[166])^(a[14] & b[167])^(a[13] & b[168])^(a[12] & b[169])^(a[11] & b[170])^(a[10] & b[171])^(a[9] & b[172])^(a[8] & b[173])^(a[7] & b[174])^(a[6] & b[175])^(a[5] & b[176])^(a[4] & b[177])^(a[3] & b[178])^(a[2] & b[179])^(a[1] & b[180])^(a[0] & b[181]);
assign y[182] = (a[182] & b[0])^(a[181] & b[1])^(a[180] & b[2])^(a[179] & b[3])^(a[178] & b[4])^(a[177] & b[5])^(a[176] & b[6])^(a[175] & b[7])^(a[174] & b[8])^(a[173] & b[9])^(a[172] & b[10])^(a[171] & b[11])^(a[170] & b[12])^(a[169] & b[13])^(a[168] & b[14])^(a[167] & b[15])^(a[166] & b[16])^(a[165] & b[17])^(a[164] & b[18])^(a[163] & b[19])^(a[162] & b[20])^(a[161] & b[21])^(a[160] & b[22])^(a[159] & b[23])^(a[158] & b[24])^(a[157] & b[25])^(a[156] & b[26])^(a[155] & b[27])^(a[154] & b[28])^(a[153] & b[29])^(a[152] & b[30])^(a[151] & b[31])^(a[150] & b[32])^(a[149] & b[33])^(a[148] & b[34])^(a[147] & b[35])^(a[146] & b[36])^(a[145] & b[37])^(a[144] & b[38])^(a[143] & b[39])^(a[142] & b[40])^(a[141] & b[41])^(a[140] & b[42])^(a[139] & b[43])^(a[138] & b[44])^(a[137] & b[45])^(a[136] & b[46])^(a[135] & b[47])^(a[134] & b[48])^(a[133] & b[49])^(a[132] & b[50])^(a[131] & b[51])^(a[130] & b[52])^(a[129] & b[53])^(a[128] & b[54])^(a[127] & b[55])^(a[126] & b[56])^(a[125] & b[57])^(a[124] & b[58])^(a[123] & b[59])^(a[122] & b[60])^(a[121] & b[61])^(a[120] & b[62])^(a[119] & b[63])^(a[118] & b[64])^(a[117] & b[65])^(a[116] & b[66])^(a[115] & b[67])^(a[114] & b[68])^(a[113] & b[69])^(a[112] & b[70])^(a[111] & b[71])^(a[110] & b[72])^(a[109] & b[73])^(a[108] & b[74])^(a[107] & b[75])^(a[106] & b[76])^(a[105] & b[77])^(a[104] & b[78])^(a[103] & b[79])^(a[102] & b[80])^(a[101] & b[81])^(a[100] & b[82])^(a[99] & b[83])^(a[98] & b[84])^(a[97] & b[85])^(a[96] & b[86])^(a[95] & b[87])^(a[94] & b[88])^(a[93] & b[89])^(a[92] & b[90])^(a[91] & b[91])^(a[90] & b[92])^(a[89] & b[93])^(a[88] & b[94])^(a[87] & b[95])^(a[86] & b[96])^(a[85] & b[97])^(a[84] & b[98])^(a[83] & b[99])^(a[82] & b[100])^(a[81] & b[101])^(a[80] & b[102])^(a[79] & b[103])^(a[78] & b[104])^(a[77] & b[105])^(a[76] & b[106])^(a[75] & b[107])^(a[74] & b[108])^(a[73] & b[109])^(a[72] & b[110])^(a[71] & b[111])^(a[70] & b[112])^(a[69] & b[113])^(a[68] & b[114])^(a[67] & b[115])^(a[66] & b[116])^(a[65] & b[117])^(a[64] & b[118])^(a[63] & b[119])^(a[62] & b[120])^(a[61] & b[121])^(a[60] & b[122])^(a[59] & b[123])^(a[58] & b[124])^(a[57] & b[125])^(a[56] & b[126])^(a[55] & b[127])^(a[54] & b[128])^(a[53] & b[129])^(a[52] & b[130])^(a[51] & b[131])^(a[50] & b[132])^(a[49] & b[133])^(a[48] & b[134])^(a[47] & b[135])^(a[46] & b[136])^(a[45] & b[137])^(a[44] & b[138])^(a[43] & b[139])^(a[42] & b[140])^(a[41] & b[141])^(a[40] & b[142])^(a[39] & b[143])^(a[38] & b[144])^(a[37] & b[145])^(a[36] & b[146])^(a[35] & b[147])^(a[34] & b[148])^(a[33] & b[149])^(a[32] & b[150])^(a[31] & b[151])^(a[30] & b[152])^(a[29] & b[153])^(a[28] & b[154])^(a[27] & b[155])^(a[26] & b[156])^(a[25] & b[157])^(a[24] & b[158])^(a[23] & b[159])^(a[22] & b[160])^(a[21] & b[161])^(a[20] & b[162])^(a[19] & b[163])^(a[18] & b[164])^(a[17] & b[165])^(a[16] & b[166])^(a[15] & b[167])^(a[14] & b[168])^(a[13] & b[169])^(a[12] & b[170])^(a[11] & b[171])^(a[10] & b[172])^(a[9] & b[173])^(a[8] & b[174])^(a[7] & b[175])^(a[6] & b[176])^(a[5] & b[177])^(a[4] & b[178])^(a[3] & b[179])^(a[2] & b[180])^(a[1] & b[181])^(a[0] & b[182]);
assign y[183] = (a[183] & b[0])^(a[182] & b[1])^(a[181] & b[2])^(a[180] & b[3])^(a[179] & b[4])^(a[178] & b[5])^(a[177] & b[6])^(a[176] & b[7])^(a[175] & b[8])^(a[174] & b[9])^(a[173] & b[10])^(a[172] & b[11])^(a[171] & b[12])^(a[170] & b[13])^(a[169] & b[14])^(a[168] & b[15])^(a[167] & b[16])^(a[166] & b[17])^(a[165] & b[18])^(a[164] & b[19])^(a[163] & b[20])^(a[162] & b[21])^(a[161] & b[22])^(a[160] & b[23])^(a[159] & b[24])^(a[158] & b[25])^(a[157] & b[26])^(a[156] & b[27])^(a[155] & b[28])^(a[154] & b[29])^(a[153] & b[30])^(a[152] & b[31])^(a[151] & b[32])^(a[150] & b[33])^(a[149] & b[34])^(a[148] & b[35])^(a[147] & b[36])^(a[146] & b[37])^(a[145] & b[38])^(a[144] & b[39])^(a[143] & b[40])^(a[142] & b[41])^(a[141] & b[42])^(a[140] & b[43])^(a[139] & b[44])^(a[138] & b[45])^(a[137] & b[46])^(a[136] & b[47])^(a[135] & b[48])^(a[134] & b[49])^(a[133] & b[50])^(a[132] & b[51])^(a[131] & b[52])^(a[130] & b[53])^(a[129] & b[54])^(a[128] & b[55])^(a[127] & b[56])^(a[126] & b[57])^(a[125] & b[58])^(a[124] & b[59])^(a[123] & b[60])^(a[122] & b[61])^(a[121] & b[62])^(a[120] & b[63])^(a[119] & b[64])^(a[118] & b[65])^(a[117] & b[66])^(a[116] & b[67])^(a[115] & b[68])^(a[114] & b[69])^(a[113] & b[70])^(a[112] & b[71])^(a[111] & b[72])^(a[110] & b[73])^(a[109] & b[74])^(a[108] & b[75])^(a[107] & b[76])^(a[106] & b[77])^(a[105] & b[78])^(a[104] & b[79])^(a[103] & b[80])^(a[102] & b[81])^(a[101] & b[82])^(a[100] & b[83])^(a[99] & b[84])^(a[98] & b[85])^(a[97] & b[86])^(a[96] & b[87])^(a[95] & b[88])^(a[94] & b[89])^(a[93] & b[90])^(a[92] & b[91])^(a[91] & b[92])^(a[90] & b[93])^(a[89] & b[94])^(a[88] & b[95])^(a[87] & b[96])^(a[86] & b[97])^(a[85] & b[98])^(a[84] & b[99])^(a[83] & b[100])^(a[82] & b[101])^(a[81] & b[102])^(a[80] & b[103])^(a[79] & b[104])^(a[78] & b[105])^(a[77] & b[106])^(a[76] & b[107])^(a[75] & b[108])^(a[74] & b[109])^(a[73] & b[110])^(a[72] & b[111])^(a[71] & b[112])^(a[70] & b[113])^(a[69] & b[114])^(a[68] & b[115])^(a[67] & b[116])^(a[66] & b[117])^(a[65] & b[118])^(a[64] & b[119])^(a[63] & b[120])^(a[62] & b[121])^(a[61] & b[122])^(a[60] & b[123])^(a[59] & b[124])^(a[58] & b[125])^(a[57] & b[126])^(a[56] & b[127])^(a[55] & b[128])^(a[54] & b[129])^(a[53] & b[130])^(a[52] & b[131])^(a[51] & b[132])^(a[50] & b[133])^(a[49] & b[134])^(a[48] & b[135])^(a[47] & b[136])^(a[46] & b[137])^(a[45] & b[138])^(a[44] & b[139])^(a[43] & b[140])^(a[42] & b[141])^(a[41] & b[142])^(a[40] & b[143])^(a[39] & b[144])^(a[38] & b[145])^(a[37] & b[146])^(a[36] & b[147])^(a[35] & b[148])^(a[34] & b[149])^(a[33] & b[150])^(a[32] & b[151])^(a[31] & b[152])^(a[30] & b[153])^(a[29] & b[154])^(a[28] & b[155])^(a[27] & b[156])^(a[26] & b[157])^(a[25] & b[158])^(a[24] & b[159])^(a[23] & b[160])^(a[22] & b[161])^(a[21] & b[162])^(a[20] & b[163])^(a[19] & b[164])^(a[18] & b[165])^(a[17] & b[166])^(a[16] & b[167])^(a[15] & b[168])^(a[14] & b[169])^(a[13] & b[170])^(a[12] & b[171])^(a[11] & b[172])^(a[10] & b[173])^(a[9] & b[174])^(a[8] & b[175])^(a[7] & b[176])^(a[6] & b[177])^(a[5] & b[178])^(a[4] & b[179])^(a[3] & b[180])^(a[2] & b[181])^(a[1] & b[182])^(a[0] & b[183]);
assign y[184] = (a[184] & b[0])^(a[183] & b[1])^(a[182] & b[2])^(a[181] & b[3])^(a[180] & b[4])^(a[179] & b[5])^(a[178] & b[6])^(a[177] & b[7])^(a[176] & b[8])^(a[175] & b[9])^(a[174] & b[10])^(a[173] & b[11])^(a[172] & b[12])^(a[171] & b[13])^(a[170] & b[14])^(a[169] & b[15])^(a[168] & b[16])^(a[167] & b[17])^(a[166] & b[18])^(a[165] & b[19])^(a[164] & b[20])^(a[163] & b[21])^(a[162] & b[22])^(a[161] & b[23])^(a[160] & b[24])^(a[159] & b[25])^(a[158] & b[26])^(a[157] & b[27])^(a[156] & b[28])^(a[155] & b[29])^(a[154] & b[30])^(a[153] & b[31])^(a[152] & b[32])^(a[151] & b[33])^(a[150] & b[34])^(a[149] & b[35])^(a[148] & b[36])^(a[147] & b[37])^(a[146] & b[38])^(a[145] & b[39])^(a[144] & b[40])^(a[143] & b[41])^(a[142] & b[42])^(a[141] & b[43])^(a[140] & b[44])^(a[139] & b[45])^(a[138] & b[46])^(a[137] & b[47])^(a[136] & b[48])^(a[135] & b[49])^(a[134] & b[50])^(a[133] & b[51])^(a[132] & b[52])^(a[131] & b[53])^(a[130] & b[54])^(a[129] & b[55])^(a[128] & b[56])^(a[127] & b[57])^(a[126] & b[58])^(a[125] & b[59])^(a[124] & b[60])^(a[123] & b[61])^(a[122] & b[62])^(a[121] & b[63])^(a[120] & b[64])^(a[119] & b[65])^(a[118] & b[66])^(a[117] & b[67])^(a[116] & b[68])^(a[115] & b[69])^(a[114] & b[70])^(a[113] & b[71])^(a[112] & b[72])^(a[111] & b[73])^(a[110] & b[74])^(a[109] & b[75])^(a[108] & b[76])^(a[107] & b[77])^(a[106] & b[78])^(a[105] & b[79])^(a[104] & b[80])^(a[103] & b[81])^(a[102] & b[82])^(a[101] & b[83])^(a[100] & b[84])^(a[99] & b[85])^(a[98] & b[86])^(a[97] & b[87])^(a[96] & b[88])^(a[95] & b[89])^(a[94] & b[90])^(a[93] & b[91])^(a[92] & b[92])^(a[91] & b[93])^(a[90] & b[94])^(a[89] & b[95])^(a[88] & b[96])^(a[87] & b[97])^(a[86] & b[98])^(a[85] & b[99])^(a[84] & b[100])^(a[83] & b[101])^(a[82] & b[102])^(a[81] & b[103])^(a[80] & b[104])^(a[79] & b[105])^(a[78] & b[106])^(a[77] & b[107])^(a[76] & b[108])^(a[75] & b[109])^(a[74] & b[110])^(a[73] & b[111])^(a[72] & b[112])^(a[71] & b[113])^(a[70] & b[114])^(a[69] & b[115])^(a[68] & b[116])^(a[67] & b[117])^(a[66] & b[118])^(a[65] & b[119])^(a[64] & b[120])^(a[63] & b[121])^(a[62] & b[122])^(a[61] & b[123])^(a[60] & b[124])^(a[59] & b[125])^(a[58] & b[126])^(a[57] & b[127])^(a[56] & b[128])^(a[55] & b[129])^(a[54] & b[130])^(a[53] & b[131])^(a[52] & b[132])^(a[51] & b[133])^(a[50] & b[134])^(a[49] & b[135])^(a[48] & b[136])^(a[47] & b[137])^(a[46] & b[138])^(a[45] & b[139])^(a[44] & b[140])^(a[43] & b[141])^(a[42] & b[142])^(a[41] & b[143])^(a[40] & b[144])^(a[39] & b[145])^(a[38] & b[146])^(a[37] & b[147])^(a[36] & b[148])^(a[35] & b[149])^(a[34] & b[150])^(a[33] & b[151])^(a[32] & b[152])^(a[31] & b[153])^(a[30] & b[154])^(a[29] & b[155])^(a[28] & b[156])^(a[27] & b[157])^(a[26] & b[158])^(a[25] & b[159])^(a[24] & b[160])^(a[23] & b[161])^(a[22] & b[162])^(a[21] & b[163])^(a[20] & b[164])^(a[19] & b[165])^(a[18] & b[166])^(a[17] & b[167])^(a[16] & b[168])^(a[15] & b[169])^(a[14] & b[170])^(a[13] & b[171])^(a[12] & b[172])^(a[11] & b[173])^(a[10] & b[174])^(a[9] & b[175])^(a[8] & b[176])^(a[7] & b[177])^(a[6] & b[178])^(a[5] & b[179])^(a[4] & b[180])^(a[3] & b[181])^(a[2] & b[182])^(a[1] & b[183])^(a[0] & b[184]);
assign y[185] = (a[185] & b[0])^(a[184] & b[1])^(a[183] & b[2])^(a[182] & b[3])^(a[181] & b[4])^(a[180] & b[5])^(a[179] & b[6])^(a[178] & b[7])^(a[177] & b[8])^(a[176] & b[9])^(a[175] & b[10])^(a[174] & b[11])^(a[173] & b[12])^(a[172] & b[13])^(a[171] & b[14])^(a[170] & b[15])^(a[169] & b[16])^(a[168] & b[17])^(a[167] & b[18])^(a[166] & b[19])^(a[165] & b[20])^(a[164] & b[21])^(a[163] & b[22])^(a[162] & b[23])^(a[161] & b[24])^(a[160] & b[25])^(a[159] & b[26])^(a[158] & b[27])^(a[157] & b[28])^(a[156] & b[29])^(a[155] & b[30])^(a[154] & b[31])^(a[153] & b[32])^(a[152] & b[33])^(a[151] & b[34])^(a[150] & b[35])^(a[149] & b[36])^(a[148] & b[37])^(a[147] & b[38])^(a[146] & b[39])^(a[145] & b[40])^(a[144] & b[41])^(a[143] & b[42])^(a[142] & b[43])^(a[141] & b[44])^(a[140] & b[45])^(a[139] & b[46])^(a[138] & b[47])^(a[137] & b[48])^(a[136] & b[49])^(a[135] & b[50])^(a[134] & b[51])^(a[133] & b[52])^(a[132] & b[53])^(a[131] & b[54])^(a[130] & b[55])^(a[129] & b[56])^(a[128] & b[57])^(a[127] & b[58])^(a[126] & b[59])^(a[125] & b[60])^(a[124] & b[61])^(a[123] & b[62])^(a[122] & b[63])^(a[121] & b[64])^(a[120] & b[65])^(a[119] & b[66])^(a[118] & b[67])^(a[117] & b[68])^(a[116] & b[69])^(a[115] & b[70])^(a[114] & b[71])^(a[113] & b[72])^(a[112] & b[73])^(a[111] & b[74])^(a[110] & b[75])^(a[109] & b[76])^(a[108] & b[77])^(a[107] & b[78])^(a[106] & b[79])^(a[105] & b[80])^(a[104] & b[81])^(a[103] & b[82])^(a[102] & b[83])^(a[101] & b[84])^(a[100] & b[85])^(a[99] & b[86])^(a[98] & b[87])^(a[97] & b[88])^(a[96] & b[89])^(a[95] & b[90])^(a[94] & b[91])^(a[93] & b[92])^(a[92] & b[93])^(a[91] & b[94])^(a[90] & b[95])^(a[89] & b[96])^(a[88] & b[97])^(a[87] & b[98])^(a[86] & b[99])^(a[85] & b[100])^(a[84] & b[101])^(a[83] & b[102])^(a[82] & b[103])^(a[81] & b[104])^(a[80] & b[105])^(a[79] & b[106])^(a[78] & b[107])^(a[77] & b[108])^(a[76] & b[109])^(a[75] & b[110])^(a[74] & b[111])^(a[73] & b[112])^(a[72] & b[113])^(a[71] & b[114])^(a[70] & b[115])^(a[69] & b[116])^(a[68] & b[117])^(a[67] & b[118])^(a[66] & b[119])^(a[65] & b[120])^(a[64] & b[121])^(a[63] & b[122])^(a[62] & b[123])^(a[61] & b[124])^(a[60] & b[125])^(a[59] & b[126])^(a[58] & b[127])^(a[57] & b[128])^(a[56] & b[129])^(a[55] & b[130])^(a[54] & b[131])^(a[53] & b[132])^(a[52] & b[133])^(a[51] & b[134])^(a[50] & b[135])^(a[49] & b[136])^(a[48] & b[137])^(a[47] & b[138])^(a[46] & b[139])^(a[45] & b[140])^(a[44] & b[141])^(a[43] & b[142])^(a[42] & b[143])^(a[41] & b[144])^(a[40] & b[145])^(a[39] & b[146])^(a[38] & b[147])^(a[37] & b[148])^(a[36] & b[149])^(a[35] & b[150])^(a[34] & b[151])^(a[33] & b[152])^(a[32] & b[153])^(a[31] & b[154])^(a[30] & b[155])^(a[29] & b[156])^(a[28] & b[157])^(a[27] & b[158])^(a[26] & b[159])^(a[25] & b[160])^(a[24] & b[161])^(a[23] & b[162])^(a[22] & b[163])^(a[21] & b[164])^(a[20] & b[165])^(a[19] & b[166])^(a[18] & b[167])^(a[17] & b[168])^(a[16] & b[169])^(a[15] & b[170])^(a[14] & b[171])^(a[13] & b[172])^(a[12] & b[173])^(a[11] & b[174])^(a[10] & b[175])^(a[9] & b[176])^(a[8] & b[177])^(a[7] & b[178])^(a[6] & b[179])^(a[5] & b[180])^(a[4] & b[181])^(a[3] & b[182])^(a[2] & b[183])^(a[1] & b[184])^(a[0] & b[185]);
assign y[186] = (a[186] & b[0])^(a[185] & b[1])^(a[184] & b[2])^(a[183] & b[3])^(a[182] & b[4])^(a[181] & b[5])^(a[180] & b[6])^(a[179] & b[7])^(a[178] & b[8])^(a[177] & b[9])^(a[176] & b[10])^(a[175] & b[11])^(a[174] & b[12])^(a[173] & b[13])^(a[172] & b[14])^(a[171] & b[15])^(a[170] & b[16])^(a[169] & b[17])^(a[168] & b[18])^(a[167] & b[19])^(a[166] & b[20])^(a[165] & b[21])^(a[164] & b[22])^(a[163] & b[23])^(a[162] & b[24])^(a[161] & b[25])^(a[160] & b[26])^(a[159] & b[27])^(a[158] & b[28])^(a[157] & b[29])^(a[156] & b[30])^(a[155] & b[31])^(a[154] & b[32])^(a[153] & b[33])^(a[152] & b[34])^(a[151] & b[35])^(a[150] & b[36])^(a[149] & b[37])^(a[148] & b[38])^(a[147] & b[39])^(a[146] & b[40])^(a[145] & b[41])^(a[144] & b[42])^(a[143] & b[43])^(a[142] & b[44])^(a[141] & b[45])^(a[140] & b[46])^(a[139] & b[47])^(a[138] & b[48])^(a[137] & b[49])^(a[136] & b[50])^(a[135] & b[51])^(a[134] & b[52])^(a[133] & b[53])^(a[132] & b[54])^(a[131] & b[55])^(a[130] & b[56])^(a[129] & b[57])^(a[128] & b[58])^(a[127] & b[59])^(a[126] & b[60])^(a[125] & b[61])^(a[124] & b[62])^(a[123] & b[63])^(a[122] & b[64])^(a[121] & b[65])^(a[120] & b[66])^(a[119] & b[67])^(a[118] & b[68])^(a[117] & b[69])^(a[116] & b[70])^(a[115] & b[71])^(a[114] & b[72])^(a[113] & b[73])^(a[112] & b[74])^(a[111] & b[75])^(a[110] & b[76])^(a[109] & b[77])^(a[108] & b[78])^(a[107] & b[79])^(a[106] & b[80])^(a[105] & b[81])^(a[104] & b[82])^(a[103] & b[83])^(a[102] & b[84])^(a[101] & b[85])^(a[100] & b[86])^(a[99] & b[87])^(a[98] & b[88])^(a[97] & b[89])^(a[96] & b[90])^(a[95] & b[91])^(a[94] & b[92])^(a[93] & b[93])^(a[92] & b[94])^(a[91] & b[95])^(a[90] & b[96])^(a[89] & b[97])^(a[88] & b[98])^(a[87] & b[99])^(a[86] & b[100])^(a[85] & b[101])^(a[84] & b[102])^(a[83] & b[103])^(a[82] & b[104])^(a[81] & b[105])^(a[80] & b[106])^(a[79] & b[107])^(a[78] & b[108])^(a[77] & b[109])^(a[76] & b[110])^(a[75] & b[111])^(a[74] & b[112])^(a[73] & b[113])^(a[72] & b[114])^(a[71] & b[115])^(a[70] & b[116])^(a[69] & b[117])^(a[68] & b[118])^(a[67] & b[119])^(a[66] & b[120])^(a[65] & b[121])^(a[64] & b[122])^(a[63] & b[123])^(a[62] & b[124])^(a[61] & b[125])^(a[60] & b[126])^(a[59] & b[127])^(a[58] & b[128])^(a[57] & b[129])^(a[56] & b[130])^(a[55] & b[131])^(a[54] & b[132])^(a[53] & b[133])^(a[52] & b[134])^(a[51] & b[135])^(a[50] & b[136])^(a[49] & b[137])^(a[48] & b[138])^(a[47] & b[139])^(a[46] & b[140])^(a[45] & b[141])^(a[44] & b[142])^(a[43] & b[143])^(a[42] & b[144])^(a[41] & b[145])^(a[40] & b[146])^(a[39] & b[147])^(a[38] & b[148])^(a[37] & b[149])^(a[36] & b[150])^(a[35] & b[151])^(a[34] & b[152])^(a[33] & b[153])^(a[32] & b[154])^(a[31] & b[155])^(a[30] & b[156])^(a[29] & b[157])^(a[28] & b[158])^(a[27] & b[159])^(a[26] & b[160])^(a[25] & b[161])^(a[24] & b[162])^(a[23] & b[163])^(a[22] & b[164])^(a[21] & b[165])^(a[20] & b[166])^(a[19] & b[167])^(a[18] & b[168])^(a[17] & b[169])^(a[16] & b[170])^(a[15] & b[171])^(a[14] & b[172])^(a[13] & b[173])^(a[12] & b[174])^(a[11] & b[175])^(a[10] & b[176])^(a[9] & b[177])^(a[8] & b[178])^(a[7] & b[179])^(a[6] & b[180])^(a[5] & b[181])^(a[4] & b[182])^(a[3] & b[183])^(a[2] & b[184])^(a[1] & b[185])^(a[0] & b[186]);
assign y[187] = (a[187] & b[0])^(a[186] & b[1])^(a[185] & b[2])^(a[184] & b[3])^(a[183] & b[4])^(a[182] & b[5])^(a[181] & b[6])^(a[180] & b[7])^(a[179] & b[8])^(a[178] & b[9])^(a[177] & b[10])^(a[176] & b[11])^(a[175] & b[12])^(a[174] & b[13])^(a[173] & b[14])^(a[172] & b[15])^(a[171] & b[16])^(a[170] & b[17])^(a[169] & b[18])^(a[168] & b[19])^(a[167] & b[20])^(a[166] & b[21])^(a[165] & b[22])^(a[164] & b[23])^(a[163] & b[24])^(a[162] & b[25])^(a[161] & b[26])^(a[160] & b[27])^(a[159] & b[28])^(a[158] & b[29])^(a[157] & b[30])^(a[156] & b[31])^(a[155] & b[32])^(a[154] & b[33])^(a[153] & b[34])^(a[152] & b[35])^(a[151] & b[36])^(a[150] & b[37])^(a[149] & b[38])^(a[148] & b[39])^(a[147] & b[40])^(a[146] & b[41])^(a[145] & b[42])^(a[144] & b[43])^(a[143] & b[44])^(a[142] & b[45])^(a[141] & b[46])^(a[140] & b[47])^(a[139] & b[48])^(a[138] & b[49])^(a[137] & b[50])^(a[136] & b[51])^(a[135] & b[52])^(a[134] & b[53])^(a[133] & b[54])^(a[132] & b[55])^(a[131] & b[56])^(a[130] & b[57])^(a[129] & b[58])^(a[128] & b[59])^(a[127] & b[60])^(a[126] & b[61])^(a[125] & b[62])^(a[124] & b[63])^(a[123] & b[64])^(a[122] & b[65])^(a[121] & b[66])^(a[120] & b[67])^(a[119] & b[68])^(a[118] & b[69])^(a[117] & b[70])^(a[116] & b[71])^(a[115] & b[72])^(a[114] & b[73])^(a[113] & b[74])^(a[112] & b[75])^(a[111] & b[76])^(a[110] & b[77])^(a[109] & b[78])^(a[108] & b[79])^(a[107] & b[80])^(a[106] & b[81])^(a[105] & b[82])^(a[104] & b[83])^(a[103] & b[84])^(a[102] & b[85])^(a[101] & b[86])^(a[100] & b[87])^(a[99] & b[88])^(a[98] & b[89])^(a[97] & b[90])^(a[96] & b[91])^(a[95] & b[92])^(a[94] & b[93])^(a[93] & b[94])^(a[92] & b[95])^(a[91] & b[96])^(a[90] & b[97])^(a[89] & b[98])^(a[88] & b[99])^(a[87] & b[100])^(a[86] & b[101])^(a[85] & b[102])^(a[84] & b[103])^(a[83] & b[104])^(a[82] & b[105])^(a[81] & b[106])^(a[80] & b[107])^(a[79] & b[108])^(a[78] & b[109])^(a[77] & b[110])^(a[76] & b[111])^(a[75] & b[112])^(a[74] & b[113])^(a[73] & b[114])^(a[72] & b[115])^(a[71] & b[116])^(a[70] & b[117])^(a[69] & b[118])^(a[68] & b[119])^(a[67] & b[120])^(a[66] & b[121])^(a[65] & b[122])^(a[64] & b[123])^(a[63] & b[124])^(a[62] & b[125])^(a[61] & b[126])^(a[60] & b[127])^(a[59] & b[128])^(a[58] & b[129])^(a[57] & b[130])^(a[56] & b[131])^(a[55] & b[132])^(a[54] & b[133])^(a[53] & b[134])^(a[52] & b[135])^(a[51] & b[136])^(a[50] & b[137])^(a[49] & b[138])^(a[48] & b[139])^(a[47] & b[140])^(a[46] & b[141])^(a[45] & b[142])^(a[44] & b[143])^(a[43] & b[144])^(a[42] & b[145])^(a[41] & b[146])^(a[40] & b[147])^(a[39] & b[148])^(a[38] & b[149])^(a[37] & b[150])^(a[36] & b[151])^(a[35] & b[152])^(a[34] & b[153])^(a[33] & b[154])^(a[32] & b[155])^(a[31] & b[156])^(a[30] & b[157])^(a[29] & b[158])^(a[28] & b[159])^(a[27] & b[160])^(a[26] & b[161])^(a[25] & b[162])^(a[24] & b[163])^(a[23] & b[164])^(a[22] & b[165])^(a[21] & b[166])^(a[20] & b[167])^(a[19] & b[168])^(a[18] & b[169])^(a[17] & b[170])^(a[16] & b[171])^(a[15] & b[172])^(a[14] & b[173])^(a[13] & b[174])^(a[12] & b[175])^(a[11] & b[176])^(a[10] & b[177])^(a[9] & b[178])^(a[8] & b[179])^(a[7] & b[180])^(a[6] & b[181])^(a[5] & b[182])^(a[4] & b[183])^(a[3] & b[184])^(a[2] & b[185])^(a[1] & b[186])^(a[0] & b[187]);
assign y[188] = (a[188] & b[0])^(a[187] & b[1])^(a[186] & b[2])^(a[185] & b[3])^(a[184] & b[4])^(a[183] & b[5])^(a[182] & b[6])^(a[181] & b[7])^(a[180] & b[8])^(a[179] & b[9])^(a[178] & b[10])^(a[177] & b[11])^(a[176] & b[12])^(a[175] & b[13])^(a[174] & b[14])^(a[173] & b[15])^(a[172] & b[16])^(a[171] & b[17])^(a[170] & b[18])^(a[169] & b[19])^(a[168] & b[20])^(a[167] & b[21])^(a[166] & b[22])^(a[165] & b[23])^(a[164] & b[24])^(a[163] & b[25])^(a[162] & b[26])^(a[161] & b[27])^(a[160] & b[28])^(a[159] & b[29])^(a[158] & b[30])^(a[157] & b[31])^(a[156] & b[32])^(a[155] & b[33])^(a[154] & b[34])^(a[153] & b[35])^(a[152] & b[36])^(a[151] & b[37])^(a[150] & b[38])^(a[149] & b[39])^(a[148] & b[40])^(a[147] & b[41])^(a[146] & b[42])^(a[145] & b[43])^(a[144] & b[44])^(a[143] & b[45])^(a[142] & b[46])^(a[141] & b[47])^(a[140] & b[48])^(a[139] & b[49])^(a[138] & b[50])^(a[137] & b[51])^(a[136] & b[52])^(a[135] & b[53])^(a[134] & b[54])^(a[133] & b[55])^(a[132] & b[56])^(a[131] & b[57])^(a[130] & b[58])^(a[129] & b[59])^(a[128] & b[60])^(a[127] & b[61])^(a[126] & b[62])^(a[125] & b[63])^(a[124] & b[64])^(a[123] & b[65])^(a[122] & b[66])^(a[121] & b[67])^(a[120] & b[68])^(a[119] & b[69])^(a[118] & b[70])^(a[117] & b[71])^(a[116] & b[72])^(a[115] & b[73])^(a[114] & b[74])^(a[113] & b[75])^(a[112] & b[76])^(a[111] & b[77])^(a[110] & b[78])^(a[109] & b[79])^(a[108] & b[80])^(a[107] & b[81])^(a[106] & b[82])^(a[105] & b[83])^(a[104] & b[84])^(a[103] & b[85])^(a[102] & b[86])^(a[101] & b[87])^(a[100] & b[88])^(a[99] & b[89])^(a[98] & b[90])^(a[97] & b[91])^(a[96] & b[92])^(a[95] & b[93])^(a[94] & b[94])^(a[93] & b[95])^(a[92] & b[96])^(a[91] & b[97])^(a[90] & b[98])^(a[89] & b[99])^(a[88] & b[100])^(a[87] & b[101])^(a[86] & b[102])^(a[85] & b[103])^(a[84] & b[104])^(a[83] & b[105])^(a[82] & b[106])^(a[81] & b[107])^(a[80] & b[108])^(a[79] & b[109])^(a[78] & b[110])^(a[77] & b[111])^(a[76] & b[112])^(a[75] & b[113])^(a[74] & b[114])^(a[73] & b[115])^(a[72] & b[116])^(a[71] & b[117])^(a[70] & b[118])^(a[69] & b[119])^(a[68] & b[120])^(a[67] & b[121])^(a[66] & b[122])^(a[65] & b[123])^(a[64] & b[124])^(a[63] & b[125])^(a[62] & b[126])^(a[61] & b[127])^(a[60] & b[128])^(a[59] & b[129])^(a[58] & b[130])^(a[57] & b[131])^(a[56] & b[132])^(a[55] & b[133])^(a[54] & b[134])^(a[53] & b[135])^(a[52] & b[136])^(a[51] & b[137])^(a[50] & b[138])^(a[49] & b[139])^(a[48] & b[140])^(a[47] & b[141])^(a[46] & b[142])^(a[45] & b[143])^(a[44] & b[144])^(a[43] & b[145])^(a[42] & b[146])^(a[41] & b[147])^(a[40] & b[148])^(a[39] & b[149])^(a[38] & b[150])^(a[37] & b[151])^(a[36] & b[152])^(a[35] & b[153])^(a[34] & b[154])^(a[33] & b[155])^(a[32] & b[156])^(a[31] & b[157])^(a[30] & b[158])^(a[29] & b[159])^(a[28] & b[160])^(a[27] & b[161])^(a[26] & b[162])^(a[25] & b[163])^(a[24] & b[164])^(a[23] & b[165])^(a[22] & b[166])^(a[21] & b[167])^(a[20] & b[168])^(a[19] & b[169])^(a[18] & b[170])^(a[17] & b[171])^(a[16] & b[172])^(a[15] & b[173])^(a[14] & b[174])^(a[13] & b[175])^(a[12] & b[176])^(a[11] & b[177])^(a[10] & b[178])^(a[9] & b[179])^(a[8] & b[180])^(a[7] & b[181])^(a[6] & b[182])^(a[5] & b[183])^(a[4] & b[184])^(a[3] & b[185])^(a[2] & b[186])^(a[1] & b[187])^(a[0] & b[188]);
assign y[189] = (a[189] & b[0])^(a[188] & b[1])^(a[187] & b[2])^(a[186] & b[3])^(a[185] & b[4])^(a[184] & b[5])^(a[183] & b[6])^(a[182] & b[7])^(a[181] & b[8])^(a[180] & b[9])^(a[179] & b[10])^(a[178] & b[11])^(a[177] & b[12])^(a[176] & b[13])^(a[175] & b[14])^(a[174] & b[15])^(a[173] & b[16])^(a[172] & b[17])^(a[171] & b[18])^(a[170] & b[19])^(a[169] & b[20])^(a[168] & b[21])^(a[167] & b[22])^(a[166] & b[23])^(a[165] & b[24])^(a[164] & b[25])^(a[163] & b[26])^(a[162] & b[27])^(a[161] & b[28])^(a[160] & b[29])^(a[159] & b[30])^(a[158] & b[31])^(a[157] & b[32])^(a[156] & b[33])^(a[155] & b[34])^(a[154] & b[35])^(a[153] & b[36])^(a[152] & b[37])^(a[151] & b[38])^(a[150] & b[39])^(a[149] & b[40])^(a[148] & b[41])^(a[147] & b[42])^(a[146] & b[43])^(a[145] & b[44])^(a[144] & b[45])^(a[143] & b[46])^(a[142] & b[47])^(a[141] & b[48])^(a[140] & b[49])^(a[139] & b[50])^(a[138] & b[51])^(a[137] & b[52])^(a[136] & b[53])^(a[135] & b[54])^(a[134] & b[55])^(a[133] & b[56])^(a[132] & b[57])^(a[131] & b[58])^(a[130] & b[59])^(a[129] & b[60])^(a[128] & b[61])^(a[127] & b[62])^(a[126] & b[63])^(a[125] & b[64])^(a[124] & b[65])^(a[123] & b[66])^(a[122] & b[67])^(a[121] & b[68])^(a[120] & b[69])^(a[119] & b[70])^(a[118] & b[71])^(a[117] & b[72])^(a[116] & b[73])^(a[115] & b[74])^(a[114] & b[75])^(a[113] & b[76])^(a[112] & b[77])^(a[111] & b[78])^(a[110] & b[79])^(a[109] & b[80])^(a[108] & b[81])^(a[107] & b[82])^(a[106] & b[83])^(a[105] & b[84])^(a[104] & b[85])^(a[103] & b[86])^(a[102] & b[87])^(a[101] & b[88])^(a[100] & b[89])^(a[99] & b[90])^(a[98] & b[91])^(a[97] & b[92])^(a[96] & b[93])^(a[95] & b[94])^(a[94] & b[95])^(a[93] & b[96])^(a[92] & b[97])^(a[91] & b[98])^(a[90] & b[99])^(a[89] & b[100])^(a[88] & b[101])^(a[87] & b[102])^(a[86] & b[103])^(a[85] & b[104])^(a[84] & b[105])^(a[83] & b[106])^(a[82] & b[107])^(a[81] & b[108])^(a[80] & b[109])^(a[79] & b[110])^(a[78] & b[111])^(a[77] & b[112])^(a[76] & b[113])^(a[75] & b[114])^(a[74] & b[115])^(a[73] & b[116])^(a[72] & b[117])^(a[71] & b[118])^(a[70] & b[119])^(a[69] & b[120])^(a[68] & b[121])^(a[67] & b[122])^(a[66] & b[123])^(a[65] & b[124])^(a[64] & b[125])^(a[63] & b[126])^(a[62] & b[127])^(a[61] & b[128])^(a[60] & b[129])^(a[59] & b[130])^(a[58] & b[131])^(a[57] & b[132])^(a[56] & b[133])^(a[55] & b[134])^(a[54] & b[135])^(a[53] & b[136])^(a[52] & b[137])^(a[51] & b[138])^(a[50] & b[139])^(a[49] & b[140])^(a[48] & b[141])^(a[47] & b[142])^(a[46] & b[143])^(a[45] & b[144])^(a[44] & b[145])^(a[43] & b[146])^(a[42] & b[147])^(a[41] & b[148])^(a[40] & b[149])^(a[39] & b[150])^(a[38] & b[151])^(a[37] & b[152])^(a[36] & b[153])^(a[35] & b[154])^(a[34] & b[155])^(a[33] & b[156])^(a[32] & b[157])^(a[31] & b[158])^(a[30] & b[159])^(a[29] & b[160])^(a[28] & b[161])^(a[27] & b[162])^(a[26] & b[163])^(a[25] & b[164])^(a[24] & b[165])^(a[23] & b[166])^(a[22] & b[167])^(a[21] & b[168])^(a[20] & b[169])^(a[19] & b[170])^(a[18] & b[171])^(a[17] & b[172])^(a[16] & b[173])^(a[15] & b[174])^(a[14] & b[175])^(a[13] & b[176])^(a[12] & b[177])^(a[11] & b[178])^(a[10] & b[179])^(a[9] & b[180])^(a[8] & b[181])^(a[7] & b[182])^(a[6] & b[183])^(a[5] & b[184])^(a[4] & b[185])^(a[3] & b[186])^(a[2] & b[187])^(a[1] & b[188])^(a[0] & b[189]);
assign y[190] = (a[190] & b[0])^(a[189] & b[1])^(a[188] & b[2])^(a[187] & b[3])^(a[186] & b[4])^(a[185] & b[5])^(a[184] & b[6])^(a[183] & b[7])^(a[182] & b[8])^(a[181] & b[9])^(a[180] & b[10])^(a[179] & b[11])^(a[178] & b[12])^(a[177] & b[13])^(a[176] & b[14])^(a[175] & b[15])^(a[174] & b[16])^(a[173] & b[17])^(a[172] & b[18])^(a[171] & b[19])^(a[170] & b[20])^(a[169] & b[21])^(a[168] & b[22])^(a[167] & b[23])^(a[166] & b[24])^(a[165] & b[25])^(a[164] & b[26])^(a[163] & b[27])^(a[162] & b[28])^(a[161] & b[29])^(a[160] & b[30])^(a[159] & b[31])^(a[158] & b[32])^(a[157] & b[33])^(a[156] & b[34])^(a[155] & b[35])^(a[154] & b[36])^(a[153] & b[37])^(a[152] & b[38])^(a[151] & b[39])^(a[150] & b[40])^(a[149] & b[41])^(a[148] & b[42])^(a[147] & b[43])^(a[146] & b[44])^(a[145] & b[45])^(a[144] & b[46])^(a[143] & b[47])^(a[142] & b[48])^(a[141] & b[49])^(a[140] & b[50])^(a[139] & b[51])^(a[138] & b[52])^(a[137] & b[53])^(a[136] & b[54])^(a[135] & b[55])^(a[134] & b[56])^(a[133] & b[57])^(a[132] & b[58])^(a[131] & b[59])^(a[130] & b[60])^(a[129] & b[61])^(a[128] & b[62])^(a[127] & b[63])^(a[126] & b[64])^(a[125] & b[65])^(a[124] & b[66])^(a[123] & b[67])^(a[122] & b[68])^(a[121] & b[69])^(a[120] & b[70])^(a[119] & b[71])^(a[118] & b[72])^(a[117] & b[73])^(a[116] & b[74])^(a[115] & b[75])^(a[114] & b[76])^(a[113] & b[77])^(a[112] & b[78])^(a[111] & b[79])^(a[110] & b[80])^(a[109] & b[81])^(a[108] & b[82])^(a[107] & b[83])^(a[106] & b[84])^(a[105] & b[85])^(a[104] & b[86])^(a[103] & b[87])^(a[102] & b[88])^(a[101] & b[89])^(a[100] & b[90])^(a[99] & b[91])^(a[98] & b[92])^(a[97] & b[93])^(a[96] & b[94])^(a[95] & b[95])^(a[94] & b[96])^(a[93] & b[97])^(a[92] & b[98])^(a[91] & b[99])^(a[90] & b[100])^(a[89] & b[101])^(a[88] & b[102])^(a[87] & b[103])^(a[86] & b[104])^(a[85] & b[105])^(a[84] & b[106])^(a[83] & b[107])^(a[82] & b[108])^(a[81] & b[109])^(a[80] & b[110])^(a[79] & b[111])^(a[78] & b[112])^(a[77] & b[113])^(a[76] & b[114])^(a[75] & b[115])^(a[74] & b[116])^(a[73] & b[117])^(a[72] & b[118])^(a[71] & b[119])^(a[70] & b[120])^(a[69] & b[121])^(a[68] & b[122])^(a[67] & b[123])^(a[66] & b[124])^(a[65] & b[125])^(a[64] & b[126])^(a[63] & b[127])^(a[62] & b[128])^(a[61] & b[129])^(a[60] & b[130])^(a[59] & b[131])^(a[58] & b[132])^(a[57] & b[133])^(a[56] & b[134])^(a[55] & b[135])^(a[54] & b[136])^(a[53] & b[137])^(a[52] & b[138])^(a[51] & b[139])^(a[50] & b[140])^(a[49] & b[141])^(a[48] & b[142])^(a[47] & b[143])^(a[46] & b[144])^(a[45] & b[145])^(a[44] & b[146])^(a[43] & b[147])^(a[42] & b[148])^(a[41] & b[149])^(a[40] & b[150])^(a[39] & b[151])^(a[38] & b[152])^(a[37] & b[153])^(a[36] & b[154])^(a[35] & b[155])^(a[34] & b[156])^(a[33] & b[157])^(a[32] & b[158])^(a[31] & b[159])^(a[30] & b[160])^(a[29] & b[161])^(a[28] & b[162])^(a[27] & b[163])^(a[26] & b[164])^(a[25] & b[165])^(a[24] & b[166])^(a[23] & b[167])^(a[22] & b[168])^(a[21] & b[169])^(a[20] & b[170])^(a[19] & b[171])^(a[18] & b[172])^(a[17] & b[173])^(a[16] & b[174])^(a[15] & b[175])^(a[14] & b[176])^(a[13] & b[177])^(a[12] & b[178])^(a[11] & b[179])^(a[10] & b[180])^(a[9] & b[181])^(a[8] & b[182])^(a[7] & b[183])^(a[6] & b[184])^(a[5] & b[185])^(a[4] & b[186])^(a[3] & b[187])^(a[2] & b[188])^(a[1] & b[189])^(a[0] & b[190]);
assign y[191] = (a[191] & b[0])^(a[190] & b[1])^(a[189] & b[2])^(a[188] & b[3])^(a[187] & b[4])^(a[186] & b[5])^(a[185] & b[6])^(a[184] & b[7])^(a[183] & b[8])^(a[182] & b[9])^(a[181] & b[10])^(a[180] & b[11])^(a[179] & b[12])^(a[178] & b[13])^(a[177] & b[14])^(a[176] & b[15])^(a[175] & b[16])^(a[174] & b[17])^(a[173] & b[18])^(a[172] & b[19])^(a[171] & b[20])^(a[170] & b[21])^(a[169] & b[22])^(a[168] & b[23])^(a[167] & b[24])^(a[166] & b[25])^(a[165] & b[26])^(a[164] & b[27])^(a[163] & b[28])^(a[162] & b[29])^(a[161] & b[30])^(a[160] & b[31])^(a[159] & b[32])^(a[158] & b[33])^(a[157] & b[34])^(a[156] & b[35])^(a[155] & b[36])^(a[154] & b[37])^(a[153] & b[38])^(a[152] & b[39])^(a[151] & b[40])^(a[150] & b[41])^(a[149] & b[42])^(a[148] & b[43])^(a[147] & b[44])^(a[146] & b[45])^(a[145] & b[46])^(a[144] & b[47])^(a[143] & b[48])^(a[142] & b[49])^(a[141] & b[50])^(a[140] & b[51])^(a[139] & b[52])^(a[138] & b[53])^(a[137] & b[54])^(a[136] & b[55])^(a[135] & b[56])^(a[134] & b[57])^(a[133] & b[58])^(a[132] & b[59])^(a[131] & b[60])^(a[130] & b[61])^(a[129] & b[62])^(a[128] & b[63])^(a[127] & b[64])^(a[126] & b[65])^(a[125] & b[66])^(a[124] & b[67])^(a[123] & b[68])^(a[122] & b[69])^(a[121] & b[70])^(a[120] & b[71])^(a[119] & b[72])^(a[118] & b[73])^(a[117] & b[74])^(a[116] & b[75])^(a[115] & b[76])^(a[114] & b[77])^(a[113] & b[78])^(a[112] & b[79])^(a[111] & b[80])^(a[110] & b[81])^(a[109] & b[82])^(a[108] & b[83])^(a[107] & b[84])^(a[106] & b[85])^(a[105] & b[86])^(a[104] & b[87])^(a[103] & b[88])^(a[102] & b[89])^(a[101] & b[90])^(a[100] & b[91])^(a[99] & b[92])^(a[98] & b[93])^(a[97] & b[94])^(a[96] & b[95])^(a[95] & b[96])^(a[94] & b[97])^(a[93] & b[98])^(a[92] & b[99])^(a[91] & b[100])^(a[90] & b[101])^(a[89] & b[102])^(a[88] & b[103])^(a[87] & b[104])^(a[86] & b[105])^(a[85] & b[106])^(a[84] & b[107])^(a[83] & b[108])^(a[82] & b[109])^(a[81] & b[110])^(a[80] & b[111])^(a[79] & b[112])^(a[78] & b[113])^(a[77] & b[114])^(a[76] & b[115])^(a[75] & b[116])^(a[74] & b[117])^(a[73] & b[118])^(a[72] & b[119])^(a[71] & b[120])^(a[70] & b[121])^(a[69] & b[122])^(a[68] & b[123])^(a[67] & b[124])^(a[66] & b[125])^(a[65] & b[126])^(a[64] & b[127])^(a[63] & b[128])^(a[62] & b[129])^(a[61] & b[130])^(a[60] & b[131])^(a[59] & b[132])^(a[58] & b[133])^(a[57] & b[134])^(a[56] & b[135])^(a[55] & b[136])^(a[54] & b[137])^(a[53] & b[138])^(a[52] & b[139])^(a[51] & b[140])^(a[50] & b[141])^(a[49] & b[142])^(a[48] & b[143])^(a[47] & b[144])^(a[46] & b[145])^(a[45] & b[146])^(a[44] & b[147])^(a[43] & b[148])^(a[42] & b[149])^(a[41] & b[150])^(a[40] & b[151])^(a[39] & b[152])^(a[38] & b[153])^(a[37] & b[154])^(a[36] & b[155])^(a[35] & b[156])^(a[34] & b[157])^(a[33] & b[158])^(a[32] & b[159])^(a[31] & b[160])^(a[30] & b[161])^(a[29] & b[162])^(a[28] & b[163])^(a[27] & b[164])^(a[26] & b[165])^(a[25] & b[166])^(a[24] & b[167])^(a[23] & b[168])^(a[22] & b[169])^(a[21] & b[170])^(a[20] & b[171])^(a[19] & b[172])^(a[18] & b[173])^(a[17] & b[174])^(a[16] & b[175])^(a[15] & b[176])^(a[14] & b[177])^(a[13] & b[178])^(a[12] & b[179])^(a[11] & b[180])^(a[10] & b[181])^(a[9] & b[182])^(a[8] & b[183])^(a[7] & b[184])^(a[6] & b[185])^(a[5] & b[186])^(a[4] & b[187])^(a[3] & b[188])^(a[2] & b[189])^(a[1] & b[190])^(a[0] & b[191]);
assign y[192] = (a[192] & b[0])^(a[191] & b[1])^(a[190] & b[2])^(a[189] & b[3])^(a[188] & b[4])^(a[187] & b[5])^(a[186] & b[6])^(a[185] & b[7])^(a[184] & b[8])^(a[183] & b[9])^(a[182] & b[10])^(a[181] & b[11])^(a[180] & b[12])^(a[179] & b[13])^(a[178] & b[14])^(a[177] & b[15])^(a[176] & b[16])^(a[175] & b[17])^(a[174] & b[18])^(a[173] & b[19])^(a[172] & b[20])^(a[171] & b[21])^(a[170] & b[22])^(a[169] & b[23])^(a[168] & b[24])^(a[167] & b[25])^(a[166] & b[26])^(a[165] & b[27])^(a[164] & b[28])^(a[163] & b[29])^(a[162] & b[30])^(a[161] & b[31])^(a[160] & b[32])^(a[159] & b[33])^(a[158] & b[34])^(a[157] & b[35])^(a[156] & b[36])^(a[155] & b[37])^(a[154] & b[38])^(a[153] & b[39])^(a[152] & b[40])^(a[151] & b[41])^(a[150] & b[42])^(a[149] & b[43])^(a[148] & b[44])^(a[147] & b[45])^(a[146] & b[46])^(a[145] & b[47])^(a[144] & b[48])^(a[143] & b[49])^(a[142] & b[50])^(a[141] & b[51])^(a[140] & b[52])^(a[139] & b[53])^(a[138] & b[54])^(a[137] & b[55])^(a[136] & b[56])^(a[135] & b[57])^(a[134] & b[58])^(a[133] & b[59])^(a[132] & b[60])^(a[131] & b[61])^(a[130] & b[62])^(a[129] & b[63])^(a[128] & b[64])^(a[127] & b[65])^(a[126] & b[66])^(a[125] & b[67])^(a[124] & b[68])^(a[123] & b[69])^(a[122] & b[70])^(a[121] & b[71])^(a[120] & b[72])^(a[119] & b[73])^(a[118] & b[74])^(a[117] & b[75])^(a[116] & b[76])^(a[115] & b[77])^(a[114] & b[78])^(a[113] & b[79])^(a[112] & b[80])^(a[111] & b[81])^(a[110] & b[82])^(a[109] & b[83])^(a[108] & b[84])^(a[107] & b[85])^(a[106] & b[86])^(a[105] & b[87])^(a[104] & b[88])^(a[103] & b[89])^(a[102] & b[90])^(a[101] & b[91])^(a[100] & b[92])^(a[99] & b[93])^(a[98] & b[94])^(a[97] & b[95])^(a[96] & b[96])^(a[95] & b[97])^(a[94] & b[98])^(a[93] & b[99])^(a[92] & b[100])^(a[91] & b[101])^(a[90] & b[102])^(a[89] & b[103])^(a[88] & b[104])^(a[87] & b[105])^(a[86] & b[106])^(a[85] & b[107])^(a[84] & b[108])^(a[83] & b[109])^(a[82] & b[110])^(a[81] & b[111])^(a[80] & b[112])^(a[79] & b[113])^(a[78] & b[114])^(a[77] & b[115])^(a[76] & b[116])^(a[75] & b[117])^(a[74] & b[118])^(a[73] & b[119])^(a[72] & b[120])^(a[71] & b[121])^(a[70] & b[122])^(a[69] & b[123])^(a[68] & b[124])^(a[67] & b[125])^(a[66] & b[126])^(a[65] & b[127])^(a[64] & b[128])^(a[63] & b[129])^(a[62] & b[130])^(a[61] & b[131])^(a[60] & b[132])^(a[59] & b[133])^(a[58] & b[134])^(a[57] & b[135])^(a[56] & b[136])^(a[55] & b[137])^(a[54] & b[138])^(a[53] & b[139])^(a[52] & b[140])^(a[51] & b[141])^(a[50] & b[142])^(a[49] & b[143])^(a[48] & b[144])^(a[47] & b[145])^(a[46] & b[146])^(a[45] & b[147])^(a[44] & b[148])^(a[43] & b[149])^(a[42] & b[150])^(a[41] & b[151])^(a[40] & b[152])^(a[39] & b[153])^(a[38] & b[154])^(a[37] & b[155])^(a[36] & b[156])^(a[35] & b[157])^(a[34] & b[158])^(a[33] & b[159])^(a[32] & b[160])^(a[31] & b[161])^(a[30] & b[162])^(a[29] & b[163])^(a[28] & b[164])^(a[27] & b[165])^(a[26] & b[166])^(a[25] & b[167])^(a[24] & b[168])^(a[23] & b[169])^(a[22] & b[170])^(a[21] & b[171])^(a[20] & b[172])^(a[19] & b[173])^(a[18] & b[174])^(a[17] & b[175])^(a[16] & b[176])^(a[15] & b[177])^(a[14] & b[178])^(a[13] & b[179])^(a[12] & b[180])^(a[11] & b[181])^(a[10] & b[182])^(a[9] & b[183])^(a[8] & b[184])^(a[7] & b[185])^(a[6] & b[186])^(a[5] & b[187])^(a[4] & b[188])^(a[3] & b[189])^(a[2] & b[190])^(a[1] & b[191])^(a[0] & b[192]);
assign y[193] = (a[193] & b[0])^(a[192] & b[1])^(a[191] & b[2])^(a[190] & b[3])^(a[189] & b[4])^(a[188] & b[5])^(a[187] & b[6])^(a[186] & b[7])^(a[185] & b[8])^(a[184] & b[9])^(a[183] & b[10])^(a[182] & b[11])^(a[181] & b[12])^(a[180] & b[13])^(a[179] & b[14])^(a[178] & b[15])^(a[177] & b[16])^(a[176] & b[17])^(a[175] & b[18])^(a[174] & b[19])^(a[173] & b[20])^(a[172] & b[21])^(a[171] & b[22])^(a[170] & b[23])^(a[169] & b[24])^(a[168] & b[25])^(a[167] & b[26])^(a[166] & b[27])^(a[165] & b[28])^(a[164] & b[29])^(a[163] & b[30])^(a[162] & b[31])^(a[161] & b[32])^(a[160] & b[33])^(a[159] & b[34])^(a[158] & b[35])^(a[157] & b[36])^(a[156] & b[37])^(a[155] & b[38])^(a[154] & b[39])^(a[153] & b[40])^(a[152] & b[41])^(a[151] & b[42])^(a[150] & b[43])^(a[149] & b[44])^(a[148] & b[45])^(a[147] & b[46])^(a[146] & b[47])^(a[145] & b[48])^(a[144] & b[49])^(a[143] & b[50])^(a[142] & b[51])^(a[141] & b[52])^(a[140] & b[53])^(a[139] & b[54])^(a[138] & b[55])^(a[137] & b[56])^(a[136] & b[57])^(a[135] & b[58])^(a[134] & b[59])^(a[133] & b[60])^(a[132] & b[61])^(a[131] & b[62])^(a[130] & b[63])^(a[129] & b[64])^(a[128] & b[65])^(a[127] & b[66])^(a[126] & b[67])^(a[125] & b[68])^(a[124] & b[69])^(a[123] & b[70])^(a[122] & b[71])^(a[121] & b[72])^(a[120] & b[73])^(a[119] & b[74])^(a[118] & b[75])^(a[117] & b[76])^(a[116] & b[77])^(a[115] & b[78])^(a[114] & b[79])^(a[113] & b[80])^(a[112] & b[81])^(a[111] & b[82])^(a[110] & b[83])^(a[109] & b[84])^(a[108] & b[85])^(a[107] & b[86])^(a[106] & b[87])^(a[105] & b[88])^(a[104] & b[89])^(a[103] & b[90])^(a[102] & b[91])^(a[101] & b[92])^(a[100] & b[93])^(a[99] & b[94])^(a[98] & b[95])^(a[97] & b[96])^(a[96] & b[97])^(a[95] & b[98])^(a[94] & b[99])^(a[93] & b[100])^(a[92] & b[101])^(a[91] & b[102])^(a[90] & b[103])^(a[89] & b[104])^(a[88] & b[105])^(a[87] & b[106])^(a[86] & b[107])^(a[85] & b[108])^(a[84] & b[109])^(a[83] & b[110])^(a[82] & b[111])^(a[81] & b[112])^(a[80] & b[113])^(a[79] & b[114])^(a[78] & b[115])^(a[77] & b[116])^(a[76] & b[117])^(a[75] & b[118])^(a[74] & b[119])^(a[73] & b[120])^(a[72] & b[121])^(a[71] & b[122])^(a[70] & b[123])^(a[69] & b[124])^(a[68] & b[125])^(a[67] & b[126])^(a[66] & b[127])^(a[65] & b[128])^(a[64] & b[129])^(a[63] & b[130])^(a[62] & b[131])^(a[61] & b[132])^(a[60] & b[133])^(a[59] & b[134])^(a[58] & b[135])^(a[57] & b[136])^(a[56] & b[137])^(a[55] & b[138])^(a[54] & b[139])^(a[53] & b[140])^(a[52] & b[141])^(a[51] & b[142])^(a[50] & b[143])^(a[49] & b[144])^(a[48] & b[145])^(a[47] & b[146])^(a[46] & b[147])^(a[45] & b[148])^(a[44] & b[149])^(a[43] & b[150])^(a[42] & b[151])^(a[41] & b[152])^(a[40] & b[153])^(a[39] & b[154])^(a[38] & b[155])^(a[37] & b[156])^(a[36] & b[157])^(a[35] & b[158])^(a[34] & b[159])^(a[33] & b[160])^(a[32] & b[161])^(a[31] & b[162])^(a[30] & b[163])^(a[29] & b[164])^(a[28] & b[165])^(a[27] & b[166])^(a[26] & b[167])^(a[25] & b[168])^(a[24] & b[169])^(a[23] & b[170])^(a[22] & b[171])^(a[21] & b[172])^(a[20] & b[173])^(a[19] & b[174])^(a[18] & b[175])^(a[17] & b[176])^(a[16] & b[177])^(a[15] & b[178])^(a[14] & b[179])^(a[13] & b[180])^(a[12] & b[181])^(a[11] & b[182])^(a[10] & b[183])^(a[9] & b[184])^(a[8] & b[185])^(a[7] & b[186])^(a[6] & b[187])^(a[5] & b[188])^(a[4] & b[189])^(a[3] & b[190])^(a[2] & b[191])^(a[1] & b[192])^(a[0] & b[193]);
assign y[194] = (a[194] & b[0])^(a[193] & b[1])^(a[192] & b[2])^(a[191] & b[3])^(a[190] & b[4])^(a[189] & b[5])^(a[188] & b[6])^(a[187] & b[7])^(a[186] & b[8])^(a[185] & b[9])^(a[184] & b[10])^(a[183] & b[11])^(a[182] & b[12])^(a[181] & b[13])^(a[180] & b[14])^(a[179] & b[15])^(a[178] & b[16])^(a[177] & b[17])^(a[176] & b[18])^(a[175] & b[19])^(a[174] & b[20])^(a[173] & b[21])^(a[172] & b[22])^(a[171] & b[23])^(a[170] & b[24])^(a[169] & b[25])^(a[168] & b[26])^(a[167] & b[27])^(a[166] & b[28])^(a[165] & b[29])^(a[164] & b[30])^(a[163] & b[31])^(a[162] & b[32])^(a[161] & b[33])^(a[160] & b[34])^(a[159] & b[35])^(a[158] & b[36])^(a[157] & b[37])^(a[156] & b[38])^(a[155] & b[39])^(a[154] & b[40])^(a[153] & b[41])^(a[152] & b[42])^(a[151] & b[43])^(a[150] & b[44])^(a[149] & b[45])^(a[148] & b[46])^(a[147] & b[47])^(a[146] & b[48])^(a[145] & b[49])^(a[144] & b[50])^(a[143] & b[51])^(a[142] & b[52])^(a[141] & b[53])^(a[140] & b[54])^(a[139] & b[55])^(a[138] & b[56])^(a[137] & b[57])^(a[136] & b[58])^(a[135] & b[59])^(a[134] & b[60])^(a[133] & b[61])^(a[132] & b[62])^(a[131] & b[63])^(a[130] & b[64])^(a[129] & b[65])^(a[128] & b[66])^(a[127] & b[67])^(a[126] & b[68])^(a[125] & b[69])^(a[124] & b[70])^(a[123] & b[71])^(a[122] & b[72])^(a[121] & b[73])^(a[120] & b[74])^(a[119] & b[75])^(a[118] & b[76])^(a[117] & b[77])^(a[116] & b[78])^(a[115] & b[79])^(a[114] & b[80])^(a[113] & b[81])^(a[112] & b[82])^(a[111] & b[83])^(a[110] & b[84])^(a[109] & b[85])^(a[108] & b[86])^(a[107] & b[87])^(a[106] & b[88])^(a[105] & b[89])^(a[104] & b[90])^(a[103] & b[91])^(a[102] & b[92])^(a[101] & b[93])^(a[100] & b[94])^(a[99] & b[95])^(a[98] & b[96])^(a[97] & b[97])^(a[96] & b[98])^(a[95] & b[99])^(a[94] & b[100])^(a[93] & b[101])^(a[92] & b[102])^(a[91] & b[103])^(a[90] & b[104])^(a[89] & b[105])^(a[88] & b[106])^(a[87] & b[107])^(a[86] & b[108])^(a[85] & b[109])^(a[84] & b[110])^(a[83] & b[111])^(a[82] & b[112])^(a[81] & b[113])^(a[80] & b[114])^(a[79] & b[115])^(a[78] & b[116])^(a[77] & b[117])^(a[76] & b[118])^(a[75] & b[119])^(a[74] & b[120])^(a[73] & b[121])^(a[72] & b[122])^(a[71] & b[123])^(a[70] & b[124])^(a[69] & b[125])^(a[68] & b[126])^(a[67] & b[127])^(a[66] & b[128])^(a[65] & b[129])^(a[64] & b[130])^(a[63] & b[131])^(a[62] & b[132])^(a[61] & b[133])^(a[60] & b[134])^(a[59] & b[135])^(a[58] & b[136])^(a[57] & b[137])^(a[56] & b[138])^(a[55] & b[139])^(a[54] & b[140])^(a[53] & b[141])^(a[52] & b[142])^(a[51] & b[143])^(a[50] & b[144])^(a[49] & b[145])^(a[48] & b[146])^(a[47] & b[147])^(a[46] & b[148])^(a[45] & b[149])^(a[44] & b[150])^(a[43] & b[151])^(a[42] & b[152])^(a[41] & b[153])^(a[40] & b[154])^(a[39] & b[155])^(a[38] & b[156])^(a[37] & b[157])^(a[36] & b[158])^(a[35] & b[159])^(a[34] & b[160])^(a[33] & b[161])^(a[32] & b[162])^(a[31] & b[163])^(a[30] & b[164])^(a[29] & b[165])^(a[28] & b[166])^(a[27] & b[167])^(a[26] & b[168])^(a[25] & b[169])^(a[24] & b[170])^(a[23] & b[171])^(a[22] & b[172])^(a[21] & b[173])^(a[20] & b[174])^(a[19] & b[175])^(a[18] & b[176])^(a[17] & b[177])^(a[16] & b[178])^(a[15] & b[179])^(a[14] & b[180])^(a[13] & b[181])^(a[12] & b[182])^(a[11] & b[183])^(a[10] & b[184])^(a[9] & b[185])^(a[8] & b[186])^(a[7] & b[187])^(a[6] & b[188])^(a[5] & b[189])^(a[4] & b[190])^(a[3] & b[191])^(a[2] & b[192])^(a[1] & b[193])^(a[0] & b[194]);
assign y[195] = (a[195] & b[0])^(a[194] & b[1])^(a[193] & b[2])^(a[192] & b[3])^(a[191] & b[4])^(a[190] & b[5])^(a[189] & b[6])^(a[188] & b[7])^(a[187] & b[8])^(a[186] & b[9])^(a[185] & b[10])^(a[184] & b[11])^(a[183] & b[12])^(a[182] & b[13])^(a[181] & b[14])^(a[180] & b[15])^(a[179] & b[16])^(a[178] & b[17])^(a[177] & b[18])^(a[176] & b[19])^(a[175] & b[20])^(a[174] & b[21])^(a[173] & b[22])^(a[172] & b[23])^(a[171] & b[24])^(a[170] & b[25])^(a[169] & b[26])^(a[168] & b[27])^(a[167] & b[28])^(a[166] & b[29])^(a[165] & b[30])^(a[164] & b[31])^(a[163] & b[32])^(a[162] & b[33])^(a[161] & b[34])^(a[160] & b[35])^(a[159] & b[36])^(a[158] & b[37])^(a[157] & b[38])^(a[156] & b[39])^(a[155] & b[40])^(a[154] & b[41])^(a[153] & b[42])^(a[152] & b[43])^(a[151] & b[44])^(a[150] & b[45])^(a[149] & b[46])^(a[148] & b[47])^(a[147] & b[48])^(a[146] & b[49])^(a[145] & b[50])^(a[144] & b[51])^(a[143] & b[52])^(a[142] & b[53])^(a[141] & b[54])^(a[140] & b[55])^(a[139] & b[56])^(a[138] & b[57])^(a[137] & b[58])^(a[136] & b[59])^(a[135] & b[60])^(a[134] & b[61])^(a[133] & b[62])^(a[132] & b[63])^(a[131] & b[64])^(a[130] & b[65])^(a[129] & b[66])^(a[128] & b[67])^(a[127] & b[68])^(a[126] & b[69])^(a[125] & b[70])^(a[124] & b[71])^(a[123] & b[72])^(a[122] & b[73])^(a[121] & b[74])^(a[120] & b[75])^(a[119] & b[76])^(a[118] & b[77])^(a[117] & b[78])^(a[116] & b[79])^(a[115] & b[80])^(a[114] & b[81])^(a[113] & b[82])^(a[112] & b[83])^(a[111] & b[84])^(a[110] & b[85])^(a[109] & b[86])^(a[108] & b[87])^(a[107] & b[88])^(a[106] & b[89])^(a[105] & b[90])^(a[104] & b[91])^(a[103] & b[92])^(a[102] & b[93])^(a[101] & b[94])^(a[100] & b[95])^(a[99] & b[96])^(a[98] & b[97])^(a[97] & b[98])^(a[96] & b[99])^(a[95] & b[100])^(a[94] & b[101])^(a[93] & b[102])^(a[92] & b[103])^(a[91] & b[104])^(a[90] & b[105])^(a[89] & b[106])^(a[88] & b[107])^(a[87] & b[108])^(a[86] & b[109])^(a[85] & b[110])^(a[84] & b[111])^(a[83] & b[112])^(a[82] & b[113])^(a[81] & b[114])^(a[80] & b[115])^(a[79] & b[116])^(a[78] & b[117])^(a[77] & b[118])^(a[76] & b[119])^(a[75] & b[120])^(a[74] & b[121])^(a[73] & b[122])^(a[72] & b[123])^(a[71] & b[124])^(a[70] & b[125])^(a[69] & b[126])^(a[68] & b[127])^(a[67] & b[128])^(a[66] & b[129])^(a[65] & b[130])^(a[64] & b[131])^(a[63] & b[132])^(a[62] & b[133])^(a[61] & b[134])^(a[60] & b[135])^(a[59] & b[136])^(a[58] & b[137])^(a[57] & b[138])^(a[56] & b[139])^(a[55] & b[140])^(a[54] & b[141])^(a[53] & b[142])^(a[52] & b[143])^(a[51] & b[144])^(a[50] & b[145])^(a[49] & b[146])^(a[48] & b[147])^(a[47] & b[148])^(a[46] & b[149])^(a[45] & b[150])^(a[44] & b[151])^(a[43] & b[152])^(a[42] & b[153])^(a[41] & b[154])^(a[40] & b[155])^(a[39] & b[156])^(a[38] & b[157])^(a[37] & b[158])^(a[36] & b[159])^(a[35] & b[160])^(a[34] & b[161])^(a[33] & b[162])^(a[32] & b[163])^(a[31] & b[164])^(a[30] & b[165])^(a[29] & b[166])^(a[28] & b[167])^(a[27] & b[168])^(a[26] & b[169])^(a[25] & b[170])^(a[24] & b[171])^(a[23] & b[172])^(a[22] & b[173])^(a[21] & b[174])^(a[20] & b[175])^(a[19] & b[176])^(a[18] & b[177])^(a[17] & b[178])^(a[16] & b[179])^(a[15] & b[180])^(a[14] & b[181])^(a[13] & b[182])^(a[12] & b[183])^(a[11] & b[184])^(a[10] & b[185])^(a[9] & b[186])^(a[8] & b[187])^(a[7] & b[188])^(a[6] & b[189])^(a[5] & b[190])^(a[4] & b[191])^(a[3] & b[192])^(a[2] & b[193])^(a[1] & b[194])^(a[0] & b[195]);
assign y[196] = (a[196] & b[0])^(a[195] & b[1])^(a[194] & b[2])^(a[193] & b[3])^(a[192] & b[4])^(a[191] & b[5])^(a[190] & b[6])^(a[189] & b[7])^(a[188] & b[8])^(a[187] & b[9])^(a[186] & b[10])^(a[185] & b[11])^(a[184] & b[12])^(a[183] & b[13])^(a[182] & b[14])^(a[181] & b[15])^(a[180] & b[16])^(a[179] & b[17])^(a[178] & b[18])^(a[177] & b[19])^(a[176] & b[20])^(a[175] & b[21])^(a[174] & b[22])^(a[173] & b[23])^(a[172] & b[24])^(a[171] & b[25])^(a[170] & b[26])^(a[169] & b[27])^(a[168] & b[28])^(a[167] & b[29])^(a[166] & b[30])^(a[165] & b[31])^(a[164] & b[32])^(a[163] & b[33])^(a[162] & b[34])^(a[161] & b[35])^(a[160] & b[36])^(a[159] & b[37])^(a[158] & b[38])^(a[157] & b[39])^(a[156] & b[40])^(a[155] & b[41])^(a[154] & b[42])^(a[153] & b[43])^(a[152] & b[44])^(a[151] & b[45])^(a[150] & b[46])^(a[149] & b[47])^(a[148] & b[48])^(a[147] & b[49])^(a[146] & b[50])^(a[145] & b[51])^(a[144] & b[52])^(a[143] & b[53])^(a[142] & b[54])^(a[141] & b[55])^(a[140] & b[56])^(a[139] & b[57])^(a[138] & b[58])^(a[137] & b[59])^(a[136] & b[60])^(a[135] & b[61])^(a[134] & b[62])^(a[133] & b[63])^(a[132] & b[64])^(a[131] & b[65])^(a[130] & b[66])^(a[129] & b[67])^(a[128] & b[68])^(a[127] & b[69])^(a[126] & b[70])^(a[125] & b[71])^(a[124] & b[72])^(a[123] & b[73])^(a[122] & b[74])^(a[121] & b[75])^(a[120] & b[76])^(a[119] & b[77])^(a[118] & b[78])^(a[117] & b[79])^(a[116] & b[80])^(a[115] & b[81])^(a[114] & b[82])^(a[113] & b[83])^(a[112] & b[84])^(a[111] & b[85])^(a[110] & b[86])^(a[109] & b[87])^(a[108] & b[88])^(a[107] & b[89])^(a[106] & b[90])^(a[105] & b[91])^(a[104] & b[92])^(a[103] & b[93])^(a[102] & b[94])^(a[101] & b[95])^(a[100] & b[96])^(a[99] & b[97])^(a[98] & b[98])^(a[97] & b[99])^(a[96] & b[100])^(a[95] & b[101])^(a[94] & b[102])^(a[93] & b[103])^(a[92] & b[104])^(a[91] & b[105])^(a[90] & b[106])^(a[89] & b[107])^(a[88] & b[108])^(a[87] & b[109])^(a[86] & b[110])^(a[85] & b[111])^(a[84] & b[112])^(a[83] & b[113])^(a[82] & b[114])^(a[81] & b[115])^(a[80] & b[116])^(a[79] & b[117])^(a[78] & b[118])^(a[77] & b[119])^(a[76] & b[120])^(a[75] & b[121])^(a[74] & b[122])^(a[73] & b[123])^(a[72] & b[124])^(a[71] & b[125])^(a[70] & b[126])^(a[69] & b[127])^(a[68] & b[128])^(a[67] & b[129])^(a[66] & b[130])^(a[65] & b[131])^(a[64] & b[132])^(a[63] & b[133])^(a[62] & b[134])^(a[61] & b[135])^(a[60] & b[136])^(a[59] & b[137])^(a[58] & b[138])^(a[57] & b[139])^(a[56] & b[140])^(a[55] & b[141])^(a[54] & b[142])^(a[53] & b[143])^(a[52] & b[144])^(a[51] & b[145])^(a[50] & b[146])^(a[49] & b[147])^(a[48] & b[148])^(a[47] & b[149])^(a[46] & b[150])^(a[45] & b[151])^(a[44] & b[152])^(a[43] & b[153])^(a[42] & b[154])^(a[41] & b[155])^(a[40] & b[156])^(a[39] & b[157])^(a[38] & b[158])^(a[37] & b[159])^(a[36] & b[160])^(a[35] & b[161])^(a[34] & b[162])^(a[33] & b[163])^(a[32] & b[164])^(a[31] & b[165])^(a[30] & b[166])^(a[29] & b[167])^(a[28] & b[168])^(a[27] & b[169])^(a[26] & b[170])^(a[25] & b[171])^(a[24] & b[172])^(a[23] & b[173])^(a[22] & b[174])^(a[21] & b[175])^(a[20] & b[176])^(a[19] & b[177])^(a[18] & b[178])^(a[17] & b[179])^(a[16] & b[180])^(a[15] & b[181])^(a[14] & b[182])^(a[13] & b[183])^(a[12] & b[184])^(a[11] & b[185])^(a[10] & b[186])^(a[9] & b[187])^(a[8] & b[188])^(a[7] & b[189])^(a[6] & b[190])^(a[5] & b[191])^(a[4] & b[192])^(a[3] & b[193])^(a[2] & b[194])^(a[1] & b[195])^(a[0] & b[196]);
assign y[197] = (a[197] & b[0])^(a[196] & b[1])^(a[195] & b[2])^(a[194] & b[3])^(a[193] & b[4])^(a[192] & b[5])^(a[191] & b[6])^(a[190] & b[7])^(a[189] & b[8])^(a[188] & b[9])^(a[187] & b[10])^(a[186] & b[11])^(a[185] & b[12])^(a[184] & b[13])^(a[183] & b[14])^(a[182] & b[15])^(a[181] & b[16])^(a[180] & b[17])^(a[179] & b[18])^(a[178] & b[19])^(a[177] & b[20])^(a[176] & b[21])^(a[175] & b[22])^(a[174] & b[23])^(a[173] & b[24])^(a[172] & b[25])^(a[171] & b[26])^(a[170] & b[27])^(a[169] & b[28])^(a[168] & b[29])^(a[167] & b[30])^(a[166] & b[31])^(a[165] & b[32])^(a[164] & b[33])^(a[163] & b[34])^(a[162] & b[35])^(a[161] & b[36])^(a[160] & b[37])^(a[159] & b[38])^(a[158] & b[39])^(a[157] & b[40])^(a[156] & b[41])^(a[155] & b[42])^(a[154] & b[43])^(a[153] & b[44])^(a[152] & b[45])^(a[151] & b[46])^(a[150] & b[47])^(a[149] & b[48])^(a[148] & b[49])^(a[147] & b[50])^(a[146] & b[51])^(a[145] & b[52])^(a[144] & b[53])^(a[143] & b[54])^(a[142] & b[55])^(a[141] & b[56])^(a[140] & b[57])^(a[139] & b[58])^(a[138] & b[59])^(a[137] & b[60])^(a[136] & b[61])^(a[135] & b[62])^(a[134] & b[63])^(a[133] & b[64])^(a[132] & b[65])^(a[131] & b[66])^(a[130] & b[67])^(a[129] & b[68])^(a[128] & b[69])^(a[127] & b[70])^(a[126] & b[71])^(a[125] & b[72])^(a[124] & b[73])^(a[123] & b[74])^(a[122] & b[75])^(a[121] & b[76])^(a[120] & b[77])^(a[119] & b[78])^(a[118] & b[79])^(a[117] & b[80])^(a[116] & b[81])^(a[115] & b[82])^(a[114] & b[83])^(a[113] & b[84])^(a[112] & b[85])^(a[111] & b[86])^(a[110] & b[87])^(a[109] & b[88])^(a[108] & b[89])^(a[107] & b[90])^(a[106] & b[91])^(a[105] & b[92])^(a[104] & b[93])^(a[103] & b[94])^(a[102] & b[95])^(a[101] & b[96])^(a[100] & b[97])^(a[99] & b[98])^(a[98] & b[99])^(a[97] & b[100])^(a[96] & b[101])^(a[95] & b[102])^(a[94] & b[103])^(a[93] & b[104])^(a[92] & b[105])^(a[91] & b[106])^(a[90] & b[107])^(a[89] & b[108])^(a[88] & b[109])^(a[87] & b[110])^(a[86] & b[111])^(a[85] & b[112])^(a[84] & b[113])^(a[83] & b[114])^(a[82] & b[115])^(a[81] & b[116])^(a[80] & b[117])^(a[79] & b[118])^(a[78] & b[119])^(a[77] & b[120])^(a[76] & b[121])^(a[75] & b[122])^(a[74] & b[123])^(a[73] & b[124])^(a[72] & b[125])^(a[71] & b[126])^(a[70] & b[127])^(a[69] & b[128])^(a[68] & b[129])^(a[67] & b[130])^(a[66] & b[131])^(a[65] & b[132])^(a[64] & b[133])^(a[63] & b[134])^(a[62] & b[135])^(a[61] & b[136])^(a[60] & b[137])^(a[59] & b[138])^(a[58] & b[139])^(a[57] & b[140])^(a[56] & b[141])^(a[55] & b[142])^(a[54] & b[143])^(a[53] & b[144])^(a[52] & b[145])^(a[51] & b[146])^(a[50] & b[147])^(a[49] & b[148])^(a[48] & b[149])^(a[47] & b[150])^(a[46] & b[151])^(a[45] & b[152])^(a[44] & b[153])^(a[43] & b[154])^(a[42] & b[155])^(a[41] & b[156])^(a[40] & b[157])^(a[39] & b[158])^(a[38] & b[159])^(a[37] & b[160])^(a[36] & b[161])^(a[35] & b[162])^(a[34] & b[163])^(a[33] & b[164])^(a[32] & b[165])^(a[31] & b[166])^(a[30] & b[167])^(a[29] & b[168])^(a[28] & b[169])^(a[27] & b[170])^(a[26] & b[171])^(a[25] & b[172])^(a[24] & b[173])^(a[23] & b[174])^(a[22] & b[175])^(a[21] & b[176])^(a[20] & b[177])^(a[19] & b[178])^(a[18] & b[179])^(a[17] & b[180])^(a[16] & b[181])^(a[15] & b[182])^(a[14] & b[183])^(a[13] & b[184])^(a[12] & b[185])^(a[11] & b[186])^(a[10] & b[187])^(a[9] & b[188])^(a[8] & b[189])^(a[7] & b[190])^(a[6] & b[191])^(a[5] & b[192])^(a[4] & b[193])^(a[3] & b[194])^(a[2] & b[195])^(a[1] & b[196])^(a[0] & b[197]);
assign y[198] = (a[198] & b[0])^(a[197] & b[1])^(a[196] & b[2])^(a[195] & b[3])^(a[194] & b[4])^(a[193] & b[5])^(a[192] & b[6])^(a[191] & b[7])^(a[190] & b[8])^(a[189] & b[9])^(a[188] & b[10])^(a[187] & b[11])^(a[186] & b[12])^(a[185] & b[13])^(a[184] & b[14])^(a[183] & b[15])^(a[182] & b[16])^(a[181] & b[17])^(a[180] & b[18])^(a[179] & b[19])^(a[178] & b[20])^(a[177] & b[21])^(a[176] & b[22])^(a[175] & b[23])^(a[174] & b[24])^(a[173] & b[25])^(a[172] & b[26])^(a[171] & b[27])^(a[170] & b[28])^(a[169] & b[29])^(a[168] & b[30])^(a[167] & b[31])^(a[166] & b[32])^(a[165] & b[33])^(a[164] & b[34])^(a[163] & b[35])^(a[162] & b[36])^(a[161] & b[37])^(a[160] & b[38])^(a[159] & b[39])^(a[158] & b[40])^(a[157] & b[41])^(a[156] & b[42])^(a[155] & b[43])^(a[154] & b[44])^(a[153] & b[45])^(a[152] & b[46])^(a[151] & b[47])^(a[150] & b[48])^(a[149] & b[49])^(a[148] & b[50])^(a[147] & b[51])^(a[146] & b[52])^(a[145] & b[53])^(a[144] & b[54])^(a[143] & b[55])^(a[142] & b[56])^(a[141] & b[57])^(a[140] & b[58])^(a[139] & b[59])^(a[138] & b[60])^(a[137] & b[61])^(a[136] & b[62])^(a[135] & b[63])^(a[134] & b[64])^(a[133] & b[65])^(a[132] & b[66])^(a[131] & b[67])^(a[130] & b[68])^(a[129] & b[69])^(a[128] & b[70])^(a[127] & b[71])^(a[126] & b[72])^(a[125] & b[73])^(a[124] & b[74])^(a[123] & b[75])^(a[122] & b[76])^(a[121] & b[77])^(a[120] & b[78])^(a[119] & b[79])^(a[118] & b[80])^(a[117] & b[81])^(a[116] & b[82])^(a[115] & b[83])^(a[114] & b[84])^(a[113] & b[85])^(a[112] & b[86])^(a[111] & b[87])^(a[110] & b[88])^(a[109] & b[89])^(a[108] & b[90])^(a[107] & b[91])^(a[106] & b[92])^(a[105] & b[93])^(a[104] & b[94])^(a[103] & b[95])^(a[102] & b[96])^(a[101] & b[97])^(a[100] & b[98])^(a[99] & b[99])^(a[98] & b[100])^(a[97] & b[101])^(a[96] & b[102])^(a[95] & b[103])^(a[94] & b[104])^(a[93] & b[105])^(a[92] & b[106])^(a[91] & b[107])^(a[90] & b[108])^(a[89] & b[109])^(a[88] & b[110])^(a[87] & b[111])^(a[86] & b[112])^(a[85] & b[113])^(a[84] & b[114])^(a[83] & b[115])^(a[82] & b[116])^(a[81] & b[117])^(a[80] & b[118])^(a[79] & b[119])^(a[78] & b[120])^(a[77] & b[121])^(a[76] & b[122])^(a[75] & b[123])^(a[74] & b[124])^(a[73] & b[125])^(a[72] & b[126])^(a[71] & b[127])^(a[70] & b[128])^(a[69] & b[129])^(a[68] & b[130])^(a[67] & b[131])^(a[66] & b[132])^(a[65] & b[133])^(a[64] & b[134])^(a[63] & b[135])^(a[62] & b[136])^(a[61] & b[137])^(a[60] & b[138])^(a[59] & b[139])^(a[58] & b[140])^(a[57] & b[141])^(a[56] & b[142])^(a[55] & b[143])^(a[54] & b[144])^(a[53] & b[145])^(a[52] & b[146])^(a[51] & b[147])^(a[50] & b[148])^(a[49] & b[149])^(a[48] & b[150])^(a[47] & b[151])^(a[46] & b[152])^(a[45] & b[153])^(a[44] & b[154])^(a[43] & b[155])^(a[42] & b[156])^(a[41] & b[157])^(a[40] & b[158])^(a[39] & b[159])^(a[38] & b[160])^(a[37] & b[161])^(a[36] & b[162])^(a[35] & b[163])^(a[34] & b[164])^(a[33] & b[165])^(a[32] & b[166])^(a[31] & b[167])^(a[30] & b[168])^(a[29] & b[169])^(a[28] & b[170])^(a[27] & b[171])^(a[26] & b[172])^(a[25] & b[173])^(a[24] & b[174])^(a[23] & b[175])^(a[22] & b[176])^(a[21] & b[177])^(a[20] & b[178])^(a[19] & b[179])^(a[18] & b[180])^(a[17] & b[181])^(a[16] & b[182])^(a[15] & b[183])^(a[14] & b[184])^(a[13] & b[185])^(a[12] & b[186])^(a[11] & b[187])^(a[10] & b[188])^(a[9] & b[189])^(a[8] & b[190])^(a[7] & b[191])^(a[6] & b[192])^(a[5] & b[193])^(a[4] & b[194])^(a[3] & b[195])^(a[2] & b[196])^(a[1] & b[197])^(a[0] & b[198]);
assign y[199] = (a[199] & b[0])^(a[198] & b[1])^(a[197] & b[2])^(a[196] & b[3])^(a[195] & b[4])^(a[194] & b[5])^(a[193] & b[6])^(a[192] & b[7])^(a[191] & b[8])^(a[190] & b[9])^(a[189] & b[10])^(a[188] & b[11])^(a[187] & b[12])^(a[186] & b[13])^(a[185] & b[14])^(a[184] & b[15])^(a[183] & b[16])^(a[182] & b[17])^(a[181] & b[18])^(a[180] & b[19])^(a[179] & b[20])^(a[178] & b[21])^(a[177] & b[22])^(a[176] & b[23])^(a[175] & b[24])^(a[174] & b[25])^(a[173] & b[26])^(a[172] & b[27])^(a[171] & b[28])^(a[170] & b[29])^(a[169] & b[30])^(a[168] & b[31])^(a[167] & b[32])^(a[166] & b[33])^(a[165] & b[34])^(a[164] & b[35])^(a[163] & b[36])^(a[162] & b[37])^(a[161] & b[38])^(a[160] & b[39])^(a[159] & b[40])^(a[158] & b[41])^(a[157] & b[42])^(a[156] & b[43])^(a[155] & b[44])^(a[154] & b[45])^(a[153] & b[46])^(a[152] & b[47])^(a[151] & b[48])^(a[150] & b[49])^(a[149] & b[50])^(a[148] & b[51])^(a[147] & b[52])^(a[146] & b[53])^(a[145] & b[54])^(a[144] & b[55])^(a[143] & b[56])^(a[142] & b[57])^(a[141] & b[58])^(a[140] & b[59])^(a[139] & b[60])^(a[138] & b[61])^(a[137] & b[62])^(a[136] & b[63])^(a[135] & b[64])^(a[134] & b[65])^(a[133] & b[66])^(a[132] & b[67])^(a[131] & b[68])^(a[130] & b[69])^(a[129] & b[70])^(a[128] & b[71])^(a[127] & b[72])^(a[126] & b[73])^(a[125] & b[74])^(a[124] & b[75])^(a[123] & b[76])^(a[122] & b[77])^(a[121] & b[78])^(a[120] & b[79])^(a[119] & b[80])^(a[118] & b[81])^(a[117] & b[82])^(a[116] & b[83])^(a[115] & b[84])^(a[114] & b[85])^(a[113] & b[86])^(a[112] & b[87])^(a[111] & b[88])^(a[110] & b[89])^(a[109] & b[90])^(a[108] & b[91])^(a[107] & b[92])^(a[106] & b[93])^(a[105] & b[94])^(a[104] & b[95])^(a[103] & b[96])^(a[102] & b[97])^(a[101] & b[98])^(a[100] & b[99])^(a[99] & b[100])^(a[98] & b[101])^(a[97] & b[102])^(a[96] & b[103])^(a[95] & b[104])^(a[94] & b[105])^(a[93] & b[106])^(a[92] & b[107])^(a[91] & b[108])^(a[90] & b[109])^(a[89] & b[110])^(a[88] & b[111])^(a[87] & b[112])^(a[86] & b[113])^(a[85] & b[114])^(a[84] & b[115])^(a[83] & b[116])^(a[82] & b[117])^(a[81] & b[118])^(a[80] & b[119])^(a[79] & b[120])^(a[78] & b[121])^(a[77] & b[122])^(a[76] & b[123])^(a[75] & b[124])^(a[74] & b[125])^(a[73] & b[126])^(a[72] & b[127])^(a[71] & b[128])^(a[70] & b[129])^(a[69] & b[130])^(a[68] & b[131])^(a[67] & b[132])^(a[66] & b[133])^(a[65] & b[134])^(a[64] & b[135])^(a[63] & b[136])^(a[62] & b[137])^(a[61] & b[138])^(a[60] & b[139])^(a[59] & b[140])^(a[58] & b[141])^(a[57] & b[142])^(a[56] & b[143])^(a[55] & b[144])^(a[54] & b[145])^(a[53] & b[146])^(a[52] & b[147])^(a[51] & b[148])^(a[50] & b[149])^(a[49] & b[150])^(a[48] & b[151])^(a[47] & b[152])^(a[46] & b[153])^(a[45] & b[154])^(a[44] & b[155])^(a[43] & b[156])^(a[42] & b[157])^(a[41] & b[158])^(a[40] & b[159])^(a[39] & b[160])^(a[38] & b[161])^(a[37] & b[162])^(a[36] & b[163])^(a[35] & b[164])^(a[34] & b[165])^(a[33] & b[166])^(a[32] & b[167])^(a[31] & b[168])^(a[30] & b[169])^(a[29] & b[170])^(a[28] & b[171])^(a[27] & b[172])^(a[26] & b[173])^(a[25] & b[174])^(a[24] & b[175])^(a[23] & b[176])^(a[22] & b[177])^(a[21] & b[178])^(a[20] & b[179])^(a[19] & b[180])^(a[18] & b[181])^(a[17] & b[182])^(a[16] & b[183])^(a[15] & b[184])^(a[14] & b[185])^(a[13] & b[186])^(a[12] & b[187])^(a[11] & b[188])^(a[10] & b[189])^(a[9] & b[190])^(a[8] & b[191])^(a[7] & b[192])^(a[6] & b[193])^(a[5] & b[194])^(a[4] & b[195])^(a[3] & b[196])^(a[2] & b[197])^(a[1] & b[198])^(a[0] & b[199]);
assign y[200] = (a[200] & b[0])^(a[199] & b[1])^(a[198] & b[2])^(a[197] & b[3])^(a[196] & b[4])^(a[195] & b[5])^(a[194] & b[6])^(a[193] & b[7])^(a[192] & b[8])^(a[191] & b[9])^(a[190] & b[10])^(a[189] & b[11])^(a[188] & b[12])^(a[187] & b[13])^(a[186] & b[14])^(a[185] & b[15])^(a[184] & b[16])^(a[183] & b[17])^(a[182] & b[18])^(a[181] & b[19])^(a[180] & b[20])^(a[179] & b[21])^(a[178] & b[22])^(a[177] & b[23])^(a[176] & b[24])^(a[175] & b[25])^(a[174] & b[26])^(a[173] & b[27])^(a[172] & b[28])^(a[171] & b[29])^(a[170] & b[30])^(a[169] & b[31])^(a[168] & b[32])^(a[167] & b[33])^(a[166] & b[34])^(a[165] & b[35])^(a[164] & b[36])^(a[163] & b[37])^(a[162] & b[38])^(a[161] & b[39])^(a[160] & b[40])^(a[159] & b[41])^(a[158] & b[42])^(a[157] & b[43])^(a[156] & b[44])^(a[155] & b[45])^(a[154] & b[46])^(a[153] & b[47])^(a[152] & b[48])^(a[151] & b[49])^(a[150] & b[50])^(a[149] & b[51])^(a[148] & b[52])^(a[147] & b[53])^(a[146] & b[54])^(a[145] & b[55])^(a[144] & b[56])^(a[143] & b[57])^(a[142] & b[58])^(a[141] & b[59])^(a[140] & b[60])^(a[139] & b[61])^(a[138] & b[62])^(a[137] & b[63])^(a[136] & b[64])^(a[135] & b[65])^(a[134] & b[66])^(a[133] & b[67])^(a[132] & b[68])^(a[131] & b[69])^(a[130] & b[70])^(a[129] & b[71])^(a[128] & b[72])^(a[127] & b[73])^(a[126] & b[74])^(a[125] & b[75])^(a[124] & b[76])^(a[123] & b[77])^(a[122] & b[78])^(a[121] & b[79])^(a[120] & b[80])^(a[119] & b[81])^(a[118] & b[82])^(a[117] & b[83])^(a[116] & b[84])^(a[115] & b[85])^(a[114] & b[86])^(a[113] & b[87])^(a[112] & b[88])^(a[111] & b[89])^(a[110] & b[90])^(a[109] & b[91])^(a[108] & b[92])^(a[107] & b[93])^(a[106] & b[94])^(a[105] & b[95])^(a[104] & b[96])^(a[103] & b[97])^(a[102] & b[98])^(a[101] & b[99])^(a[100] & b[100])^(a[99] & b[101])^(a[98] & b[102])^(a[97] & b[103])^(a[96] & b[104])^(a[95] & b[105])^(a[94] & b[106])^(a[93] & b[107])^(a[92] & b[108])^(a[91] & b[109])^(a[90] & b[110])^(a[89] & b[111])^(a[88] & b[112])^(a[87] & b[113])^(a[86] & b[114])^(a[85] & b[115])^(a[84] & b[116])^(a[83] & b[117])^(a[82] & b[118])^(a[81] & b[119])^(a[80] & b[120])^(a[79] & b[121])^(a[78] & b[122])^(a[77] & b[123])^(a[76] & b[124])^(a[75] & b[125])^(a[74] & b[126])^(a[73] & b[127])^(a[72] & b[128])^(a[71] & b[129])^(a[70] & b[130])^(a[69] & b[131])^(a[68] & b[132])^(a[67] & b[133])^(a[66] & b[134])^(a[65] & b[135])^(a[64] & b[136])^(a[63] & b[137])^(a[62] & b[138])^(a[61] & b[139])^(a[60] & b[140])^(a[59] & b[141])^(a[58] & b[142])^(a[57] & b[143])^(a[56] & b[144])^(a[55] & b[145])^(a[54] & b[146])^(a[53] & b[147])^(a[52] & b[148])^(a[51] & b[149])^(a[50] & b[150])^(a[49] & b[151])^(a[48] & b[152])^(a[47] & b[153])^(a[46] & b[154])^(a[45] & b[155])^(a[44] & b[156])^(a[43] & b[157])^(a[42] & b[158])^(a[41] & b[159])^(a[40] & b[160])^(a[39] & b[161])^(a[38] & b[162])^(a[37] & b[163])^(a[36] & b[164])^(a[35] & b[165])^(a[34] & b[166])^(a[33] & b[167])^(a[32] & b[168])^(a[31] & b[169])^(a[30] & b[170])^(a[29] & b[171])^(a[28] & b[172])^(a[27] & b[173])^(a[26] & b[174])^(a[25] & b[175])^(a[24] & b[176])^(a[23] & b[177])^(a[22] & b[178])^(a[21] & b[179])^(a[20] & b[180])^(a[19] & b[181])^(a[18] & b[182])^(a[17] & b[183])^(a[16] & b[184])^(a[15] & b[185])^(a[14] & b[186])^(a[13] & b[187])^(a[12] & b[188])^(a[11] & b[189])^(a[10] & b[190])^(a[9] & b[191])^(a[8] & b[192])^(a[7] & b[193])^(a[6] & b[194])^(a[5] & b[195])^(a[4] & b[196])^(a[3] & b[197])^(a[2] & b[198])^(a[1] & b[199])^(a[0] & b[200]);
assign y[201] = (a[201] & b[0])^(a[200] & b[1])^(a[199] & b[2])^(a[198] & b[3])^(a[197] & b[4])^(a[196] & b[5])^(a[195] & b[6])^(a[194] & b[7])^(a[193] & b[8])^(a[192] & b[9])^(a[191] & b[10])^(a[190] & b[11])^(a[189] & b[12])^(a[188] & b[13])^(a[187] & b[14])^(a[186] & b[15])^(a[185] & b[16])^(a[184] & b[17])^(a[183] & b[18])^(a[182] & b[19])^(a[181] & b[20])^(a[180] & b[21])^(a[179] & b[22])^(a[178] & b[23])^(a[177] & b[24])^(a[176] & b[25])^(a[175] & b[26])^(a[174] & b[27])^(a[173] & b[28])^(a[172] & b[29])^(a[171] & b[30])^(a[170] & b[31])^(a[169] & b[32])^(a[168] & b[33])^(a[167] & b[34])^(a[166] & b[35])^(a[165] & b[36])^(a[164] & b[37])^(a[163] & b[38])^(a[162] & b[39])^(a[161] & b[40])^(a[160] & b[41])^(a[159] & b[42])^(a[158] & b[43])^(a[157] & b[44])^(a[156] & b[45])^(a[155] & b[46])^(a[154] & b[47])^(a[153] & b[48])^(a[152] & b[49])^(a[151] & b[50])^(a[150] & b[51])^(a[149] & b[52])^(a[148] & b[53])^(a[147] & b[54])^(a[146] & b[55])^(a[145] & b[56])^(a[144] & b[57])^(a[143] & b[58])^(a[142] & b[59])^(a[141] & b[60])^(a[140] & b[61])^(a[139] & b[62])^(a[138] & b[63])^(a[137] & b[64])^(a[136] & b[65])^(a[135] & b[66])^(a[134] & b[67])^(a[133] & b[68])^(a[132] & b[69])^(a[131] & b[70])^(a[130] & b[71])^(a[129] & b[72])^(a[128] & b[73])^(a[127] & b[74])^(a[126] & b[75])^(a[125] & b[76])^(a[124] & b[77])^(a[123] & b[78])^(a[122] & b[79])^(a[121] & b[80])^(a[120] & b[81])^(a[119] & b[82])^(a[118] & b[83])^(a[117] & b[84])^(a[116] & b[85])^(a[115] & b[86])^(a[114] & b[87])^(a[113] & b[88])^(a[112] & b[89])^(a[111] & b[90])^(a[110] & b[91])^(a[109] & b[92])^(a[108] & b[93])^(a[107] & b[94])^(a[106] & b[95])^(a[105] & b[96])^(a[104] & b[97])^(a[103] & b[98])^(a[102] & b[99])^(a[101] & b[100])^(a[100] & b[101])^(a[99] & b[102])^(a[98] & b[103])^(a[97] & b[104])^(a[96] & b[105])^(a[95] & b[106])^(a[94] & b[107])^(a[93] & b[108])^(a[92] & b[109])^(a[91] & b[110])^(a[90] & b[111])^(a[89] & b[112])^(a[88] & b[113])^(a[87] & b[114])^(a[86] & b[115])^(a[85] & b[116])^(a[84] & b[117])^(a[83] & b[118])^(a[82] & b[119])^(a[81] & b[120])^(a[80] & b[121])^(a[79] & b[122])^(a[78] & b[123])^(a[77] & b[124])^(a[76] & b[125])^(a[75] & b[126])^(a[74] & b[127])^(a[73] & b[128])^(a[72] & b[129])^(a[71] & b[130])^(a[70] & b[131])^(a[69] & b[132])^(a[68] & b[133])^(a[67] & b[134])^(a[66] & b[135])^(a[65] & b[136])^(a[64] & b[137])^(a[63] & b[138])^(a[62] & b[139])^(a[61] & b[140])^(a[60] & b[141])^(a[59] & b[142])^(a[58] & b[143])^(a[57] & b[144])^(a[56] & b[145])^(a[55] & b[146])^(a[54] & b[147])^(a[53] & b[148])^(a[52] & b[149])^(a[51] & b[150])^(a[50] & b[151])^(a[49] & b[152])^(a[48] & b[153])^(a[47] & b[154])^(a[46] & b[155])^(a[45] & b[156])^(a[44] & b[157])^(a[43] & b[158])^(a[42] & b[159])^(a[41] & b[160])^(a[40] & b[161])^(a[39] & b[162])^(a[38] & b[163])^(a[37] & b[164])^(a[36] & b[165])^(a[35] & b[166])^(a[34] & b[167])^(a[33] & b[168])^(a[32] & b[169])^(a[31] & b[170])^(a[30] & b[171])^(a[29] & b[172])^(a[28] & b[173])^(a[27] & b[174])^(a[26] & b[175])^(a[25] & b[176])^(a[24] & b[177])^(a[23] & b[178])^(a[22] & b[179])^(a[21] & b[180])^(a[20] & b[181])^(a[19] & b[182])^(a[18] & b[183])^(a[17] & b[184])^(a[16] & b[185])^(a[15] & b[186])^(a[14] & b[187])^(a[13] & b[188])^(a[12] & b[189])^(a[11] & b[190])^(a[10] & b[191])^(a[9] & b[192])^(a[8] & b[193])^(a[7] & b[194])^(a[6] & b[195])^(a[5] & b[196])^(a[4] & b[197])^(a[3] & b[198])^(a[2] & b[199])^(a[1] & b[200])^(a[0] & b[201]);
assign y[202] = (a[202] & b[0])^(a[201] & b[1])^(a[200] & b[2])^(a[199] & b[3])^(a[198] & b[4])^(a[197] & b[5])^(a[196] & b[6])^(a[195] & b[7])^(a[194] & b[8])^(a[193] & b[9])^(a[192] & b[10])^(a[191] & b[11])^(a[190] & b[12])^(a[189] & b[13])^(a[188] & b[14])^(a[187] & b[15])^(a[186] & b[16])^(a[185] & b[17])^(a[184] & b[18])^(a[183] & b[19])^(a[182] & b[20])^(a[181] & b[21])^(a[180] & b[22])^(a[179] & b[23])^(a[178] & b[24])^(a[177] & b[25])^(a[176] & b[26])^(a[175] & b[27])^(a[174] & b[28])^(a[173] & b[29])^(a[172] & b[30])^(a[171] & b[31])^(a[170] & b[32])^(a[169] & b[33])^(a[168] & b[34])^(a[167] & b[35])^(a[166] & b[36])^(a[165] & b[37])^(a[164] & b[38])^(a[163] & b[39])^(a[162] & b[40])^(a[161] & b[41])^(a[160] & b[42])^(a[159] & b[43])^(a[158] & b[44])^(a[157] & b[45])^(a[156] & b[46])^(a[155] & b[47])^(a[154] & b[48])^(a[153] & b[49])^(a[152] & b[50])^(a[151] & b[51])^(a[150] & b[52])^(a[149] & b[53])^(a[148] & b[54])^(a[147] & b[55])^(a[146] & b[56])^(a[145] & b[57])^(a[144] & b[58])^(a[143] & b[59])^(a[142] & b[60])^(a[141] & b[61])^(a[140] & b[62])^(a[139] & b[63])^(a[138] & b[64])^(a[137] & b[65])^(a[136] & b[66])^(a[135] & b[67])^(a[134] & b[68])^(a[133] & b[69])^(a[132] & b[70])^(a[131] & b[71])^(a[130] & b[72])^(a[129] & b[73])^(a[128] & b[74])^(a[127] & b[75])^(a[126] & b[76])^(a[125] & b[77])^(a[124] & b[78])^(a[123] & b[79])^(a[122] & b[80])^(a[121] & b[81])^(a[120] & b[82])^(a[119] & b[83])^(a[118] & b[84])^(a[117] & b[85])^(a[116] & b[86])^(a[115] & b[87])^(a[114] & b[88])^(a[113] & b[89])^(a[112] & b[90])^(a[111] & b[91])^(a[110] & b[92])^(a[109] & b[93])^(a[108] & b[94])^(a[107] & b[95])^(a[106] & b[96])^(a[105] & b[97])^(a[104] & b[98])^(a[103] & b[99])^(a[102] & b[100])^(a[101] & b[101])^(a[100] & b[102])^(a[99] & b[103])^(a[98] & b[104])^(a[97] & b[105])^(a[96] & b[106])^(a[95] & b[107])^(a[94] & b[108])^(a[93] & b[109])^(a[92] & b[110])^(a[91] & b[111])^(a[90] & b[112])^(a[89] & b[113])^(a[88] & b[114])^(a[87] & b[115])^(a[86] & b[116])^(a[85] & b[117])^(a[84] & b[118])^(a[83] & b[119])^(a[82] & b[120])^(a[81] & b[121])^(a[80] & b[122])^(a[79] & b[123])^(a[78] & b[124])^(a[77] & b[125])^(a[76] & b[126])^(a[75] & b[127])^(a[74] & b[128])^(a[73] & b[129])^(a[72] & b[130])^(a[71] & b[131])^(a[70] & b[132])^(a[69] & b[133])^(a[68] & b[134])^(a[67] & b[135])^(a[66] & b[136])^(a[65] & b[137])^(a[64] & b[138])^(a[63] & b[139])^(a[62] & b[140])^(a[61] & b[141])^(a[60] & b[142])^(a[59] & b[143])^(a[58] & b[144])^(a[57] & b[145])^(a[56] & b[146])^(a[55] & b[147])^(a[54] & b[148])^(a[53] & b[149])^(a[52] & b[150])^(a[51] & b[151])^(a[50] & b[152])^(a[49] & b[153])^(a[48] & b[154])^(a[47] & b[155])^(a[46] & b[156])^(a[45] & b[157])^(a[44] & b[158])^(a[43] & b[159])^(a[42] & b[160])^(a[41] & b[161])^(a[40] & b[162])^(a[39] & b[163])^(a[38] & b[164])^(a[37] & b[165])^(a[36] & b[166])^(a[35] & b[167])^(a[34] & b[168])^(a[33] & b[169])^(a[32] & b[170])^(a[31] & b[171])^(a[30] & b[172])^(a[29] & b[173])^(a[28] & b[174])^(a[27] & b[175])^(a[26] & b[176])^(a[25] & b[177])^(a[24] & b[178])^(a[23] & b[179])^(a[22] & b[180])^(a[21] & b[181])^(a[20] & b[182])^(a[19] & b[183])^(a[18] & b[184])^(a[17] & b[185])^(a[16] & b[186])^(a[15] & b[187])^(a[14] & b[188])^(a[13] & b[189])^(a[12] & b[190])^(a[11] & b[191])^(a[10] & b[192])^(a[9] & b[193])^(a[8] & b[194])^(a[7] & b[195])^(a[6] & b[196])^(a[5] & b[197])^(a[4] & b[198])^(a[3] & b[199])^(a[2] & b[200])^(a[1] & b[201])^(a[0] & b[202]);
assign y[203] = (a[203] & b[0])^(a[202] & b[1])^(a[201] & b[2])^(a[200] & b[3])^(a[199] & b[4])^(a[198] & b[5])^(a[197] & b[6])^(a[196] & b[7])^(a[195] & b[8])^(a[194] & b[9])^(a[193] & b[10])^(a[192] & b[11])^(a[191] & b[12])^(a[190] & b[13])^(a[189] & b[14])^(a[188] & b[15])^(a[187] & b[16])^(a[186] & b[17])^(a[185] & b[18])^(a[184] & b[19])^(a[183] & b[20])^(a[182] & b[21])^(a[181] & b[22])^(a[180] & b[23])^(a[179] & b[24])^(a[178] & b[25])^(a[177] & b[26])^(a[176] & b[27])^(a[175] & b[28])^(a[174] & b[29])^(a[173] & b[30])^(a[172] & b[31])^(a[171] & b[32])^(a[170] & b[33])^(a[169] & b[34])^(a[168] & b[35])^(a[167] & b[36])^(a[166] & b[37])^(a[165] & b[38])^(a[164] & b[39])^(a[163] & b[40])^(a[162] & b[41])^(a[161] & b[42])^(a[160] & b[43])^(a[159] & b[44])^(a[158] & b[45])^(a[157] & b[46])^(a[156] & b[47])^(a[155] & b[48])^(a[154] & b[49])^(a[153] & b[50])^(a[152] & b[51])^(a[151] & b[52])^(a[150] & b[53])^(a[149] & b[54])^(a[148] & b[55])^(a[147] & b[56])^(a[146] & b[57])^(a[145] & b[58])^(a[144] & b[59])^(a[143] & b[60])^(a[142] & b[61])^(a[141] & b[62])^(a[140] & b[63])^(a[139] & b[64])^(a[138] & b[65])^(a[137] & b[66])^(a[136] & b[67])^(a[135] & b[68])^(a[134] & b[69])^(a[133] & b[70])^(a[132] & b[71])^(a[131] & b[72])^(a[130] & b[73])^(a[129] & b[74])^(a[128] & b[75])^(a[127] & b[76])^(a[126] & b[77])^(a[125] & b[78])^(a[124] & b[79])^(a[123] & b[80])^(a[122] & b[81])^(a[121] & b[82])^(a[120] & b[83])^(a[119] & b[84])^(a[118] & b[85])^(a[117] & b[86])^(a[116] & b[87])^(a[115] & b[88])^(a[114] & b[89])^(a[113] & b[90])^(a[112] & b[91])^(a[111] & b[92])^(a[110] & b[93])^(a[109] & b[94])^(a[108] & b[95])^(a[107] & b[96])^(a[106] & b[97])^(a[105] & b[98])^(a[104] & b[99])^(a[103] & b[100])^(a[102] & b[101])^(a[101] & b[102])^(a[100] & b[103])^(a[99] & b[104])^(a[98] & b[105])^(a[97] & b[106])^(a[96] & b[107])^(a[95] & b[108])^(a[94] & b[109])^(a[93] & b[110])^(a[92] & b[111])^(a[91] & b[112])^(a[90] & b[113])^(a[89] & b[114])^(a[88] & b[115])^(a[87] & b[116])^(a[86] & b[117])^(a[85] & b[118])^(a[84] & b[119])^(a[83] & b[120])^(a[82] & b[121])^(a[81] & b[122])^(a[80] & b[123])^(a[79] & b[124])^(a[78] & b[125])^(a[77] & b[126])^(a[76] & b[127])^(a[75] & b[128])^(a[74] & b[129])^(a[73] & b[130])^(a[72] & b[131])^(a[71] & b[132])^(a[70] & b[133])^(a[69] & b[134])^(a[68] & b[135])^(a[67] & b[136])^(a[66] & b[137])^(a[65] & b[138])^(a[64] & b[139])^(a[63] & b[140])^(a[62] & b[141])^(a[61] & b[142])^(a[60] & b[143])^(a[59] & b[144])^(a[58] & b[145])^(a[57] & b[146])^(a[56] & b[147])^(a[55] & b[148])^(a[54] & b[149])^(a[53] & b[150])^(a[52] & b[151])^(a[51] & b[152])^(a[50] & b[153])^(a[49] & b[154])^(a[48] & b[155])^(a[47] & b[156])^(a[46] & b[157])^(a[45] & b[158])^(a[44] & b[159])^(a[43] & b[160])^(a[42] & b[161])^(a[41] & b[162])^(a[40] & b[163])^(a[39] & b[164])^(a[38] & b[165])^(a[37] & b[166])^(a[36] & b[167])^(a[35] & b[168])^(a[34] & b[169])^(a[33] & b[170])^(a[32] & b[171])^(a[31] & b[172])^(a[30] & b[173])^(a[29] & b[174])^(a[28] & b[175])^(a[27] & b[176])^(a[26] & b[177])^(a[25] & b[178])^(a[24] & b[179])^(a[23] & b[180])^(a[22] & b[181])^(a[21] & b[182])^(a[20] & b[183])^(a[19] & b[184])^(a[18] & b[185])^(a[17] & b[186])^(a[16] & b[187])^(a[15] & b[188])^(a[14] & b[189])^(a[13] & b[190])^(a[12] & b[191])^(a[11] & b[192])^(a[10] & b[193])^(a[9] & b[194])^(a[8] & b[195])^(a[7] & b[196])^(a[6] & b[197])^(a[5] & b[198])^(a[4] & b[199])^(a[3] & b[200])^(a[2] & b[201])^(a[1] & b[202])^(a[0] & b[203]);
assign y[204] = (a[204] & b[0])^(a[203] & b[1])^(a[202] & b[2])^(a[201] & b[3])^(a[200] & b[4])^(a[199] & b[5])^(a[198] & b[6])^(a[197] & b[7])^(a[196] & b[8])^(a[195] & b[9])^(a[194] & b[10])^(a[193] & b[11])^(a[192] & b[12])^(a[191] & b[13])^(a[190] & b[14])^(a[189] & b[15])^(a[188] & b[16])^(a[187] & b[17])^(a[186] & b[18])^(a[185] & b[19])^(a[184] & b[20])^(a[183] & b[21])^(a[182] & b[22])^(a[181] & b[23])^(a[180] & b[24])^(a[179] & b[25])^(a[178] & b[26])^(a[177] & b[27])^(a[176] & b[28])^(a[175] & b[29])^(a[174] & b[30])^(a[173] & b[31])^(a[172] & b[32])^(a[171] & b[33])^(a[170] & b[34])^(a[169] & b[35])^(a[168] & b[36])^(a[167] & b[37])^(a[166] & b[38])^(a[165] & b[39])^(a[164] & b[40])^(a[163] & b[41])^(a[162] & b[42])^(a[161] & b[43])^(a[160] & b[44])^(a[159] & b[45])^(a[158] & b[46])^(a[157] & b[47])^(a[156] & b[48])^(a[155] & b[49])^(a[154] & b[50])^(a[153] & b[51])^(a[152] & b[52])^(a[151] & b[53])^(a[150] & b[54])^(a[149] & b[55])^(a[148] & b[56])^(a[147] & b[57])^(a[146] & b[58])^(a[145] & b[59])^(a[144] & b[60])^(a[143] & b[61])^(a[142] & b[62])^(a[141] & b[63])^(a[140] & b[64])^(a[139] & b[65])^(a[138] & b[66])^(a[137] & b[67])^(a[136] & b[68])^(a[135] & b[69])^(a[134] & b[70])^(a[133] & b[71])^(a[132] & b[72])^(a[131] & b[73])^(a[130] & b[74])^(a[129] & b[75])^(a[128] & b[76])^(a[127] & b[77])^(a[126] & b[78])^(a[125] & b[79])^(a[124] & b[80])^(a[123] & b[81])^(a[122] & b[82])^(a[121] & b[83])^(a[120] & b[84])^(a[119] & b[85])^(a[118] & b[86])^(a[117] & b[87])^(a[116] & b[88])^(a[115] & b[89])^(a[114] & b[90])^(a[113] & b[91])^(a[112] & b[92])^(a[111] & b[93])^(a[110] & b[94])^(a[109] & b[95])^(a[108] & b[96])^(a[107] & b[97])^(a[106] & b[98])^(a[105] & b[99])^(a[104] & b[100])^(a[103] & b[101])^(a[102] & b[102])^(a[101] & b[103])^(a[100] & b[104])^(a[99] & b[105])^(a[98] & b[106])^(a[97] & b[107])^(a[96] & b[108])^(a[95] & b[109])^(a[94] & b[110])^(a[93] & b[111])^(a[92] & b[112])^(a[91] & b[113])^(a[90] & b[114])^(a[89] & b[115])^(a[88] & b[116])^(a[87] & b[117])^(a[86] & b[118])^(a[85] & b[119])^(a[84] & b[120])^(a[83] & b[121])^(a[82] & b[122])^(a[81] & b[123])^(a[80] & b[124])^(a[79] & b[125])^(a[78] & b[126])^(a[77] & b[127])^(a[76] & b[128])^(a[75] & b[129])^(a[74] & b[130])^(a[73] & b[131])^(a[72] & b[132])^(a[71] & b[133])^(a[70] & b[134])^(a[69] & b[135])^(a[68] & b[136])^(a[67] & b[137])^(a[66] & b[138])^(a[65] & b[139])^(a[64] & b[140])^(a[63] & b[141])^(a[62] & b[142])^(a[61] & b[143])^(a[60] & b[144])^(a[59] & b[145])^(a[58] & b[146])^(a[57] & b[147])^(a[56] & b[148])^(a[55] & b[149])^(a[54] & b[150])^(a[53] & b[151])^(a[52] & b[152])^(a[51] & b[153])^(a[50] & b[154])^(a[49] & b[155])^(a[48] & b[156])^(a[47] & b[157])^(a[46] & b[158])^(a[45] & b[159])^(a[44] & b[160])^(a[43] & b[161])^(a[42] & b[162])^(a[41] & b[163])^(a[40] & b[164])^(a[39] & b[165])^(a[38] & b[166])^(a[37] & b[167])^(a[36] & b[168])^(a[35] & b[169])^(a[34] & b[170])^(a[33] & b[171])^(a[32] & b[172])^(a[31] & b[173])^(a[30] & b[174])^(a[29] & b[175])^(a[28] & b[176])^(a[27] & b[177])^(a[26] & b[178])^(a[25] & b[179])^(a[24] & b[180])^(a[23] & b[181])^(a[22] & b[182])^(a[21] & b[183])^(a[20] & b[184])^(a[19] & b[185])^(a[18] & b[186])^(a[17] & b[187])^(a[16] & b[188])^(a[15] & b[189])^(a[14] & b[190])^(a[13] & b[191])^(a[12] & b[192])^(a[11] & b[193])^(a[10] & b[194])^(a[9] & b[195])^(a[8] & b[196])^(a[7] & b[197])^(a[6] & b[198])^(a[5] & b[199])^(a[4] & b[200])^(a[3] & b[201])^(a[2] & b[202])^(a[1] & b[203])^(a[0] & b[204]);
assign y[205] = (a[205] & b[0])^(a[204] & b[1])^(a[203] & b[2])^(a[202] & b[3])^(a[201] & b[4])^(a[200] & b[5])^(a[199] & b[6])^(a[198] & b[7])^(a[197] & b[8])^(a[196] & b[9])^(a[195] & b[10])^(a[194] & b[11])^(a[193] & b[12])^(a[192] & b[13])^(a[191] & b[14])^(a[190] & b[15])^(a[189] & b[16])^(a[188] & b[17])^(a[187] & b[18])^(a[186] & b[19])^(a[185] & b[20])^(a[184] & b[21])^(a[183] & b[22])^(a[182] & b[23])^(a[181] & b[24])^(a[180] & b[25])^(a[179] & b[26])^(a[178] & b[27])^(a[177] & b[28])^(a[176] & b[29])^(a[175] & b[30])^(a[174] & b[31])^(a[173] & b[32])^(a[172] & b[33])^(a[171] & b[34])^(a[170] & b[35])^(a[169] & b[36])^(a[168] & b[37])^(a[167] & b[38])^(a[166] & b[39])^(a[165] & b[40])^(a[164] & b[41])^(a[163] & b[42])^(a[162] & b[43])^(a[161] & b[44])^(a[160] & b[45])^(a[159] & b[46])^(a[158] & b[47])^(a[157] & b[48])^(a[156] & b[49])^(a[155] & b[50])^(a[154] & b[51])^(a[153] & b[52])^(a[152] & b[53])^(a[151] & b[54])^(a[150] & b[55])^(a[149] & b[56])^(a[148] & b[57])^(a[147] & b[58])^(a[146] & b[59])^(a[145] & b[60])^(a[144] & b[61])^(a[143] & b[62])^(a[142] & b[63])^(a[141] & b[64])^(a[140] & b[65])^(a[139] & b[66])^(a[138] & b[67])^(a[137] & b[68])^(a[136] & b[69])^(a[135] & b[70])^(a[134] & b[71])^(a[133] & b[72])^(a[132] & b[73])^(a[131] & b[74])^(a[130] & b[75])^(a[129] & b[76])^(a[128] & b[77])^(a[127] & b[78])^(a[126] & b[79])^(a[125] & b[80])^(a[124] & b[81])^(a[123] & b[82])^(a[122] & b[83])^(a[121] & b[84])^(a[120] & b[85])^(a[119] & b[86])^(a[118] & b[87])^(a[117] & b[88])^(a[116] & b[89])^(a[115] & b[90])^(a[114] & b[91])^(a[113] & b[92])^(a[112] & b[93])^(a[111] & b[94])^(a[110] & b[95])^(a[109] & b[96])^(a[108] & b[97])^(a[107] & b[98])^(a[106] & b[99])^(a[105] & b[100])^(a[104] & b[101])^(a[103] & b[102])^(a[102] & b[103])^(a[101] & b[104])^(a[100] & b[105])^(a[99] & b[106])^(a[98] & b[107])^(a[97] & b[108])^(a[96] & b[109])^(a[95] & b[110])^(a[94] & b[111])^(a[93] & b[112])^(a[92] & b[113])^(a[91] & b[114])^(a[90] & b[115])^(a[89] & b[116])^(a[88] & b[117])^(a[87] & b[118])^(a[86] & b[119])^(a[85] & b[120])^(a[84] & b[121])^(a[83] & b[122])^(a[82] & b[123])^(a[81] & b[124])^(a[80] & b[125])^(a[79] & b[126])^(a[78] & b[127])^(a[77] & b[128])^(a[76] & b[129])^(a[75] & b[130])^(a[74] & b[131])^(a[73] & b[132])^(a[72] & b[133])^(a[71] & b[134])^(a[70] & b[135])^(a[69] & b[136])^(a[68] & b[137])^(a[67] & b[138])^(a[66] & b[139])^(a[65] & b[140])^(a[64] & b[141])^(a[63] & b[142])^(a[62] & b[143])^(a[61] & b[144])^(a[60] & b[145])^(a[59] & b[146])^(a[58] & b[147])^(a[57] & b[148])^(a[56] & b[149])^(a[55] & b[150])^(a[54] & b[151])^(a[53] & b[152])^(a[52] & b[153])^(a[51] & b[154])^(a[50] & b[155])^(a[49] & b[156])^(a[48] & b[157])^(a[47] & b[158])^(a[46] & b[159])^(a[45] & b[160])^(a[44] & b[161])^(a[43] & b[162])^(a[42] & b[163])^(a[41] & b[164])^(a[40] & b[165])^(a[39] & b[166])^(a[38] & b[167])^(a[37] & b[168])^(a[36] & b[169])^(a[35] & b[170])^(a[34] & b[171])^(a[33] & b[172])^(a[32] & b[173])^(a[31] & b[174])^(a[30] & b[175])^(a[29] & b[176])^(a[28] & b[177])^(a[27] & b[178])^(a[26] & b[179])^(a[25] & b[180])^(a[24] & b[181])^(a[23] & b[182])^(a[22] & b[183])^(a[21] & b[184])^(a[20] & b[185])^(a[19] & b[186])^(a[18] & b[187])^(a[17] & b[188])^(a[16] & b[189])^(a[15] & b[190])^(a[14] & b[191])^(a[13] & b[192])^(a[12] & b[193])^(a[11] & b[194])^(a[10] & b[195])^(a[9] & b[196])^(a[8] & b[197])^(a[7] & b[198])^(a[6] & b[199])^(a[5] & b[200])^(a[4] & b[201])^(a[3] & b[202])^(a[2] & b[203])^(a[1] & b[204])^(a[0] & b[205]);
assign y[206] = (a[206] & b[0])^(a[205] & b[1])^(a[204] & b[2])^(a[203] & b[3])^(a[202] & b[4])^(a[201] & b[5])^(a[200] & b[6])^(a[199] & b[7])^(a[198] & b[8])^(a[197] & b[9])^(a[196] & b[10])^(a[195] & b[11])^(a[194] & b[12])^(a[193] & b[13])^(a[192] & b[14])^(a[191] & b[15])^(a[190] & b[16])^(a[189] & b[17])^(a[188] & b[18])^(a[187] & b[19])^(a[186] & b[20])^(a[185] & b[21])^(a[184] & b[22])^(a[183] & b[23])^(a[182] & b[24])^(a[181] & b[25])^(a[180] & b[26])^(a[179] & b[27])^(a[178] & b[28])^(a[177] & b[29])^(a[176] & b[30])^(a[175] & b[31])^(a[174] & b[32])^(a[173] & b[33])^(a[172] & b[34])^(a[171] & b[35])^(a[170] & b[36])^(a[169] & b[37])^(a[168] & b[38])^(a[167] & b[39])^(a[166] & b[40])^(a[165] & b[41])^(a[164] & b[42])^(a[163] & b[43])^(a[162] & b[44])^(a[161] & b[45])^(a[160] & b[46])^(a[159] & b[47])^(a[158] & b[48])^(a[157] & b[49])^(a[156] & b[50])^(a[155] & b[51])^(a[154] & b[52])^(a[153] & b[53])^(a[152] & b[54])^(a[151] & b[55])^(a[150] & b[56])^(a[149] & b[57])^(a[148] & b[58])^(a[147] & b[59])^(a[146] & b[60])^(a[145] & b[61])^(a[144] & b[62])^(a[143] & b[63])^(a[142] & b[64])^(a[141] & b[65])^(a[140] & b[66])^(a[139] & b[67])^(a[138] & b[68])^(a[137] & b[69])^(a[136] & b[70])^(a[135] & b[71])^(a[134] & b[72])^(a[133] & b[73])^(a[132] & b[74])^(a[131] & b[75])^(a[130] & b[76])^(a[129] & b[77])^(a[128] & b[78])^(a[127] & b[79])^(a[126] & b[80])^(a[125] & b[81])^(a[124] & b[82])^(a[123] & b[83])^(a[122] & b[84])^(a[121] & b[85])^(a[120] & b[86])^(a[119] & b[87])^(a[118] & b[88])^(a[117] & b[89])^(a[116] & b[90])^(a[115] & b[91])^(a[114] & b[92])^(a[113] & b[93])^(a[112] & b[94])^(a[111] & b[95])^(a[110] & b[96])^(a[109] & b[97])^(a[108] & b[98])^(a[107] & b[99])^(a[106] & b[100])^(a[105] & b[101])^(a[104] & b[102])^(a[103] & b[103])^(a[102] & b[104])^(a[101] & b[105])^(a[100] & b[106])^(a[99] & b[107])^(a[98] & b[108])^(a[97] & b[109])^(a[96] & b[110])^(a[95] & b[111])^(a[94] & b[112])^(a[93] & b[113])^(a[92] & b[114])^(a[91] & b[115])^(a[90] & b[116])^(a[89] & b[117])^(a[88] & b[118])^(a[87] & b[119])^(a[86] & b[120])^(a[85] & b[121])^(a[84] & b[122])^(a[83] & b[123])^(a[82] & b[124])^(a[81] & b[125])^(a[80] & b[126])^(a[79] & b[127])^(a[78] & b[128])^(a[77] & b[129])^(a[76] & b[130])^(a[75] & b[131])^(a[74] & b[132])^(a[73] & b[133])^(a[72] & b[134])^(a[71] & b[135])^(a[70] & b[136])^(a[69] & b[137])^(a[68] & b[138])^(a[67] & b[139])^(a[66] & b[140])^(a[65] & b[141])^(a[64] & b[142])^(a[63] & b[143])^(a[62] & b[144])^(a[61] & b[145])^(a[60] & b[146])^(a[59] & b[147])^(a[58] & b[148])^(a[57] & b[149])^(a[56] & b[150])^(a[55] & b[151])^(a[54] & b[152])^(a[53] & b[153])^(a[52] & b[154])^(a[51] & b[155])^(a[50] & b[156])^(a[49] & b[157])^(a[48] & b[158])^(a[47] & b[159])^(a[46] & b[160])^(a[45] & b[161])^(a[44] & b[162])^(a[43] & b[163])^(a[42] & b[164])^(a[41] & b[165])^(a[40] & b[166])^(a[39] & b[167])^(a[38] & b[168])^(a[37] & b[169])^(a[36] & b[170])^(a[35] & b[171])^(a[34] & b[172])^(a[33] & b[173])^(a[32] & b[174])^(a[31] & b[175])^(a[30] & b[176])^(a[29] & b[177])^(a[28] & b[178])^(a[27] & b[179])^(a[26] & b[180])^(a[25] & b[181])^(a[24] & b[182])^(a[23] & b[183])^(a[22] & b[184])^(a[21] & b[185])^(a[20] & b[186])^(a[19] & b[187])^(a[18] & b[188])^(a[17] & b[189])^(a[16] & b[190])^(a[15] & b[191])^(a[14] & b[192])^(a[13] & b[193])^(a[12] & b[194])^(a[11] & b[195])^(a[10] & b[196])^(a[9] & b[197])^(a[8] & b[198])^(a[7] & b[199])^(a[6] & b[200])^(a[5] & b[201])^(a[4] & b[202])^(a[3] & b[203])^(a[2] & b[204])^(a[1] & b[205])^(a[0] & b[206]);
assign y[207] = (a[207] & b[0])^(a[206] & b[1])^(a[205] & b[2])^(a[204] & b[3])^(a[203] & b[4])^(a[202] & b[5])^(a[201] & b[6])^(a[200] & b[7])^(a[199] & b[8])^(a[198] & b[9])^(a[197] & b[10])^(a[196] & b[11])^(a[195] & b[12])^(a[194] & b[13])^(a[193] & b[14])^(a[192] & b[15])^(a[191] & b[16])^(a[190] & b[17])^(a[189] & b[18])^(a[188] & b[19])^(a[187] & b[20])^(a[186] & b[21])^(a[185] & b[22])^(a[184] & b[23])^(a[183] & b[24])^(a[182] & b[25])^(a[181] & b[26])^(a[180] & b[27])^(a[179] & b[28])^(a[178] & b[29])^(a[177] & b[30])^(a[176] & b[31])^(a[175] & b[32])^(a[174] & b[33])^(a[173] & b[34])^(a[172] & b[35])^(a[171] & b[36])^(a[170] & b[37])^(a[169] & b[38])^(a[168] & b[39])^(a[167] & b[40])^(a[166] & b[41])^(a[165] & b[42])^(a[164] & b[43])^(a[163] & b[44])^(a[162] & b[45])^(a[161] & b[46])^(a[160] & b[47])^(a[159] & b[48])^(a[158] & b[49])^(a[157] & b[50])^(a[156] & b[51])^(a[155] & b[52])^(a[154] & b[53])^(a[153] & b[54])^(a[152] & b[55])^(a[151] & b[56])^(a[150] & b[57])^(a[149] & b[58])^(a[148] & b[59])^(a[147] & b[60])^(a[146] & b[61])^(a[145] & b[62])^(a[144] & b[63])^(a[143] & b[64])^(a[142] & b[65])^(a[141] & b[66])^(a[140] & b[67])^(a[139] & b[68])^(a[138] & b[69])^(a[137] & b[70])^(a[136] & b[71])^(a[135] & b[72])^(a[134] & b[73])^(a[133] & b[74])^(a[132] & b[75])^(a[131] & b[76])^(a[130] & b[77])^(a[129] & b[78])^(a[128] & b[79])^(a[127] & b[80])^(a[126] & b[81])^(a[125] & b[82])^(a[124] & b[83])^(a[123] & b[84])^(a[122] & b[85])^(a[121] & b[86])^(a[120] & b[87])^(a[119] & b[88])^(a[118] & b[89])^(a[117] & b[90])^(a[116] & b[91])^(a[115] & b[92])^(a[114] & b[93])^(a[113] & b[94])^(a[112] & b[95])^(a[111] & b[96])^(a[110] & b[97])^(a[109] & b[98])^(a[108] & b[99])^(a[107] & b[100])^(a[106] & b[101])^(a[105] & b[102])^(a[104] & b[103])^(a[103] & b[104])^(a[102] & b[105])^(a[101] & b[106])^(a[100] & b[107])^(a[99] & b[108])^(a[98] & b[109])^(a[97] & b[110])^(a[96] & b[111])^(a[95] & b[112])^(a[94] & b[113])^(a[93] & b[114])^(a[92] & b[115])^(a[91] & b[116])^(a[90] & b[117])^(a[89] & b[118])^(a[88] & b[119])^(a[87] & b[120])^(a[86] & b[121])^(a[85] & b[122])^(a[84] & b[123])^(a[83] & b[124])^(a[82] & b[125])^(a[81] & b[126])^(a[80] & b[127])^(a[79] & b[128])^(a[78] & b[129])^(a[77] & b[130])^(a[76] & b[131])^(a[75] & b[132])^(a[74] & b[133])^(a[73] & b[134])^(a[72] & b[135])^(a[71] & b[136])^(a[70] & b[137])^(a[69] & b[138])^(a[68] & b[139])^(a[67] & b[140])^(a[66] & b[141])^(a[65] & b[142])^(a[64] & b[143])^(a[63] & b[144])^(a[62] & b[145])^(a[61] & b[146])^(a[60] & b[147])^(a[59] & b[148])^(a[58] & b[149])^(a[57] & b[150])^(a[56] & b[151])^(a[55] & b[152])^(a[54] & b[153])^(a[53] & b[154])^(a[52] & b[155])^(a[51] & b[156])^(a[50] & b[157])^(a[49] & b[158])^(a[48] & b[159])^(a[47] & b[160])^(a[46] & b[161])^(a[45] & b[162])^(a[44] & b[163])^(a[43] & b[164])^(a[42] & b[165])^(a[41] & b[166])^(a[40] & b[167])^(a[39] & b[168])^(a[38] & b[169])^(a[37] & b[170])^(a[36] & b[171])^(a[35] & b[172])^(a[34] & b[173])^(a[33] & b[174])^(a[32] & b[175])^(a[31] & b[176])^(a[30] & b[177])^(a[29] & b[178])^(a[28] & b[179])^(a[27] & b[180])^(a[26] & b[181])^(a[25] & b[182])^(a[24] & b[183])^(a[23] & b[184])^(a[22] & b[185])^(a[21] & b[186])^(a[20] & b[187])^(a[19] & b[188])^(a[18] & b[189])^(a[17] & b[190])^(a[16] & b[191])^(a[15] & b[192])^(a[14] & b[193])^(a[13] & b[194])^(a[12] & b[195])^(a[11] & b[196])^(a[10] & b[197])^(a[9] & b[198])^(a[8] & b[199])^(a[7] & b[200])^(a[6] & b[201])^(a[5] & b[202])^(a[4] & b[203])^(a[3] & b[204])^(a[2] & b[205])^(a[1] & b[206])^(a[0] & b[207]);
assign y[208] = (a[208] & b[0])^(a[207] & b[1])^(a[206] & b[2])^(a[205] & b[3])^(a[204] & b[4])^(a[203] & b[5])^(a[202] & b[6])^(a[201] & b[7])^(a[200] & b[8])^(a[199] & b[9])^(a[198] & b[10])^(a[197] & b[11])^(a[196] & b[12])^(a[195] & b[13])^(a[194] & b[14])^(a[193] & b[15])^(a[192] & b[16])^(a[191] & b[17])^(a[190] & b[18])^(a[189] & b[19])^(a[188] & b[20])^(a[187] & b[21])^(a[186] & b[22])^(a[185] & b[23])^(a[184] & b[24])^(a[183] & b[25])^(a[182] & b[26])^(a[181] & b[27])^(a[180] & b[28])^(a[179] & b[29])^(a[178] & b[30])^(a[177] & b[31])^(a[176] & b[32])^(a[175] & b[33])^(a[174] & b[34])^(a[173] & b[35])^(a[172] & b[36])^(a[171] & b[37])^(a[170] & b[38])^(a[169] & b[39])^(a[168] & b[40])^(a[167] & b[41])^(a[166] & b[42])^(a[165] & b[43])^(a[164] & b[44])^(a[163] & b[45])^(a[162] & b[46])^(a[161] & b[47])^(a[160] & b[48])^(a[159] & b[49])^(a[158] & b[50])^(a[157] & b[51])^(a[156] & b[52])^(a[155] & b[53])^(a[154] & b[54])^(a[153] & b[55])^(a[152] & b[56])^(a[151] & b[57])^(a[150] & b[58])^(a[149] & b[59])^(a[148] & b[60])^(a[147] & b[61])^(a[146] & b[62])^(a[145] & b[63])^(a[144] & b[64])^(a[143] & b[65])^(a[142] & b[66])^(a[141] & b[67])^(a[140] & b[68])^(a[139] & b[69])^(a[138] & b[70])^(a[137] & b[71])^(a[136] & b[72])^(a[135] & b[73])^(a[134] & b[74])^(a[133] & b[75])^(a[132] & b[76])^(a[131] & b[77])^(a[130] & b[78])^(a[129] & b[79])^(a[128] & b[80])^(a[127] & b[81])^(a[126] & b[82])^(a[125] & b[83])^(a[124] & b[84])^(a[123] & b[85])^(a[122] & b[86])^(a[121] & b[87])^(a[120] & b[88])^(a[119] & b[89])^(a[118] & b[90])^(a[117] & b[91])^(a[116] & b[92])^(a[115] & b[93])^(a[114] & b[94])^(a[113] & b[95])^(a[112] & b[96])^(a[111] & b[97])^(a[110] & b[98])^(a[109] & b[99])^(a[108] & b[100])^(a[107] & b[101])^(a[106] & b[102])^(a[105] & b[103])^(a[104] & b[104])^(a[103] & b[105])^(a[102] & b[106])^(a[101] & b[107])^(a[100] & b[108])^(a[99] & b[109])^(a[98] & b[110])^(a[97] & b[111])^(a[96] & b[112])^(a[95] & b[113])^(a[94] & b[114])^(a[93] & b[115])^(a[92] & b[116])^(a[91] & b[117])^(a[90] & b[118])^(a[89] & b[119])^(a[88] & b[120])^(a[87] & b[121])^(a[86] & b[122])^(a[85] & b[123])^(a[84] & b[124])^(a[83] & b[125])^(a[82] & b[126])^(a[81] & b[127])^(a[80] & b[128])^(a[79] & b[129])^(a[78] & b[130])^(a[77] & b[131])^(a[76] & b[132])^(a[75] & b[133])^(a[74] & b[134])^(a[73] & b[135])^(a[72] & b[136])^(a[71] & b[137])^(a[70] & b[138])^(a[69] & b[139])^(a[68] & b[140])^(a[67] & b[141])^(a[66] & b[142])^(a[65] & b[143])^(a[64] & b[144])^(a[63] & b[145])^(a[62] & b[146])^(a[61] & b[147])^(a[60] & b[148])^(a[59] & b[149])^(a[58] & b[150])^(a[57] & b[151])^(a[56] & b[152])^(a[55] & b[153])^(a[54] & b[154])^(a[53] & b[155])^(a[52] & b[156])^(a[51] & b[157])^(a[50] & b[158])^(a[49] & b[159])^(a[48] & b[160])^(a[47] & b[161])^(a[46] & b[162])^(a[45] & b[163])^(a[44] & b[164])^(a[43] & b[165])^(a[42] & b[166])^(a[41] & b[167])^(a[40] & b[168])^(a[39] & b[169])^(a[38] & b[170])^(a[37] & b[171])^(a[36] & b[172])^(a[35] & b[173])^(a[34] & b[174])^(a[33] & b[175])^(a[32] & b[176])^(a[31] & b[177])^(a[30] & b[178])^(a[29] & b[179])^(a[28] & b[180])^(a[27] & b[181])^(a[26] & b[182])^(a[25] & b[183])^(a[24] & b[184])^(a[23] & b[185])^(a[22] & b[186])^(a[21] & b[187])^(a[20] & b[188])^(a[19] & b[189])^(a[18] & b[190])^(a[17] & b[191])^(a[16] & b[192])^(a[15] & b[193])^(a[14] & b[194])^(a[13] & b[195])^(a[12] & b[196])^(a[11] & b[197])^(a[10] & b[198])^(a[9] & b[199])^(a[8] & b[200])^(a[7] & b[201])^(a[6] & b[202])^(a[5] & b[203])^(a[4] & b[204])^(a[3] & b[205])^(a[2] & b[206])^(a[1] & b[207])^(a[0] & b[208]);
assign y[209] = (a[209] & b[0])^(a[208] & b[1])^(a[207] & b[2])^(a[206] & b[3])^(a[205] & b[4])^(a[204] & b[5])^(a[203] & b[6])^(a[202] & b[7])^(a[201] & b[8])^(a[200] & b[9])^(a[199] & b[10])^(a[198] & b[11])^(a[197] & b[12])^(a[196] & b[13])^(a[195] & b[14])^(a[194] & b[15])^(a[193] & b[16])^(a[192] & b[17])^(a[191] & b[18])^(a[190] & b[19])^(a[189] & b[20])^(a[188] & b[21])^(a[187] & b[22])^(a[186] & b[23])^(a[185] & b[24])^(a[184] & b[25])^(a[183] & b[26])^(a[182] & b[27])^(a[181] & b[28])^(a[180] & b[29])^(a[179] & b[30])^(a[178] & b[31])^(a[177] & b[32])^(a[176] & b[33])^(a[175] & b[34])^(a[174] & b[35])^(a[173] & b[36])^(a[172] & b[37])^(a[171] & b[38])^(a[170] & b[39])^(a[169] & b[40])^(a[168] & b[41])^(a[167] & b[42])^(a[166] & b[43])^(a[165] & b[44])^(a[164] & b[45])^(a[163] & b[46])^(a[162] & b[47])^(a[161] & b[48])^(a[160] & b[49])^(a[159] & b[50])^(a[158] & b[51])^(a[157] & b[52])^(a[156] & b[53])^(a[155] & b[54])^(a[154] & b[55])^(a[153] & b[56])^(a[152] & b[57])^(a[151] & b[58])^(a[150] & b[59])^(a[149] & b[60])^(a[148] & b[61])^(a[147] & b[62])^(a[146] & b[63])^(a[145] & b[64])^(a[144] & b[65])^(a[143] & b[66])^(a[142] & b[67])^(a[141] & b[68])^(a[140] & b[69])^(a[139] & b[70])^(a[138] & b[71])^(a[137] & b[72])^(a[136] & b[73])^(a[135] & b[74])^(a[134] & b[75])^(a[133] & b[76])^(a[132] & b[77])^(a[131] & b[78])^(a[130] & b[79])^(a[129] & b[80])^(a[128] & b[81])^(a[127] & b[82])^(a[126] & b[83])^(a[125] & b[84])^(a[124] & b[85])^(a[123] & b[86])^(a[122] & b[87])^(a[121] & b[88])^(a[120] & b[89])^(a[119] & b[90])^(a[118] & b[91])^(a[117] & b[92])^(a[116] & b[93])^(a[115] & b[94])^(a[114] & b[95])^(a[113] & b[96])^(a[112] & b[97])^(a[111] & b[98])^(a[110] & b[99])^(a[109] & b[100])^(a[108] & b[101])^(a[107] & b[102])^(a[106] & b[103])^(a[105] & b[104])^(a[104] & b[105])^(a[103] & b[106])^(a[102] & b[107])^(a[101] & b[108])^(a[100] & b[109])^(a[99] & b[110])^(a[98] & b[111])^(a[97] & b[112])^(a[96] & b[113])^(a[95] & b[114])^(a[94] & b[115])^(a[93] & b[116])^(a[92] & b[117])^(a[91] & b[118])^(a[90] & b[119])^(a[89] & b[120])^(a[88] & b[121])^(a[87] & b[122])^(a[86] & b[123])^(a[85] & b[124])^(a[84] & b[125])^(a[83] & b[126])^(a[82] & b[127])^(a[81] & b[128])^(a[80] & b[129])^(a[79] & b[130])^(a[78] & b[131])^(a[77] & b[132])^(a[76] & b[133])^(a[75] & b[134])^(a[74] & b[135])^(a[73] & b[136])^(a[72] & b[137])^(a[71] & b[138])^(a[70] & b[139])^(a[69] & b[140])^(a[68] & b[141])^(a[67] & b[142])^(a[66] & b[143])^(a[65] & b[144])^(a[64] & b[145])^(a[63] & b[146])^(a[62] & b[147])^(a[61] & b[148])^(a[60] & b[149])^(a[59] & b[150])^(a[58] & b[151])^(a[57] & b[152])^(a[56] & b[153])^(a[55] & b[154])^(a[54] & b[155])^(a[53] & b[156])^(a[52] & b[157])^(a[51] & b[158])^(a[50] & b[159])^(a[49] & b[160])^(a[48] & b[161])^(a[47] & b[162])^(a[46] & b[163])^(a[45] & b[164])^(a[44] & b[165])^(a[43] & b[166])^(a[42] & b[167])^(a[41] & b[168])^(a[40] & b[169])^(a[39] & b[170])^(a[38] & b[171])^(a[37] & b[172])^(a[36] & b[173])^(a[35] & b[174])^(a[34] & b[175])^(a[33] & b[176])^(a[32] & b[177])^(a[31] & b[178])^(a[30] & b[179])^(a[29] & b[180])^(a[28] & b[181])^(a[27] & b[182])^(a[26] & b[183])^(a[25] & b[184])^(a[24] & b[185])^(a[23] & b[186])^(a[22] & b[187])^(a[21] & b[188])^(a[20] & b[189])^(a[19] & b[190])^(a[18] & b[191])^(a[17] & b[192])^(a[16] & b[193])^(a[15] & b[194])^(a[14] & b[195])^(a[13] & b[196])^(a[12] & b[197])^(a[11] & b[198])^(a[10] & b[199])^(a[9] & b[200])^(a[8] & b[201])^(a[7] & b[202])^(a[6] & b[203])^(a[5] & b[204])^(a[4] & b[205])^(a[3] & b[206])^(a[2] & b[207])^(a[1] & b[208])^(a[0] & b[209]);
assign y[210] = (a[210] & b[0])^(a[209] & b[1])^(a[208] & b[2])^(a[207] & b[3])^(a[206] & b[4])^(a[205] & b[5])^(a[204] & b[6])^(a[203] & b[7])^(a[202] & b[8])^(a[201] & b[9])^(a[200] & b[10])^(a[199] & b[11])^(a[198] & b[12])^(a[197] & b[13])^(a[196] & b[14])^(a[195] & b[15])^(a[194] & b[16])^(a[193] & b[17])^(a[192] & b[18])^(a[191] & b[19])^(a[190] & b[20])^(a[189] & b[21])^(a[188] & b[22])^(a[187] & b[23])^(a[186] & b[24])^(a[185] & b[25])^(a[184] & b[26])^(a[183] & b[27])^(a[182] & b[28])^(a[181] & b[29])^(a[180] & b[30])^(a[179] & b[31])^(a[178] & b[32])^(a[177] & b[33])^(a[176] & b[34])^(a[175] & b[35])^(a[174] & b[36])^(a[173] & b[37])^(a[172] & b[38])^(a[171] & b[39])^(a[170] & b[40])^(a[169] & b[41])^(a[168] & b[42])^(a[167] & b[43])^(a[166] & b[44])^(a[165] & b[45])^(a[164] & b[46])^(a[163] & b[47])^(a[162] & b[48])^(a[161] & b[49])^(a[160] & b[50])^(a[159] & b[51])^(a[158] & b[52])^(a[157] & b[53])^(a[156] & b[54])^(a[155] & b[55])^(a[154] & b[56])^(a[153] & b[57])^(a[152] & b[58])^(a[151] & b[59])^(a[150] & b[60])^(a[149] & b[61])^(a[148] & b[62])^(a[147] & b[63])^(a[146] & b[64])^(a[145] & b[65])^(a[144] & b[66])^(a[143] & b[67])^(a[142] & b[68])^(a[141] & b[69])^(a[140] & b[70])^(a[139] & b[71])^(a[138] & b[72])^(a[137] & b[73])^(a[136] & b[74])^(a[135] & b[75])^(a[134] & b[76])^(a[133] & b[77])^(a[132] & b[78])^(a[131] & b[79])^(a[130] & b[80])^(a[129] & b[81])^(a[128] & b[82])^(a[127] & b[83])^(a[126] & b[84])^(a[125] & b[85])^(a[124] & b[86])^(a[123] & b[87])^(a[122] & b[88])^(a[121] & b[89])^(a[120] & b[90])^(a[119] & b[91])^(a[118] & b[92])^(a[117] & b[93])^(a[116] & b[94])^(a[115] & b[95])^(a[114] & b[96])^(a[113] & b[97])^(a[112] & b[98])^(a[111] & b[99])^(a[110] & b[100])^(a[109] & b[101])^(a[108] & b[102])^(a[107] & b[103])^(a[106] & b[104])^(a[105] & b[105])^(a[104] & b[106])^(a[103] & b[107])^(a[102] & b[108])^(a[101] & b[109])^(a[100] & b[110])^(a[99] & b[111])^(a[98] & b[112])^(a[97] & b[113])^(a[96] & b[114])^(a[95] & b[115])^(a[94] & b[116])^(a[93] & b[117])^(a[92] & b[118])^(a[91] & b[119])^(a[90] & b[120])^(a[89] & b[121])^(a[88] & b[122])^(a[87] & b[123])^(a[86] & b[124])^(a[85] & b[125])^(a[84] & b[126])^(a[83] & b[127])^(a[82] & b[128])^(a[81] & b[129])^(a[80] & b[130])^(a[79] & b[131])^(a[78] & b[132])^(a[77] & b[133])^(a[76] & b[134])^(a[75] & b[135])^(a[74] & b[136])^(a[73] & b[137])^(a[72] & b[138])^(a[71] & b[139])^(a[70] & b[140])^(a[69] & b[141])^(a[68] & b[142])^(a[67] & b[143])^(a[66] & b[144])^(a[65] & b[145])^(a[64] & b[146])^(a[63] & b[147])^(a[62] & b[148])^(a[61] & b[149])^(a[60] & b[150])^(a[59] & b[151])^(a[58] & b[152])^(a[57] & b[153])^(a[56] & b[154])^(a[55] & b[155])^(a[54] & b[156])^(a[53] & b[157])^(a[52] & b[158])^(a[51] & b[159])^(a[50] & b[160])^(a[49] & b[161])^(a[48] & b[162])^(a[47] & b[163])^(a[46] & b[164])^(a[45] & b[165])^(a[44] & b[166])^(a[43] & b[167])^(a[42] & b[168])^(a[41] & b[169])^(a[40] & b[170])^(a[39] & b[171])^(a[38] & b[172])^(a[37] & b[173])^(a[36] & b[174])^(a[35] & b[175])^(a[34] & b[176])^(a[33] & b[177])^(a[32] & b[178])^(a[31] & b[179])^(a[30] & b[180])^(a[29] & b[181])^(a[28] & b[182])^(a[27] & b[183])^(a[26] & b[184])^(a[25] & b[185])^(a[24] & b[186])^(a[23] & b[187])^(a[22] & b[188])^(a[21] & b[189])^(a[20] & b[190])^(a[19] & b[191])^(a[18] & b[192])^(a[17] & b[193])^(a[16] & b[194])^(a[15] & b[195])^(a[14] & b[196])^(a[13] & b[197])^(a[12] & b[198])^(a[11] & b[199])^(a[10] & b[200])^(a[9] & b[201])^(a[8] & b[202])^(a[7] & b[203])^(a[6] & b[204])^(a[5] & b[205])^(a[4] & b[206])^(a[3] & b[207])^(a[2] & b[208])^(a[1] & b[209])^(a[0] & b[210]);
assign y[211] = (a[211] & b[0])^(a[210] & b[1])^(a[209] & b[2])^(a[208] & b[3])^(a[207] & b[4])^(a[206] & b[5])^(a[205] & b[6])^(a[204] & b[7])^(a[203] & b[8])^(a[202] & b[9])^(a[201] & b[10])^(a[200] & b[11])^(a[199] & b[12])^(a[198] & b[13])^(a[197] & b[14])^(a[196] & b[15])^(a[195] & b[16])^(a[194] & b[17])^(a[193] & b[18])^(a[192] & b[19])^(a[191] & b[20])^(a[190] & b[21])^(a[189] & b[22])^(a[188] & b[23])^(a[187] & b[24])^(a[186] & b[25])^(a[185] & b[26])^(a[184] & b[27])^(a[183] & b[28])^(a[182] & b[29])^(a[181] & b[30])^(a[180] & b[31])^(a[179] & b[32])^(a[178] & b[33])^(a[177] & b[34])^(a[176] & b[35])^(a[175] & b[36])^(a[174] & b[37])^(a[173] & b[38])^(a[172] & b[39])^(a[171] & b[40])^(a[170] & b[41])^(a[169] & b[42])^(a[168] & b[43])^(a[167] & b[44])^(a[166] & b[45])^(a[165] & b[46])^(a[164] & b[47])^(a[163] & b[48])^(a[162] & b[49])^(a[161] & b[50])^(a[160] & b[51])^(a[159] & b[52])^(a[158] & b[53])^(a[157] & b[54])^(a[156] & b[55])^(a[155] & b[56])^(a[154] & b[57])^(a[153] & b[58])^(a[152] & b[59])^(a[151] & b[60])^(a[150] & b[61])^(a[149] & b[62])^(a[148] & b[63])^(a[147] & b[64])^(a[146] & b[65])^(a[145] & b[66])^(a[144] & b[67])^(a[143] & b[68])^(a[142] & b[69])^(a[141] & b[70])^(a[140] & b[71])^(a[139] & b[72])^(a[138] & b[73])^(a[137] & b[74])^(a[136] & b[75])^(a[135] & b[76])^(a[134] & b[77])^(a[133] & b[78])^(a[132] & b[79])^(a[131] & b[80])^(a[130] & b[81])^(a[129] & b[82])^(a[128] & b[83])^(a[127] & b[84])^(a[126] & b[85])^(a[125] & b[86])^(a[124] & b[87])^(a[123] & b[88])^(a[122] & b[89])^(a[121] & b[90])^(a[120] & b[91])^(a[119] & b[92])^(a[118] & b[93])^(a[117] & b[94])^(a[116] & b[95])^(a[115] & b[96])^(a[114] & b[97])^(a[113] & b[98])^(a[112] & b[99])^(a[111] & b[100])^(a[110] & b[101])^(a[109] & b[102])^(a[108] & b[103])^(a[107] & b[104])^(a[106] & b[105])^(a[105] & b[106])^(a[104] & b[107])^(a[103] & b[108])^(a[102] & b[109])^(a[101] & b[110])^(a[100] & b[111])^(a[99] & b[112])^(a[98] & b[113])^(a[97] & b[114])^(a[96] & b[115])^(a[95] & b[116])^(a[94] & b[117])^(a[93] & b[118])^(a[92] & b[119])^(a[91] & b[120])^(a[90] & b[121])^(a[89] & b[122])^(a[88] & b[123])^(a[87] & b[124])^(a[86] & b[125])^(a[85] & b[126])^(a[84] & b[127])^(a[83] & b[128])^(a[82] & b[129])^(a[81] & b[130])^(a[80] & b[131])^(a[79] & b[132])^(a[78] & b[133])^(a[77] & b[134])^(a[76] & b[135])^(a[75] & b[136])^(a[74] & b[137])^(a[73] & b[138])^(a[72] & b[139])^(a[71] & b[140])^(a[70] & b[141])^(a[69] & b[142])^(a[68] & b[143])^(a[67] & b[144])^(a[66] & b[145])^(a[65] & b[146])^(a[64] & b[147])^(a[63] & b[148])^(a[62] & b[149])^(a[61] & b[150])^(a[60] & b[151])^(a[59] & b[152])^(a[58] & b[153])^(a[57] & b[154])^(a[56] & b[155])^(a[55] & b[156])^(a[54] & b[157])^(a[53] & b[158])^(a[52] & b[159])^(a[51] & b[160])^(a[50] & b[161])^(a[49] & b[162])^(a[48] & b[163])^(a[47] & b[164])^(a[46] & b[165])^(a[45] & b[166])^(a[44] & b[167])^(a[43] & b[168])^(a[42] & b[169])^(a[41] & b[170])^(a[40] & b[171])^(a[39] & b[172])^(a[38] & b[173])^(a[37] & b[174])^(a[36] & b[175])^(a[35] & b[176])^(a[34] & b[177])^(a[33] & b[178])^(a[32] & b[179])^(a[31] & b[180])^(a[30] & b[181])^(a[29] & b[182])^(a[28] & b[183])^(a[27] & b[184])^(a[26] & b[185])^(a[25] & b[186])^(a[24] & b[187])^(a[23] & b[188])^(a[22] & b[189])^(a[21] & b[190])^(a[20] & b[191])^(a[19] & b[192])^(a[18] & b[193])^(a[17] & b[194])^(a[16] & b[195])^(a[15] & b[196])^(a[14] & b[197])^(a[13] & b[198])^(a[12] & b[199])^(a[11] & b[200])^(a[10] & b[201])^(a[9] & b[202])^(a[8] & b[203])^(a[7] & b[204])^(a[6] & b[205])^(a[5] & b[206])^(a[4] & b[207])^(a[3] & b[208])^(a[2] & b[209])^(a[1] & b[210])^(a[0] & b[211]);
assign y[212] = (a[212] & b[0])^(a[211] & b[1])^(a[210] & b[2])^(a[209] & b[3])^(a[208] & b[4])^(a[207] & b[5])^(a[206] & b[6])^(a[205] & b[7])^(a[204] & b[8])^(a[203] & b[9])^(a[202] & b[10])^(a[201] & b[11])^(a[200] & b[12])^(a[199] & b[13])^(a[198] & b[14])^(a[197] & b[15])^(a[196] & b[16])^(a[195] & b[17])^(a[194] & b[18])^(a[193] & b[19])^(a[192] & b[20])^(a[191] & b[21])^(a[190] & b[22])^(a[189] & b[23])^(a[188] & b[24])^(a[187] & b[25])^(a[186] & b[26])^(a[185] & b[27])^(a[184] & b[28])^(a[183] & b[29])^(a[182] & b[30])^(a[181] & b[31])^(a[180] & b[32])^(a[179] & b[33])^(a[178] & b[34])^(a[177] & b[35])^(a[176] & b[36])^(a[175] & b[37])^(a[174] & b[38])^(a[173] & b[39])^(a[172] & b[40])^(a[171] & b[41])^(a[170] & b[42])^(a[169] & b[43])^(a[168] & b[44])^(a[167] & b[45])^(a[166] & b[46])^(a[165] & b[47])^(a[164] & b[48])^(a[163] & b[49])^(a[162] & b[50])^(a[161] & b[51])^(a[160] & b[52])^(a[159] & b[53])^(a[158] & b[54])^(a[157] & b[55])^(a[156] & b[56])^(a[155] & b[57])^(a[154] & b[58])^(a[153] & b[59])^(a[152] & b[60])^(a[151] & b[61])^(a[150] & b[62])^(a[149] & b[63])^(a[148] & b[64])^(a[147] & b[65])^(a[146] & b[66])^(a[145] & b[67])^(a[144] & b[68])^(a[143] & b[69])^(a[142] & b[70])^(a[141] & b[71])^(a[140] & b[72])^(a[139] & b[73])^(a[138] & b[74])^(a[137] & b[75])^(a[136] & b[76])^(a[135] & b[77])^(a[134] & b[78])^(a[133] & b[79])^(a[132] & b[80])^(a[131] & b[81])^(a[130] & b[82])^(a[129] & b[83])^(a[128] & b[84])^(a[127] & b[85])^(a[126] & b[86])^(a[125] & b[87])^(a[124] & b[88])^(a[123] & b[89])^(a[122] & b[90])^(a[121] & b[91])^(a[120] & b[92])^(a[119] & b[93])^(a[118] & b[94])^(a[117] & b[95])^(a[116] & b[96])^(a[115] & b[97])^(a[114] & b[98])^(a[113] & b[99])^(a[112] & b[100])^(a[111] & b[101])^(a[110] & b[102])^(a[109] & b[103])^(a[108] & b[104])^(a[107] & b[105])^(a[106] & b[106])^(a[105] & b[107])^(a[104] & b[108])^(a[103] & b[109])^(a[102] & b[110])^(a[101] & b[111])^(a[100] & b[112])^(a[99] & b[113])^(a[98] & b[114])^(a[97] & b[115])^(a[96] & b[116])^(a[95] & b[117])^(a[94] & b[118])^(a[93] & b[119])^(a[92] & b[120])^(a[91] & b[121])^(a[90] & b[122])^(a[89] & b[123])^(a[88] & b[124])^(a[87] & b[125])^(a[86] & b[126])^(a[85] & b[127])^(a[84] & b[128])^(a[83] & b[129])^(a[82] & b[130])^(a[81] & b[131])^(a[80] & b[132])^(a[79] & b[133])^(a[78] & b[134])^(a[77] & b[135])^(a[76] & b[136])^(a[75] & b[137])^(a[74] & b[138])^(a[73] & b[139])^(a[72] & b[140])^(a[71] & b[141])^(a[70] & b[142])^(a[69] & b[143])^(a[68] & b[144])^(a[67] & b[145])^(a[66] & b[146])^(a[65] & b[147])^(a[64] & b[148])^(a[63] & b[149])^(a[62] & b[150])^(a[61] & b[151])^(a[60] & b[152])^(a[59] & b[153])^(a[58] & b[154])^(a[57] & b[155])^(a[56] & b[156])^(a[55] & b[157])^(a[54] & b[158])^(a[53] & b[159])^(a[52] & b[160])^(a[51] & b[161])^(a[50] & b[162])^(a[49] & b[163])^(a[48] & b[164])^(a[47] & b[165])^(a[46] & b[166])^(a[45] & b[167])^(a[44] & b[168])^(a[43] & b[169])^(a[42] & b[170])^(a[41] & b[171])^(a[40] & b[172])^(a[39] & b[173])^(a[38] & b[174])^(a[37] & b[175])^(a[36] & b[176])^(a[35] & b[177])^(a[34] & b[178])^(a[33] & b[179])^(a[32] & b[180])^(a[31] & b[181])^(a[30] & b[182])^(a[29] & b[183])^(a[28] & b[184])^(a[27] & b[185])^(a[26] & b[186])^(a[25] & b[187])^(a[24] & b[188])^(a[23] & b[189])^(a[22] & b[190])^(a[21] & b[191])^(a[20] & b[192])^(a[19] & b[193])^(a[18] & b[194])^(a[17] & b[195])^(a[16] & b[196])^(a[15] & b[197])^(a[14] & b[198])^(a[13] & b[199])^(a[12] & b[200])^(a[11] & b[201])^(a[10] & b[202])^(a[9] & b[203])^(a[8] & b[204])^(a[7] & b[205])^(a[6] & b[206])^(a[5] & b[207])^(a[4] & b[208])^(a[3] & b[209])^(a[2] & b[210])^(a[1] & b[211])^(a[0] & b[212]);
assign y[213] = (a[213] & b[0])^(a[212] & b[1])^(a[211] & b[2])^(a[210] & b[3])^(a[209] & b[4])^(a[208] & b[5])^(a[207] & b[6])^(a[206] & b[7])^(a[205] & b[8])^(a[204] & b[9])^(a[203] & b[10])^(a[202] & b[11])^(a[201] & b[12])^(a[200] & b[13])^(a[199] & b[14])^(a[198] & b[15])^(a[197] & b[16])^(a[196] & b[17])^(a[195] & b[18])^(a[194] & b[19])^(a[193] & b[20])^(a[192] & b[21])^(a[191] & b[22])^(a[190] & b[23])^(a[189] & b[24])^(a[188] & b[25])^(a[187] & b[26])^(a[186] & b[27])^(a[185] & b[28])^(a[184] & b[29])^(a[183] & b[30])^(a[182] & b[31])^(a[181] & b[32])^(a[180] & b[33])^(a[179] & b[34])^(a[178] & b[35])^(a[177] & b[36])^(a[176] & b[37])^(a[175] & b[38])^(a[174] & b[39])^(a[173] & b[40])^(a[172] & b[41])^(a[171] & b[42])^(a[170] & b[43])^(a[169] & b[44])^(a[168] & b[45])^(a[167] & b[46])^(a[166] & b[47])^(a[165] & b[48])^(a[164] & b[49])^(a[163] & b[50])^(a[162] & b[51])^(a[161] & b[52])^(a[160] & b[53])^(a[159] & b[54])^(a[158] & b[55])^(a[157] & b[56])^(a[156] & b[57])^(a[155] & b[58])^(a[154] & b[59])^(a[153] & b[60])^(a[152] & b[61])^(a[151] & b[62])^(a[150] & b[63])^(a[149] & b[64])^(a[148] & b[65])^(a[147] & b[66])^(a[146] & b[67])^(a[145] & b[68])^(a[144] & b[69])^(a[143] & b[70])^(a[142] & b[71])^(a[141] & b[72])^(a[140] & b[73])^(a[139] & b[74])^(a[138] & b[75])^(a[137] & b[76])^(a[136] & b[77])^(a[135] & b[78])^(a[134] & b[79])^(a[133] & b[80])^(a[132] & b[81])^(a[131] & b[82])^(a[130] & b[83])^(a[129] & b[84])^(a[128] & b[85])^(a[127] & b[86])^(a[126] & b[87])^(a[125] & b[88])^(a[124] & b[89])^(a[123] & b[90])^(a[122] & b[91])^(a[121] & b[92])^(a[120] & b[93])^(a[119] & b[94])^(a[118] & b[95])^(a[117] & b[96])^(a[116] & b[97])^(a[115] & b[98])^(a[114] & b[99])^(a[113] & b[100])^(a[112] & b[101])^(a[111] & b[102])^(a[110] & b[103])^(a[109] & b[104])^(a[108] & b[105])^(a[107] & b[106])^(a[106] & b[107])^(a[105] & b[108])^(a[104] & b[109])^(a[103] & b[110])^(a[102] & b[111])^(a[101] & b[112])^(a[100] & b[113])^(a[99] & b[114])^(a[98] & b[115])^(a[97] & b[116])^(a[96] & b[117])^(a[95] & b[118])^(a[94] & b[119])^(a[93] & b[120])^(a[92] & b[121])^(a[91] & b[122])^(a[90] & b[123])^(a[89] & b[124])^(a[88] & b[125])^(a[87] & b[126])^(a[86] & b[127])^(a[85] & b[128])^(a[84] & b[129])^(a[83] & b[130])^(a[82] & b[131])^(a[81] & b[132])^(a[80] & b[133])^(a[79] & b[134])^(a[78] & b[135])^(a[77] & b[136])^(a[76] & b[137])^(a[75] & b[138])^(a[74] & b[139])^(a[73] & b[140])^(a[72] & b[141])^(a[71] & b[142])^(a[70] & b[143])^(a[69] & b[144])^(a[68] & b[145])^(a[67] & b[146])^(a[66] & b[147])^(a[65] & b[148])^(a[64] & b[149])^(a[63] & b[150])^(a[62] & b[151])^(a[61] & b[152])^(a[60] & b[153])^(a[59] & b[154])^(a[58] & b[155])^(a[57] & b[156])^(a[56] & b[157])^(a[55] & b[158])^(a[54] & b[159])^(a[53] & b[160])^(a[52] & b[161])^(a[51] & b[162])^(a[50] & b[163])^(a[49] & b[164])^(a[48] & b[165])^(a[47] & b[166])^(a[46] & b[167])^(a[45] & b[168])^(a[44] & b[169])^(a[43] & b[170])^(a[42] & b[171])^(a[41] & b[172])^(a[40] & b[173])^(a[39] & b[174])^(a[38] & b[175])^(a[37] & b[176])^(a[36] & b[177])^(a[35] & b[178])^(a[34] & b[179])^(a[33] & b[180])^(a[32] & b[181])^(a[31] & b[182])^(a[30] & b[183])^(a[29] & b[184])^(a[28] & b[185])^(a[27] & b[186])^(a[26] & b[187])^(a[25] & b[188])^(a[24] & b[189])^(a[23] & b[190])^(a[22] & b[191])^(a[21] & b[192])^(a[20] & b[193])^(a[19] & b[194])^(a[18] & b[195])^(a[17] & b[196])^(a[16] & b[197])^(a[15] & b[198])^(a[14] & b[199])^(a[13] & b[200])^(a[12] & b[201])^(a[11] & b[202])^(a[10] & b[203])^(a[9] & b[204])^(a[8] & b[205])^(a[7] & b[206])^(a[6] & b[207])^(a[5] & b[208])^(a[4] & b[209])^(a[3] & b[210])^(a[2] & b[211])^(a[1] & b[212])^(a[0] & b[213]);
assign y[214] = (a[214] & b[0])^(a[213] & b[1])^(a[212] & b[2])^(a[211] & b[3])^(a[210] & b[4])^(a[209] & b[5])^(a[208] & b[6])^(a[207] & b[7])^(a[206] & b[8])^(a[205] & b[9])^(a[204] & b[10])^(a[203] & b[11])^(a[202] & b[12])^(a[201] & b[13])^(a[200] & b[14])^(a[199] & b[15])^(a[198] & b[16])^(a[197] & b[17])^(a[196] & b[18])^(a[195] & b[19])^(a[194] & b[20])^(a[193] & b[21])^(a[192] & b[22])^(a[191] & b[23])^(a[190] & b[24])^(a[189] & b[25])^(a[188] & b[26])^(a[187] & b[27])^(a[186] & b[28])^(a[185] & b[29])^(a[184] & b[30])^(a[183] & b[31])^(a[182] & b[32])^(a[181] & b[33])^(a[180] & b[34])^(a[179] & b[35])^(a[178] & b[36])^(a[177] & b[37])^(a[176] & b[38])^(a[175] & b[39])^(a[174] & b[40])^(a[173] & b[41])^(a[172] & b[42])^(a[171] & b[43])^(a[170] & b[44])^(a[169] & b[45])^(a[168] & b[46])^(a[167] & b[47])^(a[166] & b[48])^(a[165] & b[49])^(a[164] & b[50])^(a[163] & b[51])^(a[162] & b[52])^(a[161] & b[53])^(a[160] & b[54])^(a[159] & b[55])^(a[158] & b[56])^(a[157] & b[57])^(a[156] & b[58])^(a[155] & b[59])^(a[154] & b[60])^(a[153] & b[61])^(a[152] & b[62])^(a[151] & b[63])^(a[150] & b[64])^(a[149] & b[65])^(a[148] & b[66])^(a[147] & b[67])^(a[146] & b[68])^(a[145] & b[69])^(a[144] & b[70])^(a[143] & b[71])^(a[142] & b[72])^(a[141] & b[73])^(a[140] & b[74])^(a[139] & b[75])^(a[138] & b[76])^(a[137] & b[77])^(a[136] & b[78])^(a[135] & b[79])^(a[134] & b[80])^(a[133] & b[81])^(a[132] & b[82])^(a[131] & b[83])^(a[130] & b[84])^(a[129] & b[85])^(a[128] & b[86])^(a[127] & b[87])^(a[126] & b[88])^(a[125] & b[89])^(a[124] & b[90])^(a[123] & b[91])^(a[122] & b[92])^(a[121] & b[93])^(a[120] & b[94])^(a[119] & b[95])^(a[118] & b[96])^(a[117] & b[97])^(a[116] & b[98])^(a[115] & b[99])^(a[114] & b[100])^(a[113] & b[101])^(a[112] & b[102])^(a[111] & b[103])^(a[110] & b[104])^(a[109] & b[105])^(a[108] & b[106])^(a[107] & b[107])^(a[106] & b[108])^(a[105] & b[109])^(a[104] & b[110])^(a[103] & b[111])^(a[102] & b[112])^(a[101] & b[113])^(a[100] & b[114])^(a[99] & b[115])^(a[98] & b[116])^(a[97] & b[117])^(a[96] & b[118])^(a[95] & b[119])^(a[94] & b[120])^(a[93] & b[121])^(a[92] & b[122])^(a[91] & b[123])^(a[90] & b[124])^(a[89] & b[125])^(a[88] & b[126])^(a[87] & b[127])^(a[86] & b[128])^(a[85] & b[129])^(a[84] & b[130])^(a[83] & b[131])^(a[82] & b[132])^(a[81] & b[133])^(a[80] & b[134])^(a[79] & b[135])^(a[78] & b[136])^(a[77] & b[137])^(a[76] & b[138])^(a[75] & b[139])^(a[74] & b[140])^(a[73] & b[141])^(a[72] & b[142])^(a[71] & b[143])^(a[70] & b[144])^(a[69] & b[145])^(a[68] & b[146])^(a[67] & b[147])^(a[66] & b[148])^(a[65] & b[149])^(a[64] & b[150])^(a[63] & b[151])^(a[62] & b[152])^(a[61] & b[153])^(a[60] & b[154])^(a[59] & b[155])^(a[58] & b[156])^(a[57] & b[157])^(a[56] & b[158])^(a[55] & b[159])^(a[54] & b[160])^(a[53] & b[161])^(a[52] & b[162])^(a[51] & b[163])^(a[50] & b[164])^(a[49] & b[165])^(a[48] & b[166])^(a[47] & b[167])^(a[46] & b[168])^(a[45] & b[169])^(a[44] & b[170])^(a[43] & b[171])^(a[42] & b[172])^(a[41] & b[173])^(a[40] & b[174])^(a[39] & b[175])^(a[38] & b[176])^(a[37] & b[177])^(a[36] & b[178])^(a[35] & b[179])^(a[34] & b[180])^(a[33] & b[181])^(a[32] & b[182])^(a[31] & b[183])^(a[30] & b[184])^(a[29] & b[185])^(a[28] & b[186])^(a[27] & b[187])^(a[26] & b[188])^(a[25] & b[189])^(a[24] & b[190])^(a[23] & b[191])^(a[22] & b[192])^(a[21] & b[193])^(a[20] & b[194])^(a[19] & b[195])^(a[18] & b[196])^(a[17] & b[197])^(a[16] & b[198])^(a[15] & b[199])^(a[14] & b[200])^(a[13] & b[201])^(a[12] & b[202])^(a[11] & b[203])^(a[10] & b[204])^(a[9] & b[205])^(a[8] & b[206])^(a[7] & b[207])^(a[6] & b[208])^(a[5] & b[209])^(a[4] & b[210])^(a[3] & b[211])^(a[2] & b[212])^(a[1] & b[213])^(a[0] & b[214]);
assign y[215] = (a[215] & b[0])^(a[214] & b[1])^(a[213] & b[2])^(a[212] & b[3])^(a[211] & b[4])^(a[210] & b[5])^(a[209] & b[6])^(a[208] & b[7])^(a[207] & b[8])^(a[206] & b[9])^(a[205] & b[10])^(a[204] & b[11])^(a[203] & b[12])^(a[202] & b[13])^(a[201] & b[14])^(a[200] & b[15])^(a[199] & b[16])^(a[198] & b[17])^(a[197] & b[18])^(a[196] & b[19])^(a[195] & b[20])^(a[194] & b[21])^(a[193] & b[22])^(a[192] & b[23])^(a[191] & b[24])^(a[190] & b[25])^(a[189] & b[26])^(a[188] & b[27])^(a[187] & b[28])^(a[186] & b[29])^(a[185] & b[30])^(a[184] & b[31])^(a[183] & b[32])^(a[182] & b[33])^(a[181] & b[34])^(a[180] & b[35])^(a[179] & b[36])^(a[178] & b[37])^(a[177] & b[38])^(a[176] & b[39])^(a[175] & b[40])^(a[174] & b[41])^(a[173] & b[42])^(a[172] & b[43])^(a[171] & b[44])^(a[170] & b[45])^(a[169] & b[46])^(a[168] & b[47])^(a[167] & b[48])^(a[166] & b[49])^(a[165] & b[50])^(a[164] & b[51])^(a[163] & b[52])^(a[162] & b[53])^(a[161] & b[54])^(a[160] & b[55])^(a[159] & b[56])^(a[158] & b[57])^(a[157] & b[58])^(a[156] & b[59])^(a[155] & b[60])^(a[154] & b[61])^(a[153] & b[62])^(a[152] & b[63])^(a[151] & b[64])^(a[150] & b[65])^(a[149] & b[66])^(a[148] & b[67])^(a[147] & b[68])^(a[146] & b[69])^(a[145] & b[70])^(a[144] & b[71])^(a[143] & b[72])^(a[142] & b[73])^(a[141] & b[74])^(a[140] & b[75])^(a[139] & b[76])^(a[138] & b[77])^(a[137] & b[78])^(a[136] & b[79])^(a[135] & b[80])^(a[134] & b[81])^(a[133] & b[82])^(a[132] & b[83])^(a[131] & b[84])^(a[130] & b[85])^(a[129] & b[86])^(a[128] & b[87])^(a[127] & b[88])^(a[126] & b[89])^(a[125] & b[90])^(a[124] & b[91])^(a[123] & b[92])^(a[122] & b[93])^(a[121] & b[94])^(a[120] & b[95])^(a[119] & b[96])^(a[118] & b[97])^(a[117] & b[98])^(a[116] & b[99])^(a[115] & b[100])^(a[114] & b[101])^(a[113] & b[102])^(a[112] & b[103])^(a[111] & b[104])^(a[110] & b[105])^(a[109] & b[106])^(a[108] & b[107])^(a[107] & b[108])^(a[106] & b[109])^(a[105] & b[110])^(a[104] & b[111])^(a[103] & b[112])^(a[102] & b[113])^(a[101] & b[114])^(a[100] & b[115])^(a[99] & b[116])^(a[98] & b[117])^(a[97] & b[118])^(a[96] & b[119])^(a[95] & b[120])^(a[94] & b[121])^(a[93] & b[122])^(a[92] & b[123])^(a[91] & b[124])^(a[90] & b[125])^(a[89] & b[126])^(a[88] & b[127])^(a[87] & b[128])^(a[86] & b[129])^(a[85] & b[130])^(a[84] & b[131])^(a[83] & b[132])^(a[82] & b[133])^(a[81] & b[134])^(a[80] & b[135])^(a[79] & b[136])^(a[78] & b[137])^(a[77] & b[138])^(a[76] & b[139])^(a[75] & b[140])^(a[74] & b[141])^(a[73] & b[142])^(a[72] & b[143])^(a[71] & b[144])^(a[70] & b[145])^(a[69] & b[146])^(a[68] & b[147])^(a[67] & b[148])^(a[66] & b[149])^(a[65] & b[150])^(a[64] & b[151])^(a[63] & b[152])^(a[62] & b[153])^(a[61] & b[154])^(a[60] & b[155])^(a[59] & b[156])^(a[58] & b[157])^(a[57] & b[158])^(a[56] & b[159])^(a[55] & b[160])^(a[54] & b[161])^(a[53] & b[162])^(a[52] & b[163])^(a[51] & b[164])^(a[50] & b[165])^(a[49] & b[166])^(a[48] & b[167])^(a[47] & b[168])^(a[46] & b[169])^(a[45] & b[170])^(a[44] & b[171])^(a[43] & b[172])^(a[42] & b[173])^(a[41] & b[174])^(a[40] & b[175])^(a[39] & b[176])^(a[38] & b[177])^(a[37] & b[178])^(a[36] & b[179])^(a[35] & b[180])^(a[34] & b[181])^(a[33] & b[182])^(a[32] & b[183])^(a[31] & b[184])^(a[30] & b[185])^(a[29] & b[186])^(a[28] & b[187])^(a[27] & b[188])^(a[26] & b[189])^(a[25] & b[190])^(a[24] & b[191])^(a[23] & b[192])^(a[22] & b[193])^(a[21] & b[194])^(a[20] & b[195])^(a[19] & b[196])^(a[18] & b[197])^(a[17] & b[198])^(a[16] & b[199])^(a[15] & b[200])^(a[14] & b[201])^(a[13] & b[202])^(a[12] & b[203])^(a[11] & b[204])^(a[10] & b[205])^(a[9] & b[206])^(a[8] & b[207])^(a[7] & b[208])^(a[6] & b[209])^(a[5] & b[210])^(a[4] & b[211])^(a[3] & b[212])^(a[2] & b[213])^(a[1] & b[214])^(a[0] & b[215]);
assign y[216] = (a[216] & b[0])^(a[215] & b[1])^(a[214] & b[2])^(a[213] & b[3])^(a[212] & b[4])^(a[211] & b[5])^(a[210] & b[6])^(a[209] & b[7])^(a[208] & b[8])^(a[207] & b[9])^(a[206] & b[10])^(a[205] & b[11])^(a[204] & b[12])^(a[203] & b[13])^(a[202] & b[14])^(a[201] & b[15])^(a[200] & b[16])^(a[199] & b[17])^(a[198] & b[18])^(a[197] & b[19])^(a[196] & b[20])^(a[195] & b[21])^(a[194] & b[22])^(a[193] & b[23])^(a[192] & b[24])^(a[191] & b[25])^(a[190] & b[26])^(a[189] & b[27])^(a[188] & b[28])^(a[187] & b[29])^(a[186] & b[30])^(a[185] & b[31])^(a[184] & b[32])^(a[183] & b[33])^(a[182] & b[34])^(a[181] & b[35])^(a[180] & b[36])^(a[179] & b[37])^(a[178] & b[38])^(a[177] & b[39])^(a[176] & b[40])^(a[175] & b[41])^(a[174] & b[42])^(a[173] & b[43])^(a[172] & b[44])^(a[171] & b[45])^(a[170] & b[46])^(a[169] & b[47])^(a[168] & b[48])^(a[167] & b[49])^(a[166] & b[50])^(a[165] & b[51])^(a[164] & b[52])^(a[163] & b[53])^(a[162] & b[54])^(a[161] & b[55])^(a[160] & b[56])^(a[159] & b[57])^(a[158] & b[58])^(a[157] & b[59])^(a[156] & b[60])^(a[155] & b[61])^(a[154] & b[62])^(a[153] & b[63])^(a[152] & b[64])^(a[151] & b[65])^(a[150] & b[66])^(a[149] & b[67])^(a[148] & b[68])^(a[147] & b[69])^(a[146] & b[70])^(a[145] & b[71])^(a[144] & b[72])^(a[143] & b[73])^(a[142] & b[74])^(a[141] & b[75])^(a[140] & b[76])^(a[139] & b[77])^(a[138] & b[78])^(a[137] & b[79])^(a[136] & b[80])^(a[135] & b[81])^(a[134] & b[82])^(a[133] & b[83])^(a[132] & b[84])^(a[131] & b[85])^(a[130] & b[86])^(a[129] & b[87])^(a[128] & b[88])^(a[127] & b[89])^(a[126] & b[90])^(a[125] & b[91])^(a[124] & b[92])^(a[123] & b[93])^(a[122] & b[94])^(a[121] & b[95])^(a[120] & b[96])^(a[119] & b[97])^(a[118] & b[98])^(a[117] & b[99])^(a[116] & b[100])^(a[115] & b[101])^(a[114] & b[102])^(a[113] & b[103])^(a[112] & b[104])^(a[111] & b[105])^(a[110] & b[106])^(a[109] & b[107])^(a[108] & b[108])^(a[107] & b[109])^(a[106] & b[110])^(a[105] & b[111])^(a[104] & b[112])^(a[103] & b[113])^(a[102] & b[114])^(a[101] & b[115])^(a[100] & b[116])^(a[99] & b[117])^(a[98] & b[118])^(a[97] & b[119])^(a[96] & b[120])^(a[95] & b[121])^(a[94] & b[122])^(a[93] & b[123])^(a[92] & b[124])^(a[91] & b[125])^(a[90] & b[126])^(a[89] & b[127])^(a[88] & b[128])^(a[87] & b[129])^(a[86] & b[130])^(a[85] & b[131])^(a[84] & b[132])^(a[83] & b[133])^(a[82] & b[134])^(a[81] & b[135])^(a[80] & b[136])^(a[79] & b[137])^(a[78] & b[138])^(a[77] & b[139])^(a[76] & b[140])^(a[75] & b[141])^(a[74] & b[142])^(a[73] & b[143])^(a[72] & b[144])^(a[71] & b[145])^(a[70] & b[146])^(a[69] & b[147])^(a[68] & b[148])^(a[67] & b[149])^(a[66] & b[150])^(a[65] & b[151])^(a[64] & b[152])^(a[63] & b[153])^(a[62] & b[154])^(a[61] & b[155])^(a[60] & b[156])^(a[59] & b[157])^(a[58] & b[158])^(a[57] & b[159])^(a[56] & b[160])^(a[55] & b[161])^(a[54] & b[162])^(a[53] & b[163])^(a[52] & b[164])^(a[51] & b[165])^(a[50] & b[166])^(a[49] & b[167])^(a[48] & b[168])^(a[47] & b[169])^(a[46] & b[170])^(a[45] & b[171])^(a[44] & b[172])^(a[43] & b[173])^(a[42] & b[174])^(a[41] & b[175])^(a[40] & b[176])^(a[39] & b[177])^(a[38] & b[178])^(a[37] & b[179])^(a[36] & b[180])^(a[35] & b[181])^(a[34] & b[182])^(a[33] & b[183])^(a[32] & b[184])^(a[31] & b[185])^(a[30] & b[186])^(a[29] & b[187])^(a[28] & b[188])^(a[27] & b[189])^(a[26] & b[190])^(a[25] & b[191])^(a[24] & b[192])^(a[23] & b[193])^(a[22] & b[194])^(a[21] & b[195])^(a[20] & b[196])^(a[19] & b[197])^(a[18] & b[198])^(a[17] & b[199])^(a[16] & b[200])^(a[15] & b[201])^(a[14] & b[202])^(a[13] & b[203])^(a[12] & b[204])^(a[11] & b[205])^(a[10] & b[206])^(a[9] & b[207])^(a[8] & b[208])^(a[7] & b[209])^(a[6] & b[210])^(a[5] & b[211])^(a[4] & b[212])^(a[3] & b[213])^(a[2] & b[214])^(a[1] & b[215])^(a[0] & b[216]);
assign y[217] = (a[217] & b[0])^(a[216] & b[1])^(a[215] & b[2])^(a[214] & b[3])^(a[213] & b[4])^(a[212] & b[5])^(a[211] & b[6])^(a[210] & b[7])^(a[209] & b[8])^(a[208] & b[9])^(a[207] & b[10])^(a[206] & b[11])^(a[205] & b[12])^(a[204] & b[13])^(a[203] & b[14])^(a[202] & b[15])^(a[201] & b[16])^(a[200] & b[17])^(a[199] & b[18])^(a[198] & b[19])^(a[197] & b[20])^(a[196] & b[21])^(a[195] & b[22])^(a[194] & b[23])^(a[193] & b[24])^(a[192] & b[25])^(a[191] & b[26])^(a[190] & b[27])^(a[189] & b[28])^(a[188] & b[29])^(a[187] & b[30])^(a[186] & b[31])^(a[185] & b[32])^(a[184] & b[33])^(a[183] & b[34])^(a[182] & b[35])^(a[181] & b[36])^(a[180] & b[37])^(a[179] & b[38])^(a[178] & b[39])^(a[177] & b[40])^(a[176] & b[41])^(a[175] & b[42])^(a[174] & b[43])^(a[173] & b[44])^(a[172] & b[45])^(a[171] & b[46])^(a[170] & b[47])^(a[169] & b[48])^(a[168] & b[49])^(a[167] & b[50])^(a[166] & b[51])^(a[165] & b[52])^(a[164] & b[53])^(a[163] & b[54])^(a[162] & b[55])^(a[161] & b[56])^(a[160] & b[57])^(a[159] & b[58])^(a[158] & b[59])^(a[157] & b[60])^(a[156] & b[61])^(a[155] & b[62])^(a[154] & b[63])^(a[153] & b[64])^(a[152] & b[65])^(a[151] & b[66])^(a[150] & b[67])^(a[149] & b[68])^(a[148] & b[69])^(a[147] & b[70])^(a[146] & b[71])^(a[145] & b[72])^(a[144] & b[73])^(a[143] & b[74])^(a[142] & b[75])^(a[141] & b[76])^(a[140] & b[77])^(a[139] & b[78])^(a[138] & b[79])^(a[137] & b[80])^(a[136] & b[81])^(a[135] & b[82])^(a[134] & b[83])^(a[133] & b[84])^(a[132] & b[85])^(a[131] & b[86])^(a[130] & b[87])^(a[129] & b[88])^(a[128] & b[89])^(a[127] & b[90])^(a[126] & b[91])^(a[125] & b[92])^(a[124] & b[93])^(a[123] & b[94])^(a[122] & b[95])^(a[121] & b[96])^(a[120] & b[97])^(a[119] & b[98])^(a[118] & b[99])^(a[117] & b[100])^(a[116] & b[101])^(a[115] & b[102])^(a[114] & b[103])^(a[113] & b[104])^(a[112] & b[105])^(a[111] & b[106])^(a[110] & b[107])^(a[109] & b[108])^(a[108] & b[109])^(a[107] & b[110])^(a[106] & b[111])^(a[105] & b[112])^(a[104] & b[113])^(a[103] & b[114])^(a[102] & b[115])^(a[101] & b[116])^(a[100] & b[117])^(a[99] & b[118])^(a[98] & b[119])^(a[97] & b[120])^(a[96] & b[121])^(a[95] & b[122])^(a[94] & b[123])^(a[93] & b[124])^(a[92] & b[125])^(a[91] & b[126])^(a[90] & b[127])^(a[89] & b[128])^(a[88] & b[129])^(a[87] & b[130])^(a[86] & b[131])^(a[85] & b[132])^(a[84] & b[133])^(a[83] & b[134])^(a[82] & b[135])^(a[81] & b[136])^(a[80] & b[137])^(a[79] & b[138])^(a[78] & b[139])^(a[77] & b[140])^(a[76] & b[141])^(a[75] & b[142])^(a[74] & b[143])^(a[73] & b[144])^(a[72] & b[145])^(a[71] & b[146])^(a[70] & b[147])^(a[69] & b[148])^(a[68] & b[149])^(a[67] & b[150])^(a[66] & b[151])^(a[65] & b[152])^(a[64] & b[153])^(a[63] & b[154])^(a[62] & b[155])^(a[61] & b[156])^(a[60] & b[157])^(a[59] & b[158])^(a[58] & b[159])^(a[57] & b[160])^(a[56] & b[161])^(a[55] & b[162])^(a[54] & b[163])^(a[53] & b[164])^(a[52] & b[165])^(a[51] & b[166])^(a[50] & b[167])^(a[49] & b[168])^(a[48] & b[169])^(a[47] & b[170])^(a[46] & b[171])^(a[45] & b[172])^(a[44] & b[173])^(a[43] & b[174])^(a[42] & b[175])^(a[41] & b[176])^(a[40] & b[177])^(a[39] & b[178])^(a[38] & b[179])^(a[37] & b[180])^(a[36] & b[181])^(a[35] & b[182])^(a[34] & b[183])^(a[33] & b[184])^(a[32] & b[185])^(a[31] & b[186])^(a[30] & b[187])^(a[29] & b[188])^(a[28] & b[189])^(a[27] & b[190])^(a[26] & b[191])^(a[25] & b[192])^(a[24] & b[193])^(a[23] & b[194])^(a[22] & b[195])^(a[21] & b[196])^(a[20] & b[197])^(a[19] & b[198])^(a[18] & b[199])^(a[17] & b[200])^(a[16] & b[201])^(a[15] & b[202])^(a[14] & b[203])^(a[13] & b[204])^(a[12] & b[205])^(a[11] & b[206])^(a[10] & b[207])^(a[9] & b[208])^(a[8] & b[209])^(a[7] & b[210])^(a[6] & b[211])^(a[5] & b[212])^(a[4] & b[213])^(a[3] & b[214])^(a[2] & b[215])^(a[1] & b[216])^(a[0] & b[217]);
assign y[218] = (a[218] & b[0])^(a[217] & b[1])^(a[216] & b[2])^(a[215] & b[3])^(a[214] & b[4])^(a[213] & b[5])^(a[212] & b[6])^(a[211] & b[7])^(a[210] & b[8])^(a[209] & b[9])^(a[208] & b[10])^(a[207] & b[11])^(a[206] & b[12])^(a[205] & b[13])^(a[204] & b[14])^(a[203] & b[15])^(a[202] & b[16])^(a[201] & b[17])^(a[200] & b[18])^(a[199] & b[19])^(a[198] & b[20])^(a[197] & b[21])^(a[196] & b[22])^(a[195] & b[23])^(a[194] & b[24])^(a[193] & b[25])^(a[192] & b[26])^(a[191] & b[27])^(a[190] & b[28])^(a[189] & b[29])^(a[188] & b[30])^(a[187] & b[31])^(a[186] & b[32])^(a[185] & b[33])^(a[184] & b[34])^(a[183] & b[35])^(a[182] & b[36])^(a[181] & b[37])^(a[180] & b[38])^(a[179] & b[39])^(a[178] & b[40])^(a[177] & b[41])^(a[176] & b[42])^(a[175] & b[43])^(a[174] & b[44])^(a[173] & b[45])^(a[172] & b[46])^(a[171] & b[47])^(a[170] & b[48])^(a[169] & b[49])^(a[168] & b[50])^(a[167] & b[51])^(a[166] & b[52])^(a[165] & b[53])^(a[164] & b[54])^(a[163] & b[55])^(a[162] & b[56])^(a[161] & b[57])^(a[160] & b[58])^(a[159] & b[59])^(a[158] & b[60])^(a[157] & b[61])^(a[156] & b[62])^(a[155] & b[63])^(a[154] & b[64])^(a[153] & b[65])^(a[152] & b[66])^(a[151] & b[67])^(a[150] & b[68])^(a[149] & b[69])^(a[148] & b[70])^(a[147] & b[71])^(a[146] & b[72])^(a[145] & b[73])^(a[144] & b[74])^(a[143] & b[75])^(a[142] & b[76])^(a[141] & b[77])^(a[140] & b[78])^(a[139] & b[79])^(a[138] & b[80])^(a[137] & b[81])^(a[136] & b[82])^(a[135] & b[83])^(a[134] & b[84])^(a[133] & b[85])^(a[132] & b[86])^(a[131] & b[87])^(a[130] & b[88])^(a[129] & b[89])^(a[128] & b[90])^(a[127] & b[91])^(a[126] & b[92])^(a[125] & b[93])^(a[124] & b[94])^(a[123] & b[95])^(a[122] & b[96])^(a[121] & b[97])^(a[120] & b[98])^(a[119] & b[99])^(a[118] & b[100])^(a[117] & b[101])^(a[116] & b[102])^(a[115] & b[103])^(a[114] & b[104])^(a[113] & b[105])^(a[112] & b[106])^(a[111] & b[107])^(a[110] & b[108])^(a[109] & b[109])^(a[108] & b[110])^(a[107] & b[111])^(a[106] & b[112])^(a[105] & b[113])^(a[104] & b[114])^(a[103] & b[115])^(a[102] & b[116])^(a[101] & b[117])^(a[100] & b[118])^(a[99] & b[119])^(a[98] & b[120])^(a[97] & b[121])^(a[96] & b[122])^(a[95] & b[123])^(a[94] & b[124])^(a[93] & b[125])^(a[92] & b[126])^(a[91] & b[127])^(a[90] & b[128])^(a[89] & b[129])^(a[88] & b[130])^(a[87] & b[131])^(a[86] & b[132])^(a[85] & b[133])^(a[84] & b[134])^(a[83] & b[135])^(a[82] & b[136])^(a[81] & b[137])^(a[80] & b[138])^(a[79] & b[139])^(a[78] & b[140])^(a[77] & b[141])^(a[76] & b[142])^(a[75] & b[143])^(a[74] & b[144])^(a[73] & b[145])^(a[72] & b[146])^(a[71] & b[147])^(a[70] & b[148])^(a[69] & b[149])^(a[68] & b[150])^(a[67] & b[151])^(a[66] & b[152])^(a[65] & b[153])^(a[64] & b[154])^(a[63] & b[155])^(a[62] & b[156])^(a[61] & b[157])^(a[60] & b[158])^(a[59] & b[159])^(a[58] & b[160])^(a[57] & b[161])^(a[56] & b[162])^(a[55] & b[163])^(a[54] & b[164])^(a[53] & b[165])^(a[52] & b[166])^(a[51] & b[167])^(a[50] & b[168])^(a[49] & b[169])^(a[48] & b[170])^(a[47] & b[171])^(a[46] & b[172])^(a[45] & b[173])^(a[44] & b[174])^(a[43] & b[175])^(a[42] & b[176])^(a[41] & b[177])^(a[40] & b[178])^(a[39] & b[179])^(a[38] & b[180])^(a[37] & b[181])^(a[36] & b[182])^(a[35] & b[183])^(a[34] & b[184])^(a[33] & b[185])^(a[32] & b[186])^(a[31] & b[187])^(a[30] & b[188])^(a[29] & b[189])^(a[28] & b[190])^(a[27] & b[191])^(a[26] & b[192])^(a[25] & b[193])^(a[24] & b[194])^(a[23] & b[195])^(a[22] & b[196])^(a[21] & b[197])^(a[20] & b[198])^(a[19] & b[199])^(a[18] & b[200])^(a[17] & b[201])^(a[16] & b[202])^(a[15] & b[203])^(a[14] & b[204])^(a[13] & b[205])^(a[12] & b[206])^(a[11] & b[207])^(a[10] & b[208])^(a[9] & b[209])^(a[8] & b[210])^(a[7] & b[211])^(a[6] & b[212])^(a[5] & b[213])^(a[4] & b[214])^(a[3] & b[215])^(a[2] & b[216])^(a[1] & b[217])^(a[0] & b[218]);
assign y[219] = (a[219] & b[0])^(a[218] & b[1])^(a[217] & b[2])^(a[216] & b[3])^(a[215] & b[4])^(a[214] & b[5])^(a[213] & b[6])^(a[212] & b[7])^(a[211] & b[8])^(a[210] & b[9])^(a[209] & b[10])^(a[208] & b[11])^(a[207] & b[12])^(a[206] & b[13])^(a[205] & b[14])^(a[204] & b[15])^(a[203] & b[16])^(a[202] & b[17])^(a[201] & b[18])^(a[200] & b[19])^(a[199] & b[20])^(a[198] & b[21])^(a[197] & b[22])^(a[196] & b[23])^(a[195] & b[24])^(a[194] & b[25])^(a[193] & b[26])^(a[192] & b[27])^(a[191] & b[28])^(a[190] & b[29])^(a[189] & b[30])^(a[188] & b[31])^(a[187] & b[32])^(a[186] & b[33])^(a[185] & b[34])^(a[184] & b[35])^(a[183] & b[36])^(a[182] & b[37])^(a[181] & b[38])^(a[180] & b[39])^(a[179] & b[40])^(a[178] & b[41])^(a[177] & b[42])^(a[176] & b[43])^(a[175] & b[44])^(a[174] & b[45])^(a[173] & b[46])^(a[172] & b[47])^(a[171] & b[48])^(a[170] & b[49])^(a[169] & b[50])^(a[168] & b[51])^(a[167] & b[52])^(a[166] & b[53])^(a[165] & b[54])^(a[164] & b[55])^(a[163] & b[56])^(a[162] & b[57])^(a[161] & b[58])^(a[160] & b[59])^(a[159] & b[60])^(a[158] & b[61])^(a[157] & b[62])^(a[156] & b[63])^(a[155] & b[64])^(a[154] & b[65])^(a[153] & b[66])^(a[152] & b[67])^(a[151] & b[68])^(a[150] & b[69])^(a[149] & b[70])^(a[148] & b[71])^(a[147] & b[72])^(a[146] & b[73])^(a[145] & b[74])^(a[144] & b[75])^(a[143] & b[76])^(a[142] & b[77])^(a[141] & b[78])^(a[140] & b[79])^(a[139] & b[80])^(a[138] & b[81])^(a[137] & b[82])^(a[136] & b[83])^(a[135] & b[84])^(a[134] & b[85])^(a[133] & b[86])^(a[132] & b[87])^(a[131] & b[88])^(a[130] & b[89])^(a[129] & b[90])^(a[128] & b[91])^(a[127] & b[92])^(a[126] & b[93])^(a[125] & b[94])^(a[124] & b[95])^(a[123] & b[96])^(a[122] & b[97])^(a[121] & b[98])^(a[120] & b[99])^(a[119] & b[100])^(a[118] & b[101])^(a[117] & b[102])^(a[116] & b[103])^(a[115] & b[104])^(a[114] & b[105])^(a[113] & b[106])^(a[112] & b[107])^(a[111] & b[108])^(a[110] & b[109])^(a[109] & b[110])^(a[108] & b[111])^(a[107] & b[112])^(a[106] & b[113])^(a[105] & b[114])^(a[104] & b[115])^(a[103] & b[116])^(a[102] & b[117])^(a[101] & b[118])^(a[100] & b[119])^(a[99] & b[120])^(a[98] & b[121])^(a[97] & b[122])^(a[96] & b[123])^(a[95] & b[124])^(a[94] & b[125])^(a[93] & b[126])^(a[92] & b[127])^(a[91] & b[128])^(a[90] & b[129])^(a[89] & b[130])^(a[88] & b[131])^(a[87] & b[132])^(a[86] & b[133])^(a[85] & b[134])^(a[84] & b[135])^(a[83] & b[136])^(a[82] & b[137])^(a[81] & b[138])^(a[80] & b[139])^(a[79] & b[140])^(a[78] & b[141])^(a[77] & b[142])^(a[76] & b[143])^(a[75] & b[144])^(a[74] & b[145])^(a[73] & b[146])^(a[72] & b[147])^(a[71] & b[148])^(a[70] & b[149])^(a[69] & b[150])^(a[68] & b[151])^(a[67] & b[152])^(a[66] & b[153])^(a[65] & b[154])^(a[64] & b[155])^(a[63] & b[156])^(a[62] & b[157])^(a[61] & b[158])^(a[60] & b[159])^(a[59] & b[160])^(a[58] & b[161])^(a[57] & b[162])^(a[56] & b[163])^(a[55] & b[164])^(a[54] & b[165])^(a[53] & b[166])^(a[52] & b[167])^(a[51] & b[168])^(a[50] & b[169])^(a[49] & b[170])^(a[48] & b[171])^(a[47] & b[172])^(a[46] & b[173])^(a[45] & b[174])^(a[44] & b[175])^(a[43] & b[176])^(a[42] & b[177])^(a[41] & b[178])^(a[40] & b[179])^(a[39] & b[180])^(a[38] & b[181])^(a[37] & b[182])^(a[36] & b[183])^(a[35] & b[184])^(a[34] & b[185])^(a[33] & b[186])^(a[32] & b[187])^(a[31] & b[188])^(a[30] & b[189])^(a[29] & b[190])^(a[28] & b[191])^(a[27] & b[192])^(a[26] & b[193])^(a[25] & b[194])^(a[24] & b[195])^(a[23] & b[196])^(a[22] & b[197])^(a[21] & b[198])^(a[20] & b[199])^(a[19] & b[200])^(a[18] & b[201])^(a[17] & b[202])^(a[16] & b[203])^(a[15] & b[204])^(a[14] & b[205])^(a[13] & b[206])^(a[12] & b[207])^(a[11] & b[208])^(a[10] & b[209])^(a[9] & b[210])^(a[8] & b[211])^(a[7] & b[212])^(a[6] & b[213])^(a[5] & b[214])^(a[4] & b[215])^(a[3] & b[216])^(a[2] & b[217])^(a[1] & b[218])^(a[0] & b[219]);
assign y[220] = (a[220] & b[0])^(a[219] & b[1])^(a[218] & b[2])^(a[217] & b[3])^(a[216] & b[4])^(a[215] & b[5])^(a[214] & b[6])^(a[213] & b[7])^(a[212] & b[8])^(a[211] & b[9])^(a[210] & b[10])^(a[209] & b[11])^(a[208] & b[12])^(a[207] & b[13])^(a[206] & b[14])^(a[205] & b[15])^(a[204] & b[16])^(a[203] & b[17])^(a[202] & b[18])^(a[201] & b[19])^(a[200] & b[20])^(a[199] & b[21])^(a[198] & b[22])^(a[197] & b[23])^(a[196] & b[24])^(a[195] & b[25])^(a[194] & b[26])^(a[193] & b[27])^(a[192] & b[28])^(a[191] & b[29])^(a[190] & b[30])^(a[189] & b[31])^(a[188] & b[32])^(a[187] & b[33])^(a[186] & b[34])^(a[185] & b[35])^(a[184] & b[36])^(a[183] & b[37])^(a[182] & b[38])^(a[181] & b[39])^(a[180] & b[40])^(a[179] & b[41])^(a[178] & b[42])^(a[177] & b[43])^(a[176] & b[44])^(a[175] & b[45])^(a[174] & b[46])^(a[173] & b[47])^(a[172] & b[48])^(a[171] & b[49])^(a[170] & b[50])^(a[169] & b[51])^(a[168] & b[52])^(a[167] & b[53])^(a[166] & b[54])^(a[165] & b[55])^(a[164] & b[56])^(a[163] & b[57])^(a[162] & b[58])^(a[161] & b[59])^(a[160] & b[60])^(a[159] & b[61])^(a[158] & b[62])^(a[157] & b[63])^(a[156] & b[64])^(a[155] & b[65])^(a[154] & b[66])^(a[153] & b[67])^(a[152] & b[68])^(a[151] & b[69])^(a[150] & b[70])^(a[149] & b[71])^(a[148] & b[72])^(a[147] & b[73])^(a[146] & b[74])^(a[145] & b[75])^(a[144] & b[76])^(a[143] & b[77])^(a[142] & b[78])^(a[141] & b[79])^(a[140] & b[80])^(a[139] & b[81])^(a[138] & b[82])^(a[137] & b[83])^(a[136] & b[84])^(a[135] & b[85])^(a[134] & b[86])^(a[133] & b[87])^(a[132] & b[88])^(a[131] & b[89])^(a[130] & b[90])^(a[129] & b[91])^(a[128] & b[92])^(a[127] & b[93])^(a[126] & b[94])^(a[125] & b[95])^(a[124] & b[96])^(a[123] & b[97])^(a[122] & b[98])^(a[121] & b[99])^(a[120] & b[100])^(a[119] & b[101])^(a[118] & b[102])^(a[117] & b[103])^(a[116] & b[104])^(a[115] & b[105])^(a[114] & b[106])^(a[113] & b[107])^(a[112] & b[108])^(a[111] & b[109])^(a[110] & b[110])^(a[109] & b[111])^(a[108] & b[112])^(a[107] & b[113])^(a[106] & b[114])^(a[105] & b[115])^(a[104] & b[116])^(a[103] & b[117])^(a[102] & b[118])^(a[101] & b[119])^(a[100] & b[120])^(a[99] & b[121])^(a[98] & b[122])^(a[97] & b[123])^(a[96] & b[124])^(a[95] & b[125])^(a[94] & b[126])^(a[93] & b[127])^(a[92] & b[128])^(a[91] & b[129])^(a[90] & b[130])^(a[89] & b[131])^(a[88] & b[132])^(a[87] & b[133])^(a[86] & b[134])^(a[85] & b[135])^(a[84] & b[136])^(a[83] & b[137])^(a[82] & b[138])^(a[81] & b[139])^(a[80] & b[140])^(a[79] & b[141])^(a[78] & b[142])^(a[77] & b[143])^(a[76] & b[144])^(a[75] & b[145])^(a[74] & b[146])^(a[73] & b[147])^(a[72] & b[148])^(a[71] & b[149])^(a[70] & b[150])^(a[69] & b[151])^(a[68] & b[152])^(a[67] & b[153])^(a[66] & b[154])^(a[65] & b[155])^(a[64] & b[156])^(a[63] & b[157])^(a[62] & b[158])^(a[61] & b[159])^(a[60] & b[160])^(a[59] & b[161])^(a[58] & b[162])^(a[57] & b[163])^(a[56] & b[164])^(a[55] & b[165])^(a[54] & b[166])^(a[53] & b[167])^(a[52] & b[168])^(a[51] & b[169])^(a[50] & b[170])^(a[49] & b[171])^(a[48] & b[172])^(a[47] & b[173])^(a[46] & b[174])^(a[45] & b[175])^(a[44] & b[176])^(a[43] & b[177])^(a[42] & b[178])^(a[41] & b[179])^(a[40] & b[180])^(a[39] & b[181])^(a[38] & b[182])^(a[37] & b[183])^(a[36] & b[184])^(a[35] & b[185])^(a[34] & b[186])^(a[33] & b[187])^(a[32] & b[188])^(a[31] & b[189])^(a[30] & b[190])^(a[29] & b[191])^(a[28] & b[192])^(a[27] & b[193])^(a[26] & b[194])^(a[25] & b[195])^(a[24] & b[196])^(a[23] & b[197])^(a[22] & b[198])^(a[21] & b[199])^(a[20] & b[200])^(a[19] & b[201])^(a[18] & b[202])^(a[17] & b[203])^(a[16] & b[204])^(a[15] & b[205])^(a[14] & b[206])^(a[13] & b[207])^(a[12] & b[208])^(a[11] & b[209])^(a[10] & b[210])^(a[9] & b[211])^(a[8] & b[212])^(a[7] & b[213])^(a[6] & b[214])^(a[5] & b[215])^(a[4] & b[216])^(a[3] & b[217])^(a[2] & b[218])^(a[1] & b[219])^(a[0] & b[220]);
assign y[221] = (a[221] & b[0])^(a[220] & b[1])^(a[219] & b[2])^(a[218] & b[3])^(a[217] & b[4])^(a[216] & b[5])^(a[215] & b[6])^(a[214] & b[7])^(a[213] & b[8])^(a[212] & b[9])^(a[211] & b[10])^(a[210] & b[11])^(a[209] & b[12])^(a[208] & b[13])^(a[207] & b[14])^(a[206] & b[15])^(a[205] & b[16])^(a[204] & b[17])^(a[203] & b[18])^(a[202] & b[19])^(a[201] & b[20])^(a[200] & b[21])^(a[199] & b[22])^(a[198] & b[23])^(a[197] & b[24])^(a[196] & b[25])^(a[195] & b[26])^(a[194] & b[27])^(a[193] & b[28])^(a[192] & b[29])^(a[191] & b[30])^(a[190] & b[31])^(a[189] & b[32])^(a[188] & b[33])^(a[187] & b[34])^(a[186] & b[35])^(a[185] & b[36])^(a[184] & b[37])^(a[183] & b[38])^(a[182] & b[39])^(a[181] & b[40])^(a[180] & b[41])^(a[179] & b[42])^(a[178] & b[43])^(a[177] & b[44])^(a[176] & b[45])^(a[175] & b[46])^(a[174] & b[47])^(a[173] & b[48])^(a[172] & b[49])^(a[171] & b[50])^(a[170] & b[51])^(a[169] & b[52])^(a[168] & b[53])^(a[167] & b[54])^(a[166] & b[55])^(a[165] & b[56])^(a[164] & b[57])^(a[163] & b[58])^(a[162] & b[59])^(a[161] & b[60])^(a[160] & b[61])^(a[159] & b[62])^(a[158] & b[63])^(a[157] & b[64])^(a[156] & b[65])^(a[155] & b[66])^(a[154] & b[67])^(a[153] & b[68])^(a[152] & b[69])^(a[151] & b[70])^(a[150] & b[71])^(a[149] & b[72])^(a[148] & b[73])^(a[147] & b[74])^(a[146] & b[75])^(a[145] & b[76])^(a[144] & b[77])^(a[143] & b[78])^(a[142] & b[79])^(a[141] & b[80])^(a[140] & b[81])^(a[139] & b[82])^(a[138] & b[83])^(a[137] & b[84])^(a[136] & b[85])^(a[135] & b[86])^(a[134] & b[87])^(a[133] & b[88])^(a[132] & b[89])^(a[131] & b[90])^(a[130] & b[91])^(a[129] & b[92])^(a[128] & b[93])^(a[127] & b[94])^(a[126] & b[95])^(a[125] & b[96])^(a[124] & b[97])^(a[123] & b[98])^(a[122] & b[99])^(a[121] & b[100])^(a[120] & b[101])^(a[119] & b[102])^(a[118] & b[103])^(a[117] & b[104])^(a[116] & b[105])^(a[115] & b[106])^(a[114] & b[107])^(a[113] & b[108])^(a[112] & b[109])^(a[111] & b[110])^(a[110] & b[111])^(a[109] & b[112])^(a[108] & b[113])^(a[107] & b[114])^(a[106] & b[115])^(a[105] & b[116])^(a[104] & b[117])^(a[103] & b[118])^(a[102] & b[119])^(a[101] & b[120])^(a[100] & b[121])^(a[99] & b[122])^(a[98] & b[123])^(a[97] & b[124])^(a[96] & b[125])^(a[95] & b[126])^(a[94] & b[127])^(a[93] & b[128])^(a[92] & b[129])^(a[91] & b[130])^(a[90] & b[131])^(a[89] & b[132])^(a[88] & b[133])^(a[87] & b[134])^(a[86] & b[135])^(a[85] & b[136])^(a[84] & b[137])^(a[83] & b[138])^(a[82] & b[139])^(a[81] & b[140])^(a[80] & b[141])^(a[79] & b[142])^(a[78] & b[143])^(a[77] & b[144])^(a[76] & b[145])^(a[75] & b[146])^(a[74] & b[147])^(a[73] & b[148])^(a[72] & b[149])^(a[71] & b[150])^(a[70] & b[151])^(a[69] & b[152])^(a[68] & b[153])^(a[67] & b[154])^(a[66] & b[155])^(a[65] & b[156])^(a[64] & b[157])^(a[63] & b[158])^(a[62] & b[159])^(a[61] & b[160])^(a[60] & b[161])^(a[59] & b[162])^(a[58] & b[163])^(a[57] & b[164])^(a[56] & b[165])^(a[55] & b[166])^(a[54] & b[167])^(a[53] & b[168])^(a[52] & b[169])^(a[51] & b[170])^(a[50] & b[171])^(a[49] & b[172])^(a[48] & b[173])^(a[47] & b[174])^(a[46] & b[175])^(a[45] & b[176])^(a[44] & b[177])^(a[43] & b[178])^(a[42] & b[179])^(a[41] & b[180])^(a[40] & b[181])^(a[39] & b[182])^(a[38] & b[183])^(a[37] & b[184])^(a[36] & b[185])^(a[35] & b[186])^(a[34] & b[187])^(a[33] & b[188])^(a[32] & b[189])^(a[31] & b[190])^(a[30] & b[191])^(a[29] & b[192])^(a[28] & b[193])^(a[27] & b[194])^(a[26] & b[195])^(a[25] & b[196])^(a[24] & b[197])^(a[23] & b[198])^(a[22] & b[199])^(a[21] & b[200])^(a[20] & b[201])^(a[19] & b[202])^(a[18] & b[203])^(a[17] & b[204])^(a[16] & b[205])^(a[15] & b[206])^(a[14] & b[207])^(a[13] & b[208])^(a[12] & b[209])^(a[11] & b[210])^(a[10] & b[211])^(a[9] & b[212])^(a[8] & b[213])^(a[7] & b[214])^(a[6] & b[215])^(a[5] & b[216])^(a[4] & b[217])^(a[3] & b[218])^(a[2] & b[219])^(a[1] & b[220])^(a[0] & b[221]);
assign y[222] = (a[222] & b[0])^(a[221] & b[1])^(a[220] & b[2])^(a[219] & b[3])^(a[218] & b[4])^(a[217] & b[5])^(a[216] & b[6])^(a[215] & b[7])^(a[214] & b[8])^(a[213] & b[9])^(a[212] & b[10])^(a[211] & b[11])^(a[210] & b[12])^(a[209] & b[13])^(a[208] & b[14])^(a[207] & b[15])^(a[206] & b[16])^(a[205] & b[17])^(a[204] & b[18])^(a[203] & b[19])^(a[202] & b[20])^(a[201] & b[21])^(a[200] & b[22])^(a[199] & b[23])^(a[198] & b[24])^(a[197] & b[25])^(a[196] & b[26])^(a[195] & b[27])^(a[194] & b[28])^(a[193] & b[29])^(a[192] & b[30])^(a[191] & b[31])^(a[190] & b[32])^(a[189] & b[33])^(a[188] & b[34])^(a[187] & b[35])^(a[186] & b[36])^(a[185] & b[37])^(a[184] & b[38])^(a[183] & b[39])^(a[182] & b[40])^(a[181] & b[41])^(a[180] & b[42])^(a[179] & b[43])^(a[178] & b[44])^(a[177] & b[45])^(a[176] & b[46])^(a[175] & b[47])^(a[174] & b[48])^(a[173] & b[49])^(a[172] & b[50])^(a[171] & b[51])^(a[170] & b[52])^(a[169] & b[53])^(a[168] & b[54])^(a[167] & b[55])^(a[166] & b[56])^(a[165] & b[57])^(a[164] & b[58])^(a[163] & b[59])^(a[162] & b[60])^(a[161] & b[61])^(a[160] & b[62])^(a[159] & b[63])^(a[158] & b[64])^(a[157] & b[65])^(a[156] & b[66])^(a[155] & b[67])^(a[154] & b[68])^(a[153] & b[69])^(a[152] & b[70])^(a[151] & b[71])^(a[150] & b[72])^(a[149] & b[73])^(a[148] & b[74])^(a[147] & b[75])^(a[146] & b[76])^(a[145] & b[77])^(a[144] & b[78])^(a[143] & b[79])^(a[142] & b[80])^(a[141] & b[81])^(a[140] & b[82])^(a[139] & b[83])^(a[138] & b[84])^(a[137] & b[85])^(a[136] & b[86])^(a[135] & b[87])^(a[134] & b[88])^(a[133] & b[89])^(a[132] & b[90])^(a[131] & b[91])^(a[130] & b[92])^(a[129] & b[93])^(a[128] & b[94])^(a[127] & b[95])^(a[126] & b[96])^(a[125] & b[97])^(a[124] & b[98])^(a[123] & b[99])^(a[122] & b[100])^(a[121] & b[101])^(a[120] & b[102])^(a[119] & b[103])^(a[118] & b[104])^(a[117] & b[105])^(a[116] & b[106])^(a[115] & b[107])^(a[114] & b[108])^(a[113] & b[109])^(a[112] & b[110])^(a[111] & b[111])^(a[110] & b[112])^(a[109] & b[113])^(a[108] & b[114])^(a[107] & b[115])^(a[106] & b[116])^(a[105] & b[117])^(a[104] & b[118])^(a[103] & b[119])^(a[102] & b[120])^(a[101] & b[121])^(a[100] & b[122])^(a[99] & b[123])^(a[98] & b[124])^(a[97] & b[125])^(a[96] & b[126])^(a[95] & b[127])^(a[94] & b[128])^(a[93] & b[129])^(a[92] & b[130])^(a[91] & b[131])^(a[90] & b[132])^(a[89] & b[133])^(a[88] & b[134])^(a[87] & b[135])^(a[86] & b[136])^(a[85] & b[137])^(a[84] & b[138])^(a[83] & b[139])^(a[82] & b[140])^(a[81] & b[141])^(a[80] & b[142])^(a[79] & b[143])^(a[78] & b[144])^(a[77] & b[145])^(a[76] & b[146])^(a[75] & b[147])^(a[74] & b[148])^(a[73] & b[149])^(a[72] & b[150])^(a[71] & b[151])^(a[70] & b[152])^(a[69] & b[153])^(a[68] & b[154])^(a[67] & b[155])^(a[66] & b[156])^(a[65] & b[157])^(a[64] & b[158])^(a[63] & b[159])^(a[62] & b[160])^(a[61] & b[161])^(a[60] & b[162])^(a[59] & b[163])^(a[58] & b[164])^(a[57] & b[165])^(a[56] & b[166])^(a[55] & b[167])^(a[54] & b[168])^(a[53] & b[169])^(a[52] & b[170])^(a[51] & b[171])^(a[50] & b[172])^(a[49] & b[173])^(a[48] & b[174])^(a[47] & b[175])^(a[46] & b[176])^(a[45] & b[177])^(a[44] & b[178])^(a[43] & b[179])^(a[42] & b[180])^(a[41] & b[181])^(a[40] & b[182])^(a[39] & b[183])^(a[38] & b[184])^(a[37] & b[185])^(a[36] & b[186])^(a[35] & b[187])^(a[34] & b[188])^(a[33] & b[189])^(a[32] & b[190])^(a[31] & b[191])^(a[30] & b[192])^(a[29] & b[193])^(a[28] & b[194])^(a[27] & b[195])^(a[26] & b[196])^(a[25] & b[197])^(a[24] & b[198])^(a[23] & b[199])^(a[22] & b[200])^(a[21] & b[201])^(a[20] & b[202])^(a[19] & b[203])^(a[18] & b[204])^(a[17] & b[205])^(a[16] & b[206])^(a[15] & b[207])^(a[14] & b[208])^(a[13] & b[209])^(a[12] & b[210])^(a[11] & b[211])^(a[10] & b[212])^(a[9] & b[213])^(a[8] & b[214])^(a[7] & b[215])^(a[6] & b[216])^(a[5] & b[217])^(a[4] & b[218])^(a[3] & b[219])^(a[2] & b[220])^(a[1] & b[221])^(a[0] & b[222]);
assign y[223] = (a[223] & b[0])^(a[222] & b[1])^(a[221] & b[2])^(a[220] & b[3])^(a[219] & b[4])^(a[218] & b[5])^(a[217] & b[6])^(a[216] & b[7])^(a[215] & b[8])^(a[214] & b[9])^(a[213] & b[10])^(a[212] & b[11])^(a[211] & b[12])^(a[210] & b[13])^(a[209] & b[14])^(a[208] & b[15])^(a[207] & b[16])^(a[206] & b[17])^(a[205] & b[18])^(a[204] & b[19])^(a[203] & b[20])^(a[202] & b[21])^(a[201] & b[22])^(a[200] & b[23])^(a[199] & b[24])^(a[198] & b[25])^(a[197] & b[26])^(a[196] & b[27])^(a[195] & b[28])^(a[194] & b[29])^(a[193] & b[30])^(a[192] & b[31])^(a[191] & b[32])^(a[190] & b[33])^(a[189] & b[34])^(a[188] & b[35])^(a[187] & b[36])^(a[186] & b[37])^(a[185] & b[38])^(a[184] & b[39])^(a[183] & b[40])^(a[182] & b[41])^(a[181] & b[42])^(a[180] & b[43])^(a[179] & b[44])^(a[178] & b[45])^(a[177] & b[46])^(a[176] & b[47])^(a[175] & b[48])^(a[174] & b[49])^(a[173] & b[50])^(a[172] & b[51])^(a[171] & b[52])^(a[170] & b[53])^(a[169] & b[54])^(a[168] & b[55])^(a[167] & b[56])^(a[166] & b[57])^(a[165] & b[58])^(a[164] & b[59])^(a[163] & b[60])^(a[162] & b[61])^(a[161] & b[62])^(a[160] & b[63])^(a[159] & b[64])^(a[158] & b[65])^(a[157] & b[66])^(a[156] & b[67])^(a[155] & b[68])^(a[154] & b[69])^(a[153] & b[70])^(a[152] & b[71])^(a[151] & b[72])^(a[150] & b[73])^(a[149] & b[74])^(a[148] & b[75])^(a[147] & b[76])^(a[146] & b[77])^(a[145] & b[78])^(a[144] & b[79])^(a[143] & b[80])^(a[142] & b[81])^(a[141] & b[82])^(a[140] & b[83])^(a[139] & b[84])^(a[138] & b[85])^(a[137] & b[86])^(a[136] & b[87])^(a[135] & b[88])^(a[134] & b[89])^(a[133] & b[90])^(a[132] & b[91])^(a[131] & b[92])^(a[130] & b[93])^(a[129] & b[94])^(a[128] & b[95])^(a[127] & b[96])^(a[126] & b[97])^(a[125] & b[98])^(a[124] & b[99])^(a[123] & b[100])^(a[122] & b[101])^(a[121] & b[102])^(a[120] & b[103])^(a[119] & b[104])^(a[118] & b[105])^(a[117] & b[106])^(a[116] & b[107])^(a[115] & b[108])^(a[114] & b[109])^(a[113] & b[110])^(a[112] & b[111])^(a[111] & b[112])^(a[110] & b[113])^(a[109] & b[114])^(a[108] & b[115])^(a[107] & b[116])^(a[106] & b[117])^(a[105] & b[118])^(a[104] & b[119])^(a[103] & b[120])^(a[102] & b[121])^(a[101] & b[122])^(a[100] & b[123])^(a[99] & b[124])^(a[98] & b[125])^(a[97] & b[126])^(a[96] & b[127])^(a[95] & b[128])^(a[94] & b[129])^(a[93] & b[130])^(a[92] & b[131])^(a[91] & b[132])^(a[90] & b[133])^(a[89] & b[134])^(a[88] & b[135])^(a[87] & b[136])^(a[86] & b[137])^(a[85] & b[138])^(a[84] & b[139])^(a[83] & b[140])^(a[82] & b[141])^(a[81] & b[142])^(a[80] & b[143])^(a[79] & b[144])^(a[78] & b[145])^(a[77] & b[146])^(a[76] & b[147])^(a[75] & b[148])^(a[74] & b[149])^(a[73] & b[150])^(a[72] & b[151])^(a[71] & b[152])^(a[70] & b[153])^(a[69] & b[154])^(a[68] & b[155])^(a[67] & b[156])^(a[66] & b[157])^(a[65] & b[158])^(a[64] & b[159])^(a[63] & b[160])^(a[62] & b[161])^(a[61] & b[162])^(a[60] & b[163])^(a[59] & b[164])^(a[58] & b[165])^(a[57] & b[166])^(a[56] & b[167])^(a[55] & b[168])^(a[54] & b[169])^(a[53] & b[170])^(a[52] & b[171])^(a[51] & b[172])^(a[50] & b[173])^(a[49] & b[174])^(a[48] & b[175])^(a[47] & b[176])^(a[46] & b[177])^(a[45] & b[178])^(a[44] & b[179])^(a[43] & b[180])^(a[42] & b[181])^(a[41] & b[182])^(a[40] & b[183])^(a[39] & b[184])^(a[38] & b[185])^(a[37] & b[186])^(a[36] & b[187])^(a[35] & b[188])^(a[34] & b[189])^(a[33] & b[190])^(a[32] & b[191])^(a[31] & b[192])^(a[30] & b[193])^(a[29] & b[194])^(a[28] & b[195])^(a[27] & b[196])^(a[26] & b[197])^(a[25] & b[198])^(a[24] & b[199])^(a[23] & b[200])^(a[22] & b[201])^(a[21] & b[202])^(a[20] & b[203])^(a[19] & b[204])^(a[18] & b[205])^(a[17] & b[206])^(a[16] & b[207])^(a[15] & b[208])^(a[14] & b[209])^(a[13] & b[210])^(a[12] & b[211])^(a[11] & b[212])^(a[10] & b[213])^(a[9] & b[214])^(a[8] & b[215])^(a[7] & b[216])^(a[6] & b[217])^(a[5] & b[218])^(a[4] & b[219])^(a[3] & b[220])^(a[2] & b[221])^(a[1] & b[222])^(a[0] & b[223]);
assign y[224] = (a[224] & b[0])^(a[223] & b[1])^(a[222] & b[2])^(a[221] & b[3])^(a[220] & b[4])^(a[219] & b[5])^(a[218] & b[6])^(a[217] & b[7])^(a[216] & b[8])^(a[215] & b[9])^(a[214] & b[10])^(a[213] & b[11])^(a[212] & b[12])^(a[211] & b[13])^(a[210] & b[14])^(a[209] & b[15])^(a[208] & b[16])^(a[207] & b[17])^(a[206] & b[18])^(a[205] & b[19])^(a[204] & b[20])^(a[203] & b[21])^(a[202] & b[22])^(a[201] & b[23])^(a[200] & b[24])^(a[199] & b[25])^(a[198] & b[26])^(a[197] & b[27])^(a[196] & b[28])^(a[195] & b[29])^(a[194] & b[30])^(a[193] & b[31])^(a[192] & b[32])^(a[191] & b[33])^(a[190] & b[34])^(a[189] & b[35])^(a[188] & b[36])^(a[187] & b[37])^(a[186] & b[38])^(a[185] & b[39])^(a[184] & b[40])^(a[183] & b[41])^(a[182] & b[42])^(a[181] & b[43])^(a[180] & b[44])^(a[179] & b[45])^(a[178] & b[46])^(a[177] & b[47])^(a[176] & b[48])^(a[175] & b[49])^(a[174] & b[50])^(a[173] & b[51])^(a[172] & b[52])^(a[171] & b[53])^(a[170] & b[54])^(a[169] & b[55])^(a[168] & b[56])^(a[167] & b[57])^(a[166] & b[58])^(a[165] & b[59])^(a[164] & b[60])^(a[163] & b[61])^(a[162] & b[62])^(a[161] & b[63])^(a[160] & b[64])^(a[159] & b[65])^(a[158] & b[66])^(a[157] & b[67])^(a[156] & b[68])^(a[155] & b[69])^(a[154] & b[70])^(a[153] & b[71])^(a[152] & b[72])^(a[151] & b[73])^(a[150] & b[74])^(a[149] & b[75])^(a[148] & b[76])^(a[147] & b[77])^(a[146] & b[78])^(a[145] & b[79])^(a[144] & b[80])^(a[143] & b[81])^(a[142] & b[82])^(a[141] & b[83])^(a[140] & b[84])^(a[139] & b[85])^(a[138] & b[86])^(a[137] & b[87])^(a[136] & b[88])^(a[135] & b[89])^(a[134] & b[90])^(a[133] & b[91])^(a[132] & b[92])^(a[131] & b[93])^(a[130] & b[94])^(a[129] & b[95])^(a[128] & b[96])^(a[127] & b[97])^(a[126] & b[98])^(a[125] & b[99])^(a[124] & b[100])^(a[123] & b[101])^(a[122] & b[102])^(a[121] & b[103])^(a[120] & b[104])^(a[119] & b[105])^(a[118] & b[106])^(a[117] & b[107])^(a[116] & b[108])^(a[115] & b[109])^(a[114] & b[110])^(a[113] & b[111])^(a[112] & b[112])^(a[111] & b[113])^(a[110] & b[114])^(a[109] & b[115])^(a[108] & b[116])^(a[107] & b[117])^(a[106] & b[118])^(a[105] & b[119])^(a[104] & b[120])^(a[103] & b[121])^(a[102] & b[122])^(a[101] & b[123])^(a[100] & b[124])^(a[99] & b[125])^(a[98] & b[126])^(a[97] & b[127])^(a[96] & b[128])^(a[95] & b[129])^(a[94] & b[130])^(a[93] & b[131])^(a[92] & b[132])^(a[91] & b[133])^(a[90] & b[134])^(a[89] & b[135])^(a[88] & b[136])^(a[87] & b[137])^(a[86] & b[138])^(a[85] & b[139])^(a[84] & b[140])^(a[83] & b[141])^(a[82] & b[142])^(a[81] & b[143])^(a[80] & b[144])^(a[79] & b[145])^(a[78] & b[146])^(a[77] & b[147])^(a[76] & b[148])^(a[75] & b[149])^(a[74] & b[150])^(a[73] & b[151])^(a[72] & b[152])^(a[71] & b[153])^(a[70] & b[154])^(a[69] & b[155])^(a[68] & b[156])^(a[67] & b[157])^(a[66] & b[158])^(a[65] & b[159])^(a[64] & b[160])^(a[63] & b[161])^(a[62] & b[162])^(a[61] & b[163])^(a[60] & b[164])^(a[59] & b[165])^(a[58] & b[166])^(a[57] & b[167])^(a[56] & b[168])^(a[55] & b[169])^(a[54] & b[170])^(a[53] & b[171])^(a[52] & b[172])^(a[51] & b[173])^(a[50] & b[174])^(a[49] & b[175])^(a[48] & b[176])^(a[47] & b[177])^(a[46] & b[178])^(a[45] & b[179])^(a[44] & b[180])^(a[43] & b[181])^(a[42] & b[182])^(a[41] & b[183])^(a[40] & b[184])^(a[39] & b[185])^(a[38] & b[186])^(a[37] & b[187])^(a[36] & b[188])^(a[35] & b[189])^(a[34] & b[190])^(a[33] & b[191])^(a[32] & b[192])^(a[31] & b[193])^(a[30] & b[194])^(a[29] & b[195])^(a[28] & b[196])^(a[27] & b[197])^(a[26] & b[198])^(a[25] & b[199])^(a[24] & b[200])^(a[23] & b[201])^(a[22] & b[202])^(a[21] & b[203])^(a[20] & b[204])^(a[19] & b[205])^(a[18] & b[206])^(a[17] & b[207])^(a[16] & b[208])^(a[15] & b[209])^(a[14] & b[210])^(a[13] & b[211])^(a[12] & b[212])^(a[11] & b[213])^(a[10] & b[214])^(a[9] & b[215])^(a[8] & b[216])^(a[7] & b[217])^(a[6] & b[218])^(a[5] & b[219])^(a[4] & b[220])^(a[3] & b[221])^(a[2] & b[222])^(a[1] & b[223])^(a[0] & b[224]);
assign y[225] = (a[225] & b[0])^(a[224] & b[1])^(a[223] & b[2])^(a[222] & b[3])^(a[221] & b[4])^(a[220] & b[5])^(a[219] & b[6])^(a[218] & b[7])^(a[217] & b[8])^(a[216] & b[9])^(a[215] & b[10])^(a[214] & b[11])^(a[213] & b[12])^(a[212] & b[13])^(a[211] & b[14])^(a[210] & b[15])^(a[209] & b[16])^(a[208] & b[17])^(a[207] & b[18])^(a[206] & b[19])^(a[205] & b[20])^(a[204] & b[21])^(a[203] & b[22])^(a[202] & b[23])^(a[201] & b[24])^(a[200] & b[25])^(a[199] & b[26])^(a[198] & b[27])^(a[197] & b[28])^(a[196] & b[29])^(a[195] & b[30])^(a[194] & b[31])^(a[193] & b[32])^(a[192] & b[33])^(a[191] & b[34])^(a[190] & b[35])^(a[189] & b[36])^(a[188] & b[37])^(a[187] & b[38])^(a[186] & b[39])^(a[185] & b[40])^(a[184] & b[41])^(a[183] & b[42])^(a[182] & b[43])^(a[181] & b[44])^(a[180] & b[45])^(a[179] & b[46])^(a[178] & b[47])^(a[177] & b[48])^(a[176] & b[49])^(a[175] & b[50])^(a[174] & b[51])^(a[173] & b[52])^(a[172] & b[53])^(a[171] & b[54])^(a[170] & b[55])^(a[169] & b[56])^(a[168] & b[57])^(a[167] & b[58])^(a[166] & b[59])^(a[165] & b[60])^(a[164] & b[61])^(a[163] & b[62])^(a[162] & b[63])^(a[161] & b[64])^(a[160] & b[65])^(a[159] & b[66])^(a[158] & b[67])^(a[157] & b[68])^(a[156] & b[69])^(a[155] & b[70])^(a[154] & b[71])^(a[153] & b[72])^(a[152] & b[73])^(a[151] & b[74])^(a[150] & b[75])^(a[149] & b[76])^(a[148] & b[77])^(a[147] & b[78])^(a[146] & b[79])^(a[145] & b[80])^(a[144] & b[81])^(a[143] & b[82])^(a[142] & b[83])^(a[141] & b[84])^(a[140] & b[85])^(a[139] & b[86])^(a[138] & b[87])^(a[137] & b[88])^(a[136] & b[89])^(a[135] & b[90])^(a[134] & b[91])^(a[133] & b[92])^(a[132] & b[93])^(a[131] & b[94])^(a[130] & b[95])^(a[129] & b[96])^(a[128] & b[97])^(a[127] & b[98])^(a[126] & b[99])^(a[125] & b[100])^(a[124] & b[101])^(a[123] & b[102])^(a[122] & b[103])^(a[121] & b[104])^(a[120] & b[105])^(a[119] & b[106])^(a[118] & b[107])^(a[117] & b[108])^(a[116] & b[109])^(a[115] & b[110])^(a[114] & b[111])^(a[113] & b[112])^(a[112] & b[113])^(a[111] & b[114])^(a[110] & b[115])^(a[109] & b[116])^(a[108] & b[117])^(a[107] & b[118])^(a[106] & b[119])^(a[105] & b[120])^(a[104] & b[121])^(a[103] & b[122])^(a[102] & b[123])^(a[101] & b[124])^(a[100] & b[125])^(a[99] & b[126])^(a[98] & b[127])^(a[97] & b[128])^(a[96] & b[129])^(a[95] & b[130])^(a[94] & b[131])^(a[93] & b[132])^(a[92] & b[133])^(a[91] & b[134])^(a[90] & b[135])^(a[89] & b[136])^(a[88] & b[137])^(a[87] & b[138])^(a[86] & b[139])^(a[85] & b[140])^(a[84] & b[141])^(a[83] & b[142])^(a[82] & b[143])^(a[81] & b[144])^(a[80] & b[145])^(a[79] & b[146])^(a[78] & b[147])^(a[77] & b[148])^(a[76] & b[149])^(a[75] & b[150])^(a[74] & b[151])^(a[73] & b[152])^(a[72] & b[153])^(a[71] & b[154])^(a[70] & b[155])^(a[69] & b[156])^(a[68] & b[157])^(a[67] & b[158])^(a[66] & b[159])^(a[65] & b[160])^(a[64] & b[161])^(a[63] & b[162])^(a[62] & b[163])^(a[61] & b[164])^(a[60] & b[165])^(a[59] & b[166])^(a[58] & b[167])^(a[57] & b[168])^(a[56] & b[169])^(a[55] & b[170])^(a[54] & b[171])^(a[53] & b[172])^(a[52] & b[173])^(a[51] & b[174])^(a[50] & b[175])^(a[49] & b[176])^(a[48] & b[177])^(a[47] & b[178])^(a[46] & b[179])^(a[45] & b[180])^(a[44] & b[181])^(a[43] & b[182])^(a[42] & b[183])^(a[41] & b[184])^(a[40] & b[185])^(a[39] & b[186])^(a[38] & b[187])^(a[37] & b[188])^(a[36] & b[189])^(a[35] & b[190])^(a[34] & b[191])^(a[33] & b[192])^(a[32] & b[193])^(a[31] & b[194])^(a[30] & b[195])^(a[29] & b[196])^(a[28] & b[197])^(a[27] & b[198])^(a[26] & b[199])^(a[25] & b[200])^(a[24] & b[201])^(a[23] & b[202])^(a[22] & b[203])^(a[21] & b[204])^(a[20] & b[205])^(a[19] & b[206])^(a[18] & b[207])^(a[17] & b[208])^(a[16] & b[209])^(a[15] & b[210])^(a[14] & b[211])^(a[13] & b[212])^(a[12] & b[213])^(a[11] & b[214])^(a[10] & b[215])^(a[9] & b[216])^(a[8] & b[217])^(a[7] & b[218])^(a[6] & b[219])^(a[5] & b[220])^(a[4] & b[221])^(a[3] & b[222])^(a[2] & b[223])^(a[1] & b[224])^(a[0] & b[225]);
assign y[226] = (a[226] & b[0])^(a[225] & b[1])^(a[224] & b[2])^(a[223] & b[3])^(a[222] & b[4])^(a[221] & b[5])^(a[220] & b[6])^(a[219] & b[7])^(a[218] & b[8])^(a[217] & b[9])^(a[216] & b[10])^(a[215] & b[11])^(a[214] & b[12])^(a[213] & b[13])^(a[212] & b[14])^(a[211] & b[15])^(a[210] & b[16])^(a[209] & b[17])^(a[208] & b[18])^(a[207] & b[19])^(a[206] & b[20])^(a[205] & b[21])^(a[204] & b[22])^(a[203] & b[23])^(a[202] & b[24])^(a[201] & b[25])^(a[200] & b[26])^(a[199] & b[27])^(a[198] & b[28])^(a[197] & b[29])^(a[196] & b[30])^(a[195] & b[31])^(a[194] & b[32])^(a[193] & b[33])^(a[192] & b[34])^(a[191] & b[35])^(a[190] & b[36])^(a[189] & b[37])^(a[188] & b[38])^(a[187] & b[39])^(a[186] & b[40])^(a[185] & b[41])^(a[184] & b[42])^(a[183] & b[43])^(a[182] & b[44])^(a[181] & b[45])^(a[180] & b[46])^(a[179] & b[47])^(a[178] & b[48])^(a[177] & b[49])^(a[176] & b[50])^(a[175] & b[51])^(a[174] & b[52])^(a[173] & b[53])^(a[172] & b[54])^(a[171] & b[55])^(a[170] & b[56])^(a[169] & b[57])^(a[168] & b[58])^(a[167] & b[59])^(a[166] & b[60])^(a[165] & b[61])^(a[164] & b[62])^(a[163] & b[63])^(a[162] & b[64])^(a[161] & b[65])^(a[160] & b[66])^(a[159] & b[67])^(a[158] & b[68])^(a[157] & b[69])^(a[156] & b[70])^(a[155] & b[71])^(a[154] & b[72])^(a[153] & b[73])^(a[152] & b[74])^(a[151] & b[75])^(a[150] & b[76])^(a[149] & b[77])^(a[148] & b[78])^(a[147] & b[79])^(a[146] & b[80])^(a[145] & b[81])^(a[144] & b[82])^(a[143] & b[83])^(a[142] & b[84])^(a[141] & b[85])^(a[140] & b[86])^(a[139] & b[87])^(a[138] & b[88])^(a[137] & b[89])^(a[136] & b[90])^(a[135] & b[91])^(a[134] & b[92])^(a[133] & b[93])^(a[132] & b[94])^(a[131] & b[95])^(a[130] & b[96])^(a[129] & b[97])^(a[128] & b[98])^(a[127] & b[99])^(a[126] & b[100])^(a[125] & b[101])^(a[124] & b[102])^(a[123] & b[103])^(a[122] & b[104])^(a[121] & b[105])^(a[120] & b[106])^(a[119] & b[107])^(a[118] & b[108])^(a[117] & b[109])^(a[116] & b[110])^(a[115] & b[111])^(a[114] & b[112])^(a[113] & b[113])^(a[112] & b[114])^(a[111] & b[115])^(a[110] & b[116])^(a[109] & b[117])^(a[108] & b[118])^(a[107] & b[119])^(a[106] & b[120])^(a[105] & b[121])^(a[104] & b[122])^(a[103] & b[123])^(a[102] & b[124])^(a[101] & b[125])^(a[100] & b[126])^(a[99] & b[127])^(a[98] & b[128])^(a[97] & b[129])^(a[96] & b[130])^(a[95] & b[131])^(a[94] & b[132])^(a[93] & b[133])^(a[92] & b[134])^(a[91] & b[135])^(a[90] & b[136])^(a[89] & b[137])^(a[88] & b[138])^(a[87] & b[139])^(a[86] & b[140])^(a[85] & b[141])^(a[84] & b[142])^(a[83] & b[143])^(a[82] & b[144])^(a[81] & b[145])^(a[80] & b[146])^(a[79] & b[147])^(a[78] & b[148])^(a[77] & b[149])^(a[76] & b[150])^(a[75] & b[151])^(a[74] & b[152])^(a[73] & b[153])^(a[72] & b[154])^(a[71] & b[155])^(a[70] & b[156])^(a[69] & b[157])^(a[68] & b[158])^(a[67] & b[159])^(a[66] & b[160])^(a[65] & b[161])^(a[64] & b[162])^(a[63] & b[163])^(a[62] & b[164])^(a[61] & b[165])^(a[60] & b[166])^(a[59] & b[167])^(a[58] & b[168])^(a[57] & b[169])^(a[56] & b[170])^(a[55] & b[171])^(a[54] & b[172])^(a[53] & b[173])^(a[52] & b[174])^(a[51] & b[175])^(a[50] & b[176])^(a[49] & b[177])^(a[48] & b[178])^(a[47] & b[179])^(a[46] & b[180])^(a[45] & b[181])^(a[44] & b[182])^(a[43] & b[183])^(a[42] & b[184])^(a[41] & b[185])^(a[40] & b[186])^(a[39] & b[187])^(a[38] & b[188])^(a[37] & b[189])^(a[36] & b[190])^(a[35] & b[191])^(a[34] & b[192])^(a[33] & b[193])^(a[32] & b[194])^(a[31] & b[195])^(a[30] & b[196])^(a[29] & b[197])^(a[28] & b[198])^(a[27] & b[199])^(a[26] & b[200])^(a[25] & b[201])^(a[24] & b[202])^(a[23] & b[203])^(a[22] & b[204])^(a[21] & b[205])^(a[20] & b[206])^(a[19] & b[207])^(a[18] & b[208])^(a[17] & b[209])^(a[16] & b[210])^(a[15] & b[211])^(a[14] & b[212])^(a[13] & b[213])^(a[12] & b[214])^(a[11] & b[215])^(a[10] & b[216])^(a[9] & b[217])^(a[8] & b[218])^(a[7] & b[219])^(a[6] & b[220])^(a[5] & b[221])^(a[4] & b[222])^(a[3] & b[223])^(a[2] & b[224])^(a[1] & b[225])^(a[0] & b[226]);
assign y[227] = (a[227] & b[0])^(a[226] & b[1])^(a[225] & b[2])^(a[224] & b[3])^(a[223] & b[4])^(a[222] & b[5])^(a[221] & b[6])^(a[220] & b[7])^(a[219] & b[8])^(a[218] & b[9])^(a[217] & b[10])^(a[216] & b[11])^(a[215] & b[12])^(a[214] & b[13])^(a[213] & b[14])^(a[212] & b[15])^(a[211] & b[16])^(a[210] & b[17])^(a[209] & b[18])^(a[208] & b[19])^(a[207] & b[20])^(a[206] & b[21])^(a[205] & b[22])^(a[204] & b[23])^(a[203] & b[24])^(a[202] & b[25])^(a[201] & b[26])^(a[200] & b[27])^(a[199] & b[28])^(a[198] & b[29])^(a[197] & b[30])^(a[196] & b[31])^(a[195] & b[32])^(a[194] & b[33])^(a[193] & b[34])^(a[192] & b[35])^(a[191] & b[36])^(a[190] & b[37])^(a[189] & b[38])^(a[188] & b[39])^(a[187] & b[40])^(a[186] & b[41])^(a[185] & b[42])^(a[184] & b[43])^(a[183] & b[44])^(a[182] & b[45])^(a[181] & b[46])^(a[180] & b[47])^(a[179] & b[48])^(a[178] & b[49])^(a[177] & b[50])^(a[176] & b[51])^(a[175] & b[52])^(a[174] & b[53])^(a[173] & b[54])^(a[172] & b[55])^(a[171] & b[56])^(a[170] & b[57])^(a[169] & b[58])^(a[168] & b[59])^(a[167] & b[60])^(a[166] & b[61])^(a[165] & b[62])^(a[164] & b[63])^(a[163] & b[64])^(a[162] & b[65])^(a[161] & b[66])^(a[160] & b[67])^(a[159] & b[68])^(a[158] & b[69])^(a[157] & b[70])^(a[156] & b[71])^(a[155] & b[72])^(a[154] & b[73])^(a[153] & b[74])^(a[152] & b[75])^(a[151] & b[76])^(a[150] & b[77])^(a[149] & b[78])^(a[148] & b[79])^(a[147] & b[80])^(a[146] & b[81])^(a[145] & b[82])^(a[144] & b[83])^(a[143] & b[84])^(a[142] & b[85])^(a[141] & b[86])^(a[140] & b[87])^(a[139] & b[88])^(a[138] & b[89])^(a[137] & b[90])^(a[136] & b[91])^(a[135] & b[92])^(a[134] & b[93])^(a[133] & b[94])^(a[132] & b[95])^(a[131] & b[96])^(a[130] & b[97])^(a[129] & b[98])^(a[128] & b[99])^(a[127] & b[100])^(a[126] & b[101])^(a[125] & b[102])^(a[124] & b[103])^(a[123] & b[104])^(a[122] & b[105])^(a[121] & b[106])^(a[120] & b[107])^(a[119] & b[108])^(a[118] & b[109])^(a[117] & b[110])^(a[116] & b[111])^(a[115] & b[112])^(a[114] & b[113])^(a[113] & b[114])^(a[112] & b[115])^(a[111] & b[116])^(a[110] & b[117])^(a[109] & b[118])^(a[108] & b[119])^(a[107] & b[120])^(a[106] & b[121])^(a[105] & b[122])^(a[104] & b[123])^(a[103] & b[124])^(a[102] & b[125])^(a[101] & b[126])^(a[100] & b[127])^(a[99] & b[128])^(a[98] & b[129])^(a[97] & b[130])^(a[96] & b[131])^(a[95] & b[132])^(a[94] & b[133])^(a[93] & b[134])^(a[92] & b[135])^(a[91] & b[136])^(a[90] & b[137])^(a[89] & b[138])^(a[88] & b[139])^(a[87] & b[140])^(a[86] & b[141])^(a[85] & b[142])^(a[84] & b[143])^(a[83] & b[144])^(a[82] & b[145])^(a[81] & b[146])^(a[80] & b[147])^(a[79] & b[148])^(a[78] & b[149])^(a[77] & b[150])^(a[76] & b[151])^(a[75] & b[152])^(a[74] & b[153])^(a[73] & b[154])^(a[72] & b[155])^(a[71] & b[156])^(a[70] & b[157])^(a[69] & b[158])^(a[68] & b[159])^(a[67] & b[160])^(a[66] & b[161])^(a[65] & b[162])^(a[64] & b[163])^(a[63] & b[164])^(a[62] & b[165])^(a[61] & b[166])^(a[60] & b[167])^(a[59] & b[168])^(a[58] & b[169])^(a[57] & b[170])^(a[56] & b[171])^(a[55] & b[172])^(a[54] & b[173])^(a[53] & b[174])^(a[52] & b[175])^(a[51] & b[176])^(a[50] & b[177])^(a[49] & b[178])^(a[48] & b[179])^(a[47] & b[180])^(a[46] & b[181])^(a[45] & b[182])^(a[44] & b[183])^(a[43] & b[184])^(a[42] & b[185])^(a[41] & b[186])^(a[40] & b[187])^(a[39] & b[188])^(a[38] & b[189])^(a[37] & b[190])^(a[36] & b[191])^(a[35] & b[192])^(a[34] & b[193])^(a[33] & b[194])^(a[32] & b[195])^(a[31] & b[196])^(a[30] & b[197])^(a[29] & b[198])^(a[28] & b[199])^(a[27] & b[200])^(a[26] & b[201])^(a[25] & b[202])^(a[24] & b[203])^(a[23] & b[204])^(a[22] & b[205])^(a[21] & b[206])^(a[20] & b[207])^(a[19] & b[208])^(a[18] & b[209])^(a[17] & b[210])^(a[16] & b[211])^(a[15] & b[212])^(a[14] & b[213])^(a[13] & b[214])^(a[12] & b[215])^(a[11] & b[216])^(a[10] & b[217])^(a[9] & b[218])^(a[8] & b[219])^(a[7] & b[220])^(a[6] & b[221])^(a[5] & b[222])^(a[4] & b[223])^(a[3] & b[224])^(a[2] & b[225])^(a[1] & b[226])^(a[0] & b[227]);
assign y[228] = (a[228] & b[0])^(a[227] & b[1])^(a[226] & b[2])^(a[225] & b[3])^(a[224] & b[4])^(a[223] & b[5])^(a[222] & b[6])^(a[221] & b[7])^(a[220] & b[8])^(a[219] & b[9])^(a[218] & b[10])^(a[217] & b[11])^(a[216] & b[12])^(a[215] & b[13])^(a[214] & b[14])^(a[213] & b[15])^(a[212] & b[16])^(a[211] & b[17])^(a[210] & b[18])^(a[209] & b[19])^(a[208] & b[20])^(a[207] & b[21])^(a[206] & b[22])^(a[205] & b[23])^(a[204] & b[24])^(a[203] & b[25])^(a[202] & b[26])^(a[201] & b[27])^(a[200] & b[28])^(a[199] & b[29])^(a[198] & b[30])^(a[197] & b[31])^(a[196] & b[32])^(a[195] & b[33])^(a[194] & b[34])^(a[193] & b[35])^(a[192] & b[36])^(a[191] & b[37])^(a[190] & b[38])^(a[189] & b[39])^(a[188] & b[40])^(a[187] & b[41])^(a[186] & b[42])^(a[185] & b[43])^(a[184] & b[44])^(a[183] & b[45])^(a[182] & b[46])^(a[181] & b[47])^(a[180] & b[48])^(a[179] & b[49])^(a[178] & b[50])^(a[177] & b[51])^(a[176] & b[52])^(a[175] & b[53])^(a[174] & b[54])^(a[173] & b[55])^(a[172] & b[56])^(a[171] & b[57])^(a[170] & b[58])^(a[169] & b[59])^(a[168] & b[60])^(a[167] & b[61])^(a[166] & b[62])^(a[165] & b[63])^(a[164] & b[64])^(a[163] & b[65])^(a[162] & b[66])^(a[161] & b[67])^(a[160] & b[68])^(a[159] & b[69])^(a[158] & b[70])^(a[157] & b[71])^(a[156] & b[72])^(a[155] & b[73])^(a[154] & b[74])^(a[153] & b[75])^(a[152] & b[76])^(a[151] & b[77])^(a[150] & b[78])^(a[149] & b[79])^(a[148] & b[80])^(a[147] & b[81])^(a[146] & b[82])^(a[145] & b[83])^(a[144] & b[84])^(a[143] & b[85])^(a[142] & b[86])^(a[141] & b[87])^(a[140] & b[88])^(a[139] & b[89])^(a[138] & b[90])^(a[137] & b[91])^(a[136] & b[92])^(a[135] & b[93])^(a[134] & b[94])^(a[133] & b[95])^(a[132] & b[96])^(a[131] & b[97])^(a[130] & b[98])^(a[129] & b[99])^(a[128] & b[100])^(a[127] & b[101])^(a[126] & b[102])^(a[125] & b[103])^(a[124] & b[104])^(a[123] & b[105])^(a[122] & b[106])^(a[121] & b[107])^(a[120] & b[108])^(a[119] & b[109])^(a[118] & b[110])^(a[117] & b[111])^(a[116] & b[112])^(a[115] & b[113])^(a[114] & b[114])^(a[113] & b[115])^(a[112] & b[116])^(a[111] & b[117])^(a[110] & b[118])^(a[109] & b[119])^(a[108] & b[120])^(a[107] & b[121])^(a[106] & b[122])^(a[105] & b[123])^(a[104] & b[124])^(a[103] & b[125])^(a[102] & b[126])^(a[101] & b[127])^(a[100] & b[128])^(a[99] & b[129])^(a[98] & b[130])^(a[97] & b[131])^(a[96] & b[132])^(a[95] & b[133])^(a[94] & b[134])^(a[93] & b[135])^(a[92] & b[136])^(a[91] & b[137])^(a[90] & b[138])^(a[89] & b[139])^(a[88] & b[140])^(a[87] & b[141])^(a[86] & b[142])^(a[85] & b[143])^(a[84] & b[144])^(a[83] & b[145])^(a[82] & b[146])^(a[81] & b[147])^(a[80] & b[148])^(a[79] & b[149])^(a[78] & b[150])^(a[77] & b[151])^(a[76] & b[152])^(a[75] & b[153])^(a[74] & b[154])^(a[73] & b[155])^(a[72] & b[156])^(a[71] & b[157])^(a[70] & b[158])^(a[69] & b[159])^(a[68] & b[160])^(a[67] & b[161])^(a[66] & b[162])^(a[65] & b[163])^(a[64] & b[164])^(a[63] & b[165])^(a[62] & b[166])^(a[61] & b[167])^(a[60] & b[168])^(a[59] & b[169])^(a[58] & b[170])^(a[57] & b[171])^(a[56] & b[172])^(a[55] & b[173])^(a[54] & b[174])^(a[53] & b[175])^(a[52] & b[176])^(a[51] & b[177])^(a[50] & b[178])^(a[49] & b[179])^(a[48] & b[180])^(a[47] & b[181])^(a[46] & b[182])^(a[45] & b[183])^(a[44] & b[184])^(a[43] & b[185])^(a[42] & b[186])^(a[41] & b[187])^(a[40] & b[188])^(a[39] & b[189])^(a[38] & b[190])^(a[37] & b[191])^(a[36] & b[192])^(a[35] & b[193])^(a[34] & b[194])^(a[33] & b[195])^(a[32] & b[196])^(a[31] & b[197])^(a[30] & b[198])^(a[29] & b[199])^(a[28] & b[200])^(a[27] & b[201])^(a[26] & b[202])^(a[25] & b[203])^(a[24] & b[204])^(a[23] & b[205])^(a[22] & b[206])^(a[21] & b[207])^(a[20] & b[208])^(a[19] & b[209])^(a[18] & b[210])^(a[17] & b[211])^(a[16] & b[212])^(a[15] & b[213])^(a[14] & b[214])^(a[13] & b[215])^(a[12] & b[216])^(a[11] & b[217])^(a[10] & b[218])^(a[9] & b[219])^(a[8] & b[220])^(a[7] & b[221])^(a[6] & b[222])^(a[5] & b[223])^(a[4] & b[224])^(a[3] & b[225])^(a[2] & b[226])^(a[1] & b[227])^(a[0] & b[228]);
assign y[229] = (a[229] & b[0])^(a[228] & b[1])^(a[227] & b[2])^(a[226] & b[3])^(a[225] & b[4])^(a[224] & b[5])^(a[223] & b[6])^(a[222] & b[7])^(a[221] & b[8])^(a[220] & b[9])^(a[219] & b[10])^(a[218] & b[11])^(a[217] & b[12])^(a[216] & b[13])^(a[215] & b[14])^(a[214] & b[15])^(a[213] & b[16])^(a[212] & b[17])^(a[211] & b[18])^(a[210] & b[19])^(a[209] & b[20])^(a[208] & b[21])^(a[207] & b[22])^(a[206] & b[23])^(a[205] & b[24])^(a[204] & b[25])^(a[203] & b[26])^(a[202] & b[27])^(a[201] & b[28])^(a[200] & b[29])^(a[199] & b[30])^(a[198] & b[31])^(a[197] & b[32])^(a[196] & b[33])^(a[195] & b[34])^(a[194] & b[35])^(a[193] & b[36])^(a[192] & b[37])^(a[191] & b[38])^(a[190] & b[39])^(a[189] & b[40])^(a[188] & b[41])^(a[187] & b[42])^(a[186] & b[43])^(a[185] & b[44])^(a[184] & b[45])^(a[183] & b[46])^(a[182] & b[47])^(a[181] & b[48])^(a[180] & b[49])^(a[179] & b[50])^(a[178] & b[51])^(a[177] & b[52])^(a[176] & b[53])^(a[175] & b[54])^(a[174] & b[55])^(a[173] & b[56])^(a[172] & b[57])^(a[171] & b[58])^(a[170] & b[59])^(a[169] & b[60])^(a[168] & b[61])^(a[167] & b[62])^(a[166] & b[63])^(a[165] & b[64])^(a[164] & b[65])^(a[163] & b[66])^(a[162] & b[67])^(a[161] & b[68])^(a[160] & b[69])^(a[159] & b[70])^(a[158] & b[71])^(a[157] & b[72])^(a[156] & b[73])^(a[155] & b[74])^(a[154] & b[75])^(a[153] & b[76])^(a[152] & b[77])^(a[151] & b[78])^(a[150] & b[79])^(a[149] & b[80])^(a[148] & b[81])^(a[147] & b[82])^(a[146] & b[83])^(a[145] & b[84])^(a[144] & b[85])^(a[143] & b[86])^(a[142] & b[87])^(a[141] & b[88])^(a[140] & b[89])^(a[139] & b[90])^(a[138] & b[91])^(a[137] & b[92])^(a[136] & b[93])^(a[135] & b[94])^(a[134] & b[95])^(a[133] & b[96])^(a[132] & b[97])^(a[131] & b[98])^(a[130] & b[99])^(a[129] & b[100])^(a[128] & b[101])^(a[127] & b[102])^(a[126] & b[103])^(a[125] & b[104])^(a[124] & b[105])^(a[123] & b[106])^(a[122] & b[107])^(a[121] & b[108])^(a[120] & b[109])^(a[119] & b[110])^(a[118] & b[111])^(a[117] & b[112])^(a[116] & b[113])^(a[115] & b[114])^(a[114] & b[115])^(a[113] & b[116])^(a[112] & b[117])^(a[111] & b[118])^(a[110] & b[119])^(a[109] & b[120])^(a[108] & b[121])^(a[107] & b[122])^(a[106] & b[123])^(a[105] & b[124])^(a[104] & b[125])^(a[103] & b[126])^(a[102] & b[127])^(a[101] & b[128])^(a[100] & b[129])^(a[99] & b[130])^(a[98] & b[131])^(a[97] & b[132])^(a[96] & b[133])^(a[95] & b[134])^(a[94] & b[135])^(a[93] & b[136])^(a[92] & b[137])^(a[91] & b[138])^(a[90] & b[139])^(a[89] & b[140])^(a[88] & b[141])^(a[87] & b[142])^(a[86] & b[143])^(a[85] & b[144])^(a[84] & b[145])^(a[83] & b[146])^(a[82] & b[147])^(a[81] & b[148])^(a[80] & b[149])^(a[79] & b[150])^(a[78] & b[151])^(a[77] & b[152])^(a[76] & b[153])^(a[75] & b[154])^(a[74] & b[155])^(a[73] & b[156])^(a[72] & b[157])^(a[71] & b[158])^(a[70] & b[159])^(a[69] & b[160])^(a[68] & b[161])^(a[67] & b[162])^(a[66] & b[163])^(a[65] & b[164])^(a[64] & b[165])^(a[63] & b[166])^(a[62] & b[167])^(a[61] & b[168])^(a[60] & b[169])^(a[59] & b[170])^(a[58] & b[171])^(a[57] & b[172])^(a[56] & b[173])^(a[55] & b[174])^(a[54] & b[175])^(a[53] & b[176])^(a[52] & b[177])^(a[51] & b[178])^(a[50] & b[179])^(a[49] & b[180])^(a[48] & b[181])^(a[47] & b[182])^(a[46] & b[183])^(a[45] & b[184])^(a[44] & b[185])^(a[43] & b[186])^(a[42] & b[187])^(a[41] & b[188])^(a[40] & b[189])^(a[39] & b[190])^(a[38] & b[191])^(a[37] & b[192])^(a[36] & b[193])^(a[35] & b[194])^(a[34] & b[195])^(a[33] & b[196])^(a[32] & b[197])^(a[31] & b[198])^(a[30] & b[199])^(a[29] & b[200])^(a[28] & b[201])^(a[27] & b[202])^(a[26] & b[203])^(a[25] & b[204])^(a[24] & b[205])^(a[23] & b[206])^(a[22] & b[207])^(a[21] & b[208])^(a[20] & b[209])^(a[19] & b[210])^(a[18] & b[211])^(a[17] & b[212])^(a[16] & b[213])^(a[15] & b[214])^(a[14] & b[215])^(a[13] & b[216])^(a[12] & b[217])^(a[11] & b[218])^(a[10] & b[219])^(a[9] & b[220])^(a[8] & b[221])^(a[7] & b[222])^(a[6] & b[223])^(a[5] & b[224])^(a[4] & b[225])^(a[3] & b[226])^(a[2] & b[227])^(a[1] & b[228])^(a[0] & b[229]);
assign y[230] = (a[230] & b[0])^(a[229] & b[1])^(a[228] & b[2])^(a[227] & b[3])^(a[226] & b[4])^(a[225] & b[5])^(a[224] & b[6])^(a[223] & b[7])^(a[222] & b[8])^(a[221] & b[9])^(a[220] & b[10])^(a[219] & b[11])^(a[218] & b[12])^(a[217] & b[13])^(a[216] & b[14])^(a[215] & b[15])^(a[214] & b[16])^(a[213] & b[17])^(a[212] & b[18])^(a[211] & b[19])^(a[210] & b[20])^(a[209] & b[21])^(a[208] & b[22])^(a[207] & b[23])^(a[206] & b[24])^(a[205] & b[25])^(a[204] & b[26])^(a[203] & b[27])^(a[202] & b[28])^(a[201] & b[29])^(a[200] & b[30])^(a[199] & b[31])^(a[198] & b[32])^(a[197] & b[33])^(a[196] & b[34])^(a[195] & b[35])^(a[194] & b[36])^(a[193] & b[37])^(a[192] & b[38])^(a[191] & b[39])^(a[190] & b[40])^(a[189] & b[41])^(a[188] & b[42])^(a[187] & b[43])^(a[186] & b[44])^(a[185] & b[45])^(a[184] & b[46])^(a[183] & b[47])^(a[182] & b[48])^(a[181] & b[49])^(a[180] & b[50])^(a[179] & b[51])^(a[178] & b[52])^(a[177] & b[53])^(a[176] & b[54])^(a[175] & b[55])^(a[174] & b[56])^(a[173] & b[57])^(a[172] & b[58])^(a[171] & b[59])^(a[170] & b[60])^(a[169] & b[61])^(a[168] & b[62])^(a[167] & b[63])^(a[166] & b[64])^(a[165] & b[65])^(a[164] & b[66])^(a[163] & b[67])^(a[162] & b[68])^(a[161] & b[69])^(a[160] & b[70])^(a[159] & b[71])^(a[158] & b[72])^(a[157] & b[73])^(a[156] & b[74])^(a[155] & b[75])^(a[154] & b[76])^(a[153] & b[77])^(a[152] & b[78])^(a[151] & b[79])^(a[150] & b[80])^(a[149] & b[81])^(a[148] & b[82])^(a[147] & b[83])^(a[146] & b[84])^(a[145] & b[85])^(a[144] & b[86])^(a[143] & b[87])^(a[142] & b[88])^(a[141] & b[89])^(a[140] & b[90])^(a[139] & b[91])^(a[138] & b[92])^(a[137] & b[93])^(a[136] & b[94])^(a[135] & b[95])^(a[134] & b[96])^(a[133] & b[97])^(a[132] & b[98])^(a[131] & b[99])^(a[130] & b[100])^(a[129] & b[101])^(a[128] & b[102])^(a[127] & b[103])^(a[126] & b[104])^(a[125] & b[105])^(a[124] & b[106])^(a[123] & b[107])^(a[122] & b[108])^(a[121] & b[109])^(a[120] & b[110])^(a[119] & b[111])^(a[118] & b[112])^(a[117] & b[113])^(a[116] & b[114])^(a[115] & b[115])^(a[114] & b[116])^(a[113] & b[117])^(a[112] & b[118])^(a[111] & b[119])^(a[110] & b[120])^(a[109] & b[121])^(a[108] & b[122])^(a[107] & b[123])^(a[106] & b[124])^(a[105] & b[125])^(a[104] & b[126])^(a[103] & b[127])^(a[102] & b[128])^(a[101] & b[129])^(a[100] & b[130])^(a[99] & b[131])^(a[98] & b[132])^(a[97] & b[133])^(a[96] & b[134])^(a[95] & b[135])^(a[94] & b[136])^(a[93] & b[137])^(a[92] & b[138])^(a[91] & b[139])^(a[90] & b[140])^(a[89] & b[141])^(a[88] & b[142])^(a[87] & b[143])^(a[86] & b[144])^(a[85] & b[145])^(a[84] & b[146])^(a[83] & b[147])^(a[82] & b[148])^(a[81] & b[149])^(a[80] & b[150])^(a[79] & b[151])^(a[78] & b[152])^(a[77] & b[153])^(a[76] & b[154])^(a[75] & b[155])^(a[74] & b[156])^(a[73] & b[157])^(a[72] & b[158])^(a[71] & b[159])^(a[70] & b[160])^(a[69] & b[161])^(a[68] & b[162])^(a[67] & b[163])^(a[66] & b[164])^(a[65] & b[165])^(a[64] & b[166])^(a[63] & b[167])^(a[62] & b[168])^(a[61] & b[169])^(a[60] & b[170])^(a[59] & b[171])^(a[58] & b[172])^(a[57] & b[173])^(a[56] & b[174])^(a[55] & b[175])^(a[54] & b[176])^(a[53] & b[177])^(a[52] & b[178])^(a[51] & b[179])^(a[50] & b[180])^(a[49] & b[181])^(a[48] & b[182])^(a[47] & b[183])^(a[46] & b[184])^(a[45] & b[185])^(a[44] & b[186])^(a[43] & b[187])^(a[42] & b[188])^(a[41] & b[189])^(a[40] & b[190])^(a[39] & b[191])^(a[38] & b[192])^(a[37] & b[193])^(a[36] & b[194])^(a[35] & b[195])^(a[34] & b[196])^(a[33] & b[197])^(a[32] & b[198])^(a[31] & b[199])^(a[30] & b[200])^(a[29] & b[201])^(a[28] & b[202])^(a[27] & b[203])^(a[26] & b[204])^(a[25] & b[205])^(a[24] & b[206])^(a[23] & b[207])^(a[22] & b[208])^(a[21] & b[209])^(a[20] & b[210])^(a[19] & b[211])^(a[18] & b[212])^(a[17] & b[213])^(a[16] & b[214])^(a[15] & b[215])^(a[14] & b[216])^(a[13] & b[217])^(a[12] & b[218])^(a[11] & b[219])^(a[10] & b[220])^(a[9] & b[221])^(a[8] & b[222])^(a[7] & b[223])^(a[6] & b[224])^(a[5] & b[225])^(a[4] & b[226])^(a[3] & b[227])^(a[2] & b[228])^(a[1] & b[229])^(a[0] & b[230]);
assign y[231] = (a[231] & b[0])^(a[230] & b[1])^(a[229] & b[2])^(a[228] & b[3])^(a[227] & b[4])^(a[226] & b[5])^(a[225] & b[6])^(a[224] & b[7])^(a[223] & b[8])^(a[222] & b[9])^(a[221] & b[10])^(a[220] & b[11])^(a[219] & b[12])^(a[218] & b[13])^(a[217] & b[14])^(a[216] & b[15])^(a[215] & b[16])^(a[214] & b[17])^(a[213] & b[18])^(a[212] & b[19])^(a[211] & b[20])^(a[210] & b[21])^(a[209] & b[22])^(a[208] & b[23])^(a[207] & b[24])^(a[206] & b[25])^(a[205] & b[26])^(a[204] & b[27])^(a[203] & b[28])^(a[202] & b[29])^(a[201] & b[30])^(a[200] & b[31])^(a[199] & b[32])^(a[198] & b[33])^(a[197] & b[34])^(a[196] & b[35])^(a[195] & b[36])^(a[194] & b[37])^(a[193] & b[38])^(a[192] & b[39])^(a[191] & b[40])^(a[190] & b[41])^(a[189] & b[42])^(a[188] & b[43])^(a[187] & b[44])^(a[186] & b[45])^(a[185] & b[46])^(a[184] & b[47])^(a[183] & b[48])^(a[182] & b[49])^(a[181] & b[50])^(a[180] & b[51])^(a[179] & b[52])^(a[178] & b[53])^(a[177] & b[54])^(a[176] & b[55])^(a[175] & b[56])^(a[174] & b[57])^(a[173] & b[58])^(a[172] & b[59])^(a[171] & b[60])^(a[170] & b[61])^(a[169] & b[62])^(a[168] & b[63])^(a[167] & b[64])^(a[166] & b[65])^(a[165] & b[66])^(a[164] & b[67])^(a[163] & b[68])^(a[162] & b[69])^(a[161] & b[70])^(a[160] & b[71])^(a[159] & b[72])^(a[158] & b[73])^(a[157] & b[74])^(a[156] & b[75])^(a[155] & b[76])^(a[154] & b[77])^(a[153] & b[78])^(a[152] & b[79])^(a[151] & b[80])^(a[150] & b[81])^(a[149] & b[82])^(a[148] & b[83])^(a[147] & b[84])^(a[146] & b[85])^(a[145] & b[86])^(a[144] & b[87])^(a[143] & b[88])^(a[142] & b[89])^(a[141] & b[90])^(a[140] & b[91])^(a[139] & b[92])^(a[138] & b[93])^(a[137] & b[94])^(a[136] & b[95])^(a[135] & b[96])^(a[134] & b[97])^(a[133] & b[98])^(a[132] & b[99])^(a[131] & b[100])^(a[130] & b[101])^(a[129] & b[102])^(a[128] & b[103])^(a[127] & b[104])^(a[126] & b[105])^(a[125] & b[106])^(a[124] & b[107])^(a[123] & b[108])^(a[122] & b[109])^(a[121] & b[110])^(a[120] & b[111])^(a[119] & b[112])^(a[118] & b[113])^(a[117] & b[114])^(a[116] & b[115])^(a[115] & b[116])^(a[114] & b[117])^(a[113] & b[118])^(a[112] & b[119])^(a[111] & b[120])^(a[110] & b[121])^(a[109] & b[122])^(a[108] & b[123])^(a[107] & b[124])^(a[106] & b[125])^(a[105] & b[126])^(a[104] & b[127])^(a[103] & b[128])^(a[102] & b[129])^(a[101] & b[130])^(a[100] & b[131])^(a[99] & b[132])^(a[98] & b[133])^(a[97] & b[134])^(a[96] & b[135])^(a[95] & b[136])^(a[94] & b[137])^(a[93] & b[138])^(a[92] & b[139])^(a[91] & b[140])^(a[90] & b[141])^(a[89] & b[142])^(a[88] & b[143])^(a[87] & b[144])^(a[86] & b[145])^(a[85] & b[146])^(a[84] & b[147])^(a[83] & b[148])^(a[82] & b[149])^(a[81] & b[150])^(a[80] & b[151])^(a[79] & b[152])^(a[78] & b[153])^(a[77] & b[154])^(a[76] & b[155])^(a[75] & b[156])^(a[74] & b[157])^(a[73] & b[158])^(a[72] & b[159])^(a[71] & b[160])^(a[70] & b[161])^(a[69] & b[162])^(a[68] & b[163])^(a[67] & b[164])^(a[66] & b[165])^(a[65] & b[166])^(a[64] & b[167])^(a[63] & b[168])^(a[62] & b[169])^(a[61] & b[170])^(a[60] & b[171])^(a[59] & b[172])^(a[58] & b[173])^(a[57] & b[174])^(a[56] & b[175])^(a[55] & b[176])^(a[54] & b[177])^(a[53] & b[178])^(a[52] & b[179])^(a[51] & b[180])^(a[50] & b[181])^(a[49] & b[182])^(a[48] & b[183])^(a[47] & b[184])^(a[46] & b[185])^(a[45] & b[186])^(a[44] & b[187])^(a[43] & b[188])^(a[42] & b[189])^(a[41] & b[190])^(a[40] & b[191])^(a[39] & b[192])^(a[38] & b[193])^(a[37] & b[194])^(a[36] & b[195])^(a[35] & b[196])^(a[34] & b[197])^(a[33] & b[198])^(a[32] & b[199])^(a[31] & b[200])^(a[30] & b[201])^(a[29] & b[202])^(a[28] & b[203])^(a[27] & b[204])^(a[26] & b[205])^(a[25] & b[206])^(a[24] & b[207])^(a[23] & b[208])^(a[22] & b[209])^(a[21] & b[210])^(a[20] & b[211])^(a[19] & b[212])^(a[18] & b[213])^(a[17] & b[214])^(a[16] & b[215])^(a[15] & b[216])^(a[14] & b[217])^(a[13] & b[218])^(a[12] & b[219])^(a[11] & b[220])^(a[10] & b[221])^(a[9] & b[222])^(a[8] & b[223])^(a[7] & b[224])^(a[6] & b[225])^(a[5] & b[226])^(a[4] & b[227])^(a[3] & b[228])^(a[2] & b[229])^(a[1] & b[230])^(a[0] & b[231]);
assign y[232] = (a[232] & b[0])^(a[231] & b[1])^(a[230] & b[2])^(a[229] & b[3])^(a[228] & b[4])^(a[227] & b[5])^(a[226] & b[6])^(a[225] & b[7])^(a[224] & b[8])^(a[223] & b[9])^(a[222] & b[10])^(a[221] & b[11])^(a[220] & b[12])^(a[219] & b[13])^(a[218] & b[14])^(a[217] & b[15])^(a[216] & b[16])^(a[215] & b[17])^(a[214] & b[18])^(a[213] & b[19])^(a[212] & b[20])^(a[211] & b[21])^(a[210] & b[22])^(a[209] & b[23])^(a[208] & b[24])^(a[207] & b[25])^(a[206] & b[26])^(a[205] & b[27])^(a[204] & b[28])^(a[203] & b[29])^(a[202] & b[30])^(a[201] & b[31])^(a[200] & b[32])^(a[199] & b[33])^(a[198] & b[34])^(a[197] & b[35])^(a[196] & b[36])^(a[195] & b[37])^(a[194] & b[38])^(a[193] & b[39])^(a[192] & b[40])^(a[191] & b[41])^(a[190] & b[42])^(a[189] & b[43])^(a[188] & b[44])^(a[187] & b[45])^(a[186] & b[46])^(a[185] & b[47])^(a[184] & b[48])^(a[183] & b[49])^(a[182] & b[50])^(a[181] & b[51])^(a[180] & b[52])^(a[179] & b[53])^(a[178] & b[54])^(a[177] & b[55])^(a[176] & b[56])^(a[175] & b[57])^(a[174] & b[58])^(a[173] & b[59])^(a[172] & b[60])^(a[171] & b[61])^(a[170] & b[62])^(a[169] & b[63])^(a[168] & b[64])^(a[167] & b[65])^(a[166] & b[66])^(a[165] & b[67])^(a[164] & b[68])^(a[163] & b[69])^(a[162] & b[70])^(a[161] & b[71])^(a[160] & b[72])^(a[159] & b[73])^(a[158] & b[74])^(a[157] & b[75])^(a[156] & b[76])^(a[155] & b[77])^(a[154] & b[78])^(a[153] & b[79])^(a[152] & b[80])^(a[151] & b[81])^(a[150] & b[82])^(a[149] & b[83])^(a[148] & b[84])^(a[147] & b[85])^(a[146] & b[86])^(a[145] & b[87])^(a[144] & b[88])^(a[143] & b[89])^(a[142] & b[90])^(a[141] & b[91])^(a[140] & b[92])^(a[139] & b[93])^(a[138] & b[94])^(a[137] & b[95])^(a[136] & b[96])^(a[135] & b[97])^(a[134] & b[98])^(a[133] & b[99])^(a[132] & b[100])^(a[131] & b[101])^(a[130] & b[102])^(a[129] & b[103])^(a[128] & b[104])^(a[127] & b[105])^(a[126] & b[106])^(a[125] & b[107])^(a[124] & b[108])^(a[123] & b[109])^(a[122] & b[110])^(a[121] & b[111])^(a[120] & b[112])^(a[119] & b[113])^(a[118] & b[114])^(a[117] & b[115])^(a[116] & b[116])^(a[115] & b[117])^(a[114] & b[118])^(a[113] & b[119])^(a[112] & b[120])^(a[111] & b[121])^(a[110] & b[122])^(a[109] & b[123])^(a[108] & b[124])^(a[107] & b[125])^(a[106] & b[126])^(a[105] & b[127])^(a[104] & b[128])^(a[103] & b[129])^(a[102] & b[130])^(a[101] & b[131])^(a[100] & b[132])^(a[99] & b[133])^(a[98] & b[134])^(a[97] & b[135])^(a[96] & b[136])^(a[95] & b[137])^(a[94] & b[138])^(a[93] & b[139])^(a[92] & b[140])^(a[91] & b[141])^(a[90] & b[142])^(a[89] & b[143])^(a[88] & b[144])^(a[87] & b[145])^(a[86] & b[146])^(a[85] & b[147])^(a[84] & b[148])^(a[83] & b[149])^(a[82] & b[150])^(a[81] & b[151])^(a[80] & b[152])^(a[79] & b[153])^(a[78] & b[154])^(a[77] & b[155])^(a[76] & b[156])^(a[75] & b[157])^(a[74] & b[158])^(a[73] & b[159])^(a[72] & b[160])^(a[71] & b[161])^(a[70] & b[162])^(a[69] & b[163])^(a[68] & b[164])^(a[67] & b[165])^(a[66] & b[166])^(a[65] & b[167])^(a[64] & b[168])^(a[63] & b[169])^(a[62] & b[170])^(a[61] & b[171])^(a[60] & b[172])^(a[59] & b[173])^(a[58] & b[174])^(a[57] & b[175])^(a[56] & b[176])^(a[55] & b[177])^(a[54] & b[178])^(a[53] & b[179])^(a[52] & b[180])^(a[51] & b[181])^(a[50] & b[182])^(a[49] & b[183])^(a[48] & b[184])^(a[47] & b[185])^(a[46] & b[186])^(a[45] & b[187])^(a[44] & b[188])^(a[43] & b[189])^(a[42] & b[190])^(a[41] & b[191])^(a[40] & b[192])^(a[39] & b[193])^(a[38] & b[194])^(a[37] & b[195])^(a[36] & b[196])^(a[35] & b[197])^(a[34] & b[198])^(a[33] & b[199])^(a[32] & b[200])^(a[31] & b[201])^(a[30] & b[202])^(a[29] & b[203])^(a[28] & b[204])^(a[27] & b[205])^(a[26] & b[206])^(a[25] & b[207])^(a[24] & b[208])^(a[23] & b[209])^(a[22] & b[210])^(a[21] & b[211])^(a[20] & b[212])^(a[19] & b[213])^(a[18] & b[214])^(a[17] & b[215])^(a[16] & b[216])^(a[15] & b[217])^(a[14] & b[218])^(a[13] & b[219])^(a[12] & b[220])^(a[11] & b[221])^(a[10] & b[222])^(a[9] & b[223])^(a[8] & b[224])^(a[7] & b[225])^(a[6] & b[226])^(a[5] & b[227])^(a[4] & b[228])^(a[3] & b[229])^(a[2] & b[230])^(a[1] & b[231])^(a[0] & b[232]);
assign y[233] = (a[232] & b[1])^(a[231] & b[2])^(a[230] & b[3])^(a[229] & b[4])^(a[228] & b[5])^(a[227] & b[6])^(a[226] & b[7])^(a[225] & b[8])^(a[224] & b[9])^(a[223] & b[10])^(a[222] & b[11])^(a[221] & b[12])^(a[220] & b[13])^(a[219] & b[14])^(a[218] & b[15])^(a[217] & b[16])^(a[216] & b[17])^(a[215] & b[18])^(a[214] & b[19])^(a[213] & b[20])^(a[212] & b[21])^(a[211] & b[22])^(a[210] & b[23])^(a[209] & b[24])^(a[208] & b[25])^(a[207] & b[26])^(a[206] & b[27])^(a[205] & b[28])^(a[204] & b[29])^(a[203] & b[30])^(a[202] & b[31])^(a[201] & b[32])^(a[200] & b[33])^(a[199] & b[34])^(a[198] & b[35])^(a[197] & b[36])^(a[196] & b[37])^(a[195] & b[38])^(a[194] & b[39])^(a[193] & b[40])^(a[192] & b[41])^(a[191] & b[42])^(a[190] & b[43])^(a[189] & b[44])^(a[188] & b[45])^(a[187] & b[46])^(a[186] & b[47])^(a[185] & b[48])^(a[184] & b[49])^(a[183] & b[50])^(a[182] & b[51])^(a[181] & b[52])^(a[180] & b[53])^(a[179] & b[54])^(a[178] & b[55])^(a[177] & b[56])^(a[176] & b[57])^(a[175] & b[58])^(a[174] & b[59])^(a[173] & b[60])^(a[172] & b[61])^(a[171] & b[62])^(a[170] & b[63])^(a[169] & b[64])^(a[168] & b[65])^(a[167] & b[66])^(a[166] & b[67])^(a[165] & b[68])^(a[164] & b[69])^(a[163] & b[70])^(a[162] & b[71])^(a[161] & b[72])^(a[160] & b[73])^(a[159] & b[74])^(a[158] & b[75])^(a[157] & b[76])^(a[156] & b[77])^(a[155] & b[78])^(a[154] & b[79])^(a[153] & b[80])^(a[152] & b[81])^(a[151] & b[82])^(a[150] & b[83])^(a[149] & b[84])^(a[148] & b[85])^(a[147] & b[86])^(a[146] & b[87])^(a[145] & b[88])^(a[144] & b[89])^(a[143] & b[90])^(a[142] & b[91])^(a[141] & b[92])^(a[140] & b[93])^(a[139] & b[94])^(a[138] & b[95])^(a[137] & b[96])^(a[136] & b[97])^(a[135] & b[98])^(a[134] & b[99])^(a[133] & b[100])^(a[132] & b[101])^(a[131] & b[102])^(a[130] & b[103])^(a[129] & b[104])^(a[128] & b[105])^(a[127] & b[106])^(a[126] & b[107])^(a[125] & b[108])^(a[124] & b[109])^(a[123] & b[110])^(a[122] & b[111])^(a[121] & b[112])^(a[120] & b[113])^(a[119] & b[114])^(a[118] & b[115])^(a[117] & b[116])^(a[116] & b[117])^(a[115] & b[118])^(a[114] & b[119])^(a[113] & b[120])^(a[112] & b[121])^(a[111] & b[122])^(a[110] & b[123])^(a[109] & b[124])^(a[108] & b[125])^(a[107] & b[126])^(a[106] & b[127])^(a[105] & b[128])^(a[104] & b[129])^(a[103] & b[130])^(a[102] & b[131])^(a[101] & b[132])^(a[100] & b[133])^(a[99] & b[134])^(a[98] & b[135])^(a[97] & b[136])^(a[96] & b[137])^(a[95] & b[138])^(a[94] & b[139])^(a[93] & b[140])^(a[92] & b[141])^(a[91] & b[142])^(a[90] & b[143])^(a[89] & b[144])^(a[88] & b[145])^(a[87] & b[146])^(a[86] & b[147])^(a[85] & b[148])^(a[84] & b[149])^(a[83] & b[150])^(a[82] & b[151])^(a[81] & b[152])^(a[80] & b[153])^(a[79] & b[154])^(a[78] & b[155])^(a[77] & b[156])^(a[76] & b[157])^(a[75] & b[158])^(a[74] & b[159])^(a[73] & b[160])^(a[72] & b[161])^(a[71] & b[162])^(a[70] & b[163])^(a[69] & b[164])^(a[68] & b[165])^(a[67] & b[166])^(a[66] & b[167])^(a[65] & b[168])^(a[64] & b[169])^(a[63] & b[170])^(a[62] & b[171])^(a[61] & b[172])^(a[60] & b[173])^(a[59] & b[174])^(a[58] & b[175])^(a[57] & b[176])^(a[56] & b[177])^(a[55] & b[178])^(a[54] & b[179])^(a[53] & b[180])^(a[52] & b[181])^(a[51] & b[182])^(a[50] & b[183])^(a[49] & b[184])^(a[48] & b[185])^(a[47] & b[186])^(a[46] & b[187])^(a[45] & b[188])^(a[44] & b[189])^(a[43] & b[190])^(a[42] & b[191])^(a[41] & b[192])^(a[40] & b[193])^(a[39] & b[194])^(a[38] & b[195])^(a[37] & b[196])^(a[36] & b[197])^(a[35] & b[198])^(a[34] & b[199])^(a[33] & b[200])^(a[32] & b[201])^(a[31] & b[202])^(a[30] & b[203])^(a[29] & b[204])^(a[28] & b[205])^(a[27] & b[206])^(a[26] & b[207])^(a[25] & b[208])^(a[24] & b[209])^(a[23] & b[210])^(a[22] & b[211])^(a[21] & b[212])^(a[20] & b[213])^(a[19] & b[214])^(a[18] & b[215])^(a[17] & b[216])^(a[16] & b[217])^(a[15] & b[218])^(a[14] & b[219])^(a[13] & b[220])^(a[12] & b[221])^(a[11] & b[222])^(a[10] & b[223])^(a[9] & b[224])^(a[8] & b[225])^(a[7] & b[226])^(a[6] & b[227])^(a[5] & b[228])^(a[4] & b[229])^(a[3] & b[230])^(a[2] & b[231])^(a[1] & b[232]);
assign y[234] = (a[232] & b[2])^(a[231] & b[3])^(a[230] & b[4])^(a[229] & b[5])^(a[228] & b[6])^(a[227] & b[7])^(a[226] & b[8])^(a[225] & b[9])^(a[224] & b[10])^(a[223] & b[11])^(a[222] & b[12])^(a[221] & b[13])^(a[220] & b[14])^(a[219] & b[15])^(a[218] & b[16])^(a[217] & b[17])^(a[216] & b[18])^(a[215] & b[19])^(a[214] & b[20])^(a[213] & b[21])^(a[212] & b[22])^(a[211] & b[23])^(a[210] & b[24])^(a[209] & b[25])^(a[208] & b[26])^(a[207] & b[27])^(a[206] & b[28])^(a[205] & b[29])^(a[204] & b[30])^(a[203] & b[31])^(a[202] & b[32])^(a[201] & b[33])^(a[200] & b[34])^(a[199] & b[35])^(a[198] & b[36])^(a[197] & b[37])^(a[196] & b[38])^(a[195] & b[39])^(a[194] & b[40])^(a[193] & b[41])^(a[192] & b[42])^(a[191] & b[43])^(a[190] & b[44])^(a[189] & b[45])^(a[188] & b[46])^(a[187] & b[47])^(a[186] & b[48])^(a[185] & b[49])^(a[184] & b[50])^(a[183] & b[51])^(a[182] & b[52])^(a[181] & b[53])^(a[180] & b[54])^(a[179] & b[55])^(a[178] & b[56])^(a[177] & b[57])^(a[176] & b[58])^(a[175] & b[59])^(a[174] & b[60])^(a[173] & b[61])^(a[172] & b[62])^(a[171] & b[63])^(a[170] & b[64])^(a[169] & b[65])^(a[168] & b[66])^(a[167] & b[67])^(a[166] & b[68])^(a[165] & b[69])^(a[164] & b[70])^(a[163] & b[71])^(a[162] & b[72])^(a[161] & b[73])^(a[160] & b[74])^(a[159] & b[75])^(a[158] & b[76])^(a[157] & b[77])^(a[156] & b[78])^(a[155] & b[79])^(a[154] & b[80])^(a[153] & b[81])^(a[152] & b[82])^(a[151] & b[83])^(a[150] & b[84])^(a[149] & b[85])^(a[148] & b[86])^(a[147] & b[87])^(a[146] & b[88])^(a[145] & b[89])^(a[144] & b[90])^(a[143] & b[91])^(a[142] & b[92])^(a[141] & b[93])^(a[140] & b[94])^(a[139] & b[95])^(a[138] & b[96])^(a[137] & b[97])^(a[136] & b[98])^(a[135] & b[99])^(a[134] & b[100])^(a[133] & b[101])^(a[132] & b[102])^(a[131] & b[103])^(a[130] & b[104])^(a[129] & b[105])^(a[128] & b[106])^(a[127] & b[107])^(a[126] & b[108])^(a[125] & b[109])^(a[124] & b[110])^(a[123] & b[111])^(a[122] & b[112])^(a[121] & b[113])^(a[120] & b[114])^(a[119] & b[115])^(a[118] & b[116])^(a[117] & b[117])^(a[116] & b[118])^(a[115] & b[119])^(a[114] & b[120])^(a[113] & b[121])^(a[112] & b[122])^(a[111] & b[123])^(a[110] & b[124])^(a[109] & b[125])^(a[108] & b[126])^(a[107] & b[127])^(a[106] & b[128])^(a[105] & b[129])^(a[104] & b[130])^(a[103] & b[131])^(a[102] & b[132])^(a[101] & b[133])^(a[100] & b[134])^(a[99] & b[135])^(a[98] & b[136])^(a[97] & b[137])^(a[96] & b[138])^(a[95] & b[139])^(a[94] & b[140])^(a[93] & b[141])^(a[92] & b[142])^(a[91] & b[143])^(a[90] & b[144])^(a[89] & b[145])^(a[88] & b[146])^(a[87] & b[147])^(a[86] & b[148])^(a[85] & b[149])^(a[84] & b[150])^(a[83] & b[151])^(a[82] & b[152])^(a[81] & b[153])^(a[80] & b[154])^(a[79] & b[155])^(a[78] & b[156])^(a[77] & b[157])^(a[76] & b[158])^(a[75] & b[159])^(a[74] & b[160])^(a[73] & b[161])^(a[72] & b[162])^(a[71] & b[163])^(a[70] & b[164])^(a[69] & b[165])^(a[68] & b[166])^(a[67] & b[167])^(a[66] & b[168])^(a[65] & b[169])^(a[64] & b[170])^(a[63] & b[171])^(a[62] & b[172])^(a[61] & b[173])^(a[60] & b[174])^(a[59] & b[175])^(a[58] & b[176])^(a[57] & b[177])^(a[56] & b[178])^(a[55] & b[179])^(a[54] & b[180])^(a[53] & b[181])^(a[52] & b[182])^(a[51] & b[183])^(a[50] & b[184])^(a[49] & b[185])^(a[48] & b[186])^(a[47] & b[187])^(a[46] & b[188])^(a[45] & b[189])^(a[44] & b[190])^(a[43] & b[191])^(a[42] & b[192])^(a[41] & b[193])^(a[40] & b[194])^(a[39] & b[195])^(a[38] & b[196])^(a[37] & b[197])^(a[36] & b[198])^(a[35] & b[199])^(a[34] & b[200])^(a[33] & b[201])^(a[32] & b[202])^(a[31] & b[203])^(a[30] & b[204])^(a[29] & b[205])^(a[28] & b[206])^(a[27] & b[207])^(a[26] & b[208])^(a[25] & b[209])^(a[24] & b[210])^(a[23] & b[211])^(a[22] & b[212])^(a[21] & b[213])^(a[20] & b[214])^(a[19] & b[215])^(a[18] & b[216])^(a[17] & b[217])^(a[16] & b[218])^(a[15] & b[219])^(a[14] & b[220])^(a[13] & b[221])^(a[12] & b[222])^(a[11] & b[223])^(a[10] & b[224])^(a[9] & b[225])^(a[8] & b[226])^(a[7] & b[227])^(a[6] & b[228])^(a[5] & b[229])^(a[4] & b[230])^(a[3] & b[231])^(a[2] & b[232]);
assign y[235] = (a[232] & b[3])^(a[231] & b[4])^(a[230] & b[5])^(a[229] & b[6])^(a[228] & b[7])^(a[227] & b[8])^(a[226] & b[9])^(a[225] & b[10])^(a[224] & b[11])^(a[223] & b[12])^(a[222] & b[13])^(a[221] & b[14])^(a[220] & b[15])^(a[219] & b[16])^(a[218] & b[17])^(a[217] & b[18])^(a[216] & b[19])^(a[215] & b[20])^(a[214] & b[21])^(a[213] & b[22])^(a[212] & b[23])^(a[211] & b[24])^(a[210] & b[25])^(a[209] & b[26])^(a[208] & b[27])^(a[207] & b[28])^(a[206] & b[29])^(a[205] & b[30])^(a[204] & b[31])^(a[203] & b[32])^(a[202] & b[33])^(a[201] & b[34])^(a[200] & b[35])^(a[199] & b[36])^(a[198] & b[37])^(a[197] & b[38])^(a[196] & b[39])^(a[195] & b[40])^(a[194] & b[41])^(a[193] & b[42])^(a[192] & b[43])^(a[191] & b[44])^(a[190] & b[45])^(a[189] & b[46])^(a[188] & b[47])^(a[187] & b[48])^(a[186] & b[49])^(a[185] & b[50])^(a[184] & b[51])^(a[183] & b[52])^(a[182] & b[53])^(a[181] & b[54])^(a[180] & b[55])^(a[179] & b[56])^(a[178] & b[57])^(a[177] & b[58])^(a[176] & b[59])^(a[175] & b[60])^(a[174] & b[61])^(a[173] & b[62])^(a[172] & b[63])^(a[171] & b[64])^(a[170] & b[65])^(a[169] & b[66])^(a[168] & b[67])^(a[167] & b[68])^(a[166] & b[69])^(a[165] & b[70])^(a[164] & b[71])^(a[163] & b[72])^(a[162] & b[73])^(a[161] & b[74])^(a[160] & b[75])^(a[159] & b[76])^(a[158] & b[77])^(a[157] & b[78])^(a[156] & b[79])^(a[155] & b[80])^(a[154] & b[81])^(a[153] & b[82])^(a[152] & b[83])^(a[151] & b[84])^(a[150] & b[85])^(a[149] & b[86])^(a[148] & b[87])^(a[147] & b[88])^(a[146] & b[89])^(a[145] & b[90])^(a[144] & b[91])^(a[143] & b[92])^(a[142] & b[93])^(a[141] & b[94])^(a[140] & b[95])^(a[139] & b[96])^(a[138] & b[97])^(a[137] & b[98])^(a[136] & b[99])^(a[135] & b[100])^(a[134] & b[101])^(a[133] & b[102])^(a[132] & b[103])^(a[131] & b[104])^(a[130] & b[105])^(a[129] & b[106])^(a[128] & b[107])^(a[127] & b[108])^(a[126] & b[109])^(a[125] & b[110])^(a[124] & b[111])^(a[123] & b[112])^(a[122] & b[113])^(a[121] & b[114])^(a[120] & b[115])^(a[119] & b[116])^(a[118] & b[117])^(a[117] & b[118])^(a[116] & b[119])^(a[115] & b[120])^(a[114] & b[121])^(a[113] & b[122])^(a[112] & b[123])^(a[111] & b[124])^(a[110] & b[125])^(a[109] & b[126])^(a[108] & b[127])^(a[107] & b[128])^(a[106] & b[129])^(a[105] & b[130])^(a[104] & b[131])^(a[103] & b[132])^(a[102] & b[133])^(a[101] & b[134])^(a[100] & b[135])^(a[99] & b[136])^(a[98] & b[137])^(a[97] & b[138])^(a[96] & b[139])^(a[95] & b[140])^(a[94] & b[141])^(a[93] & b[142])^(a[92] & b[143])^(a[91] & b[144])^(a[90] & b[145])^(a[89] & b[146])^(a[88] & b[147])^(a[87] & b[148])^(a[86] & b[149])^(a[85] & b[150])^(a[84] & b[151])^(a[83] & b[152])^(a[82] & b[153])^(a[81] & b[154])^(a[80] & b[155])^(a[79] & b[156])^(a[78] & b[157])^(a[77] & b[158])^(a[76] & b[159])^(a[75] & b[160])^(a[74] & b[161])^(a[73] & b[162])^(a[72] & b[163])^(a[71] & b[164])^(a[70] & b[165])^(a[69] & b[166])^(a[68] & b[167])^(a[67] & b[168])^(a[66] & b[169])^(a[65] & b[170])^(a[64] & b[171])^(a[63] & b[172])^(a[62] & b[173])^(a[61] & b[174])^(a[60] & b[175])^(a[59] & b[176])^(a[58] & b[177])^(a[57] & b[178])^(a[56] & b[179])^(a[55] & b[180])^(a[54] & b[181])^(a[53] & b[182])^(a[52] & b[183])^(a[51] & b[184])^(a[50] & b[185])^(a[49] & b[186])^(a[48] & b[187])^(a[47] & b[188])^(a[46] & b[189])^(a[45] & b[190])^(a[44] & b[191])^(a[43] & b[192])^(a[42] & b[193])^(a[41] & b[194])^(a[40] & b[195])^(a[39] & b[196])^(a[38] & b[197])^(a[37] & b[198])^(a[36] & b[199])^(a[35] & b[200])^(a[34] & b[201])^(a[33] & b[202])^(a[32] & b[203])^(a[31] & b[204])^(a[30] & b[205])^(a[29] & b[206])^(a[28] & b[207])^(a[27] & b[208])^(a[26] & b[209])^(a[25] & b[210])^(a[24] & b[211])^(a[23] & b[212])^(a[22] & b[213])^(a[21] & b[214])^(a[20] & b[215])^(a[19] & b[216])^(a[18] & b[217])^(a[17] & b[218])^(a[16] & b[219])^(a[15] & b[220])^(a[14] & b[221])^(a[13] & b[222])^(a[12] & b[223])^(a[11] & b[224])^(a[10] & b[225])^(a[9] & b[226])^(a[8] & b[227])^(a[7] & b[228])^(a[6] & b[229])^(a[5] & b[230])^(a[4] & b[231])^(a[3] & b[232]);
assign y[236] = (a[232] & b[4])^(a[231] & b[5])^(a[230] & b[6])^(a[229] & b[7])^(a[228] & b[8])^(a[227] & b[9])^(a[226] & b[10])^(a[225] & b[11])^(a[224] & b[12])^(a[223] & b[13])^(a[222] & b[14])^(a[221] & b[15])^(a[220] & b[16])^(a[219] & b[17])^(a[218] & b[18])^(a[217] & b[19])^(a[216] & b[20])^(a[215] & b[21])^(a[214] & b[22])^(a[213] & b[23])^(a[212] & b[24])^(a[211] & b[25])^(a[210] & b[26])^(a[209] & b[27])^(a[208] & b[28])^(a[207] & b[29])^(a[206] & b[30])^(a[205] & b[31])^(a[204] & b[32])^(a[203] & b[33])^(a[202] & b[34])^(a[201] & b[35])^(a[200] & b[36])^(a[199] & b[37])^(a[198] & b[38])^(a[197] & b[39])^(a[196] & b[40])^(a[195] & b[41])^(a[194] & b[42])^(a[193] & b[43])^(a[192] & b[44])^(a[191] & b[45])^(a[190] & b[46])^(a[189] & b[47])^(a[188] & b[48])^(a[187] & b[49])^(a[186] & b[50])^(a[185] & b[51])^(a[184] & b[52])^(a[183] & b[53])^(a[182] & b[54])^(a[181] & b[55])^(a[180] & b[56])^(a[179] & b[57])^(a[178] & b[58])^(a[177] & b[59])^(a[176] & b[60])^(a[175] & b[61])^(a[174] & b[62])^(a[173] & b[63])^(a[172] & b[64])^(a[171] & b[65])^(a[170] & b[66])^(a[169] & b[67])^(a[168] & b[68])^(a[167] & b[69])^(a[166] & b[70])^(a[165] & b[71])^(a[164] & b[72])^(a[163] & b[73])^(a[162] & b[74])^(a[161] & b[75])^(a[160] & b[76])^(a[159] & b[77])^(a[158] & b[78])^(a[157] & b[79])^(a[156] & b[80])^(a[155] & b[81])^(a[154] & b[82])^(a[153] & b[83])^(a[152] & b[84])^(a[151] & b[85])^(a[150] & b[86])^(a[149] & b[87])^(a[148] & b[88])^(a[147] & b[89])^(a[146] & b[90])^(a[145] & b[91])^(a[144] & b[92])^(a[143] & b[93])^(a[142] & b[94])^(a[141] & b[95])^(a[140] & b[96])^(a[139] & b[97])^(a[138] & b[98])^(a[137] & b[99])^(a[136] & b[100])^(a[135] & b[101])^(a[134] & b[102])^(a[133] & b[103])^(a[132] & b[104])^(a[131] & b[105])^(a[130] & b[106])^(a[129] & b[107])^(a[128] & b[108])^(a[127] & b[109])^(a[126] & b[110])^(a[125] & b[111])^(a[124] & b[112])^(a[123] & b[113])^(a[122] & b[114])^(a[121] & b[115])^(a[120] & b[116])^(a[119] & b[117])^(a[118] & b[118])^(a[117] & b[119])^(a[116] & b[120])^(a[115] & b[121])^(a[114] & b[122])^(a[113] & b[123])^(a[112] & b[124])^(a[111] & b[125])^(a[110] & b[126])^(a[109] & b[127])^(a[108] & b[128])^(a[107] & b[129])^(a[106] & b[130])^(a[105] & b[131])^(a[104] & b[132])^(a[103] & b[133])^(a[102] & b[134])^(a[101] & b[135])^(a[100] & b[136])^(a[99] & b[137])^(a[98] & b[138])^(a[97] & b[139])^(a[96] & b[140])^(a[95] & b[141])^(a[94] & b[142])^(a[93] & b[143])^(a[92] & b[144])^(a[91] & b[145])^(a[90] & b[146])^(a[89] & b[147])^(a[88] & b[148])^(a[87] & b[149])^(a[86] & b[150])^(a[85] & b[151])^(a[84] & b[152])^(a[83] & b[153])^(a[82] & b[154])^(a[81] & b[155])^(a[80] & b[156])^(a[79] & b[157])^(a[78] & b[158])^(a[77] & b[159])^(a[76] & b[160])^(a[75] & b[161])^(a[74] & b[162])^(a[73] & b[163])^(a[72] & b[164])^(a[71] & b[165])^(a[70] & b[166])^(a[69] & b[167])^(a[68] & b[168])^(a[67] & b[169])^(a[66] & b[170])^(a[65] & b[171])^(a[64] & b[172])^(a[63] & b[173])^(a[62] & b[174])^(a[61] & b[175])^(a[60] & b[176])^(a[59] & b[177])^(a[58] & b[178])^(a[57] & b[179])^(a[56] & b[180])^(a[55] & b[181])^(a[54] & b[182])^(a[53] & b[183])^(a[52] & b[184])^(a[51] & b[185])^(a[50] & b[186])^(a[49] & b[187])^(a[48] & b[188])^(a[47] & b[189])^(a[46] & b[190])^(a[45] & b[191])^(a[44] & b[192])^(a[43] & b[193])^(a[42] & b[194])^(a[41] & b[195])^(a[40] & b[196])^(a[39] & b[197])^(a[38] & b[198])^(a[37] & b[199])^(a[36] & b[200])^(a[35] & b[201])^(a[34] & b[202])^(a[33] & b[203])^(a[32] & b[204])^(a[31] & b[205])^(a[30] & b[206])^(a[29] & b[207])^(a[28] & b[208])^(a[27] & b[209])^(a[26] & b[210])^(a[25] & b[211])^(a[24] & b[212])^(a[23] & b[213])^(a[22] & b[214])^(a[21] & b[215])^(a[20] & b[216])^(a[19] & b[217])^(a[18] & b[218])^(a[17] & b[219])^(a[16] & b[220])^(a[15] & b[221])^(a[14] & b[222])^(a[13] & b[223])^(a[12] & b[224])^(a[11] & b[225])^(a[10] & b[226])^(a[9] & b[227])^(a[8] & b[228])^(a[7] & b[229])^(a[6] & b[230])^(a[5] & b[231])^(a[4] & b[232]);
assign y[237] = (a[232] & b[5])^(a[231] & b[6])^(a[230] & b[7])^(a[229] & b[8])^(a[228] & b[9])^(a[227] & b[10])^(a[226] & b[11])^(a[225] & b[12])^(a[224] & b[13])^(a[223] & b[14])^(a[222] & b[15])^(a[221] & b[16])^(a[220] & b[17])^(a[219] & b[18])^(a[218] & b[19])^(a[217] & b[20])^(a[216] & b[21])^(a[215] & b[22])^(a[214] & b[23])^(a[213] & b[24])^(a[212] & b[25])^(a[211] & b[26])^(a[210] & b[27])^(a[209] & b[28])^(a[208] & b[29])^(a[207] & b[30])^(a[206] & b[31])^(a[205] & b[32])^(a[204] & b[33])^(a[203] & b[34])^(a[202] & b[35])^(a[201] & b[36])^(a[200] & b[37])^(a[199] & b[38])^(a[198] & b[39])^(a[197] & b[40])^(a[196] & b[41])^(a[195] & b[42])^(a[194] & b[43])^(a[193] & b[44])^(a[192] & b[45])^(a[191] & b[46])^(a[190] & b[47])^(a[189] & b[48])^(a[188] & b[49])^(a[187] & b[50])^(a[186] & b[51])^(a[185] & b[52])^(a[184] & b[53])^(a[183] & b[54])^(a[182] & b[55])^(a[181] & b[56])^(a[180] & b[57])^(a[179] & b[58])^(a[178] & b[59])^(a[177] & b[60])^(a[176] & b[61])^(a[175] & b[62])^(a[174] & b[63])^(a[173] & b[64])^(a[172] & b[65])^(a[171] & b[66])^(a[170] & b[67])^(a[169] & b[68])^(a[168] & b[69])^(a[167] & b[70])^(a[166] & b[71])^(a[165] & b[72])^(a[164] & b[73])^(a[163] & b[74])^(a[162] & b[75])^(a[161] & b[76])^(a[160] & b[77])^(a[159] & b[78])^(a[158] & b[79])^(a[157] & b[80])^(a[156] & b[81])^(a[155] & b[82])^(a[154] & b[83])^(a[153] & b[84])^(a[152] & b[85])^(a[151] & b[86])^(a[150] & b[87])^(a[149] & b[88])^(a[148] & b[89])^(a[147] & b[90])^(a[146] & b[91])^(a[145] & b[92])^(a[144] & b[93])^(a[143] & b[94])^(a[142] & b[95])^(a[141] & b[96])^(a[140] & b[97])^(a[139] & b[98])^(a[138] & b[99])^(a[137] & b[100])^(a[136] & b[101])^(a[135] & b[102])^(a[134] & b[103])^(a[133] & b[104])^(a[132] & b[105])^(a[131] & b[106])^(a[130] & b[107])^(a[129] & b[108])^(a[128] & b[109])^(a[127] & b[110])^(a[126] & b[111])^(a[125] & b[112])^(a[124] & b[113])^(a[123] & b[114])^(a[122] & b[115])^(a[121] & b[116])^(a[120] & b[117])^(a[119] & b[118])^(a[118] & b[119])^(a[117] & b[120])^(a[116] & b[121])^(a[115] & b[122])^(a[114] & b[123])^(a[113] & b[124])^(a[112] & b[125])^(a[111] & b[126])^(a[110] & b[127])^(a[109] & b[128])^(a[108] & b[129])^(a[107] & b[130])^(a[106] & b[131])^(a[105] & b[132])^(a[104] & b[133])^(a[103] & b[134])^(a[102] & b[135])^(a[101] & b[136])^(a[100] & b[137])^(a[99] & b[138])^(a[98] & b[139])^(a[97] & b[140])^(a[96] & b[141])^(a[95] & b[142])^(a[94] & b[143])^(a[93] & b[144])^(a[92] & b[145])^(a[91] & b[146])^(a[90] & b[147])^(a[89] & b[148])^(a[88] & b[149])^(a[87] & b[150])^(a[86] & b[151])^(a[85] & b[152])^(a[84] & b[153])^(a[83] & b[154])^(a[82] & b[155])^(a[81] & b[156])^(a[80] & b[157])^(a[79] & b[158])^(a[78] & b[159])^(a[77] & b[160])^(a[76] & b[161])^(a[75] & b[162])^(a[74] & b[163])^(a[73] & b[164])^(a[72] & b[165])^(a[71] & b[166])^(a[70] & b[167])^(a[69] & b[168])^(a[68] & b[169])^(a[67] & b[170])^(a[66] & b[171])^(a[65] & b[172])^(a[64] & b[173])^(a[63] & b[174])^(a[62] & b[175])^(a[61] & b[176])^(a[60] & b[177])^(a[59] & b[178])^(a[58] & b[179])^(a[57] & b[180])^(a[56] & b[181])^(a[55] & b[182])^(a[54] & b[183])^(a[53] & b[184])^(a[52] & b[185])^(a[51] & b[186])^(a[50] & b[187])^(a[49] & b[188])^(a[48] & b[189])^(a[47] & b[190])^(a[46] & b[191])^(a[45] & b[192])^(a[44] & b[193])^(a[43] & b[194])^(a[42] & b[195])^(a[41] & b[196])^(a[40] & b[197])^(a[39] & b[198])^(a[38] & b[199])^(a[37] & b[200])^(a[36] & b[201])^(a[35] & b[202])^(a[34] & b[203])^(a[33] & b[204])^(a[32] & b[205])^(a[31] & b[206])^(a[30] & b[207])^(a[29] & b[208])^(a[28] & b[209])^(a[27] & b[210])^(a[26] & b[211])^(a[25] & b[212])^(a[24] & b[213])^(a[23] & b[214])^(a[22] & b[215])^(a[21] & b[216])^(a[20] & b[217])^(a[19] & b[218])^(a[18] & b[219])^(a[17] & b[220])^(a[16] & b[221])^(a[15] & b[222])^(a[14] & b[223])^(a[13] & b[224])^(a[12] & b[225])^(a[11] & b[226])^(a[10] & b[227])^(a[9] & b[228])^(a[8] & b[229])^(a[7] & b[230])^(a[6] & b[231])^(a[5] & b[232]);
assign y[238] = (a[232] & b[6])^(a[231] & b[7])^(a[230] & b[8])^(a[229] & b[9])^(a[228] & b[10])^(a[227] & b[11])^(a[226] & b[12])^(a[225] & b[13])^(a[224] & b[14])^(a[223] & b[15])^(a[222] & b[16])^(a[221] & b[17])^(a[220] & b[18])^(a[219] & b[19])^(a[218] & b[20])^(a[217] & b[21])^(a[216] & b[22])^(a[215] & b[23])^(a[214] & b[24])^(a[213] & b[25])^(a[212] & b[26])^(a[211] & b[27])^(a[210] & b[28])^(a[209] & b[29])^(a[208] & b[30])^(a[207] & b[31])^(a[206] & b[32])^(a[205] & b[33])^(a[204] & b[34])^(a[203] & b[35])^(a[202] & b[36])^(a[201] & b[37])^(a[200] & b[38])^(a[199] & b[39])^(a[198] & b[40])^(a[197] & b[41])^(a[196] & b[42])^(a[195] & b[43])^(a[194] & b[44])^(a[193] & b[45])^(a[192] & b[46])^(a[191] & b[47])^(a[190] & b[48])^(a[189] & b[49])^(a[188] & b[50])^(a[187] & b[51])^(a[186] & b[52])^(a[185] & b[53])^(a[184] & b[54])^(a[183] & b[55])^(a[182] & b[56])^(a[181] & b[57])^(a[180] & b[58])^(a[179] & b[59])^(a[178] & b[60])^(a[177] & b[61])^(a[176] & b[62])^(a[175] & b[63])^(a[174] & b[64])^(a[173] & b[65])^(a[172] & b[66])^(a[171] & b[67])^(a[170] & b[68])^(a[169] & b[69])^(a[168] & b[70])^(a[167] & b[71])^(a[166] & b[72])^(a[165] & b[73])^(a[164] & b[74])^(a[163] & b[75])^(a[162] & b[76])^(a[161] & b[77])^(a[160] & b[78])^(a[159] & b[79])^(a[158] & b[80])^(a[157] & b[81])^(a[156] & b[82])^(a[155] & b[83])^(a[154] & b[84])^(a[153] & b[85])^(a[152] & b[86])^(a[151] & b[87])^(a[150] & b[88])^(a[149] & b[89])^(a[148] & b[90])^(a[147] & b[91])^(a[146] & b[92])^(a[145] & b[93])^(a[144] & b[94])^(a[143] & b[95])^(a[142] & b[96])^(a[141] & b[97])^(a[140] & b[98])^(a[139] & b[99])^(a[138] & b[100])^(a[137] & b[101])^(a[136] & b[102])^(a[135] & b[103])^(a[134] & b[104])^(a[133] & b[105])^(a[132] & b[106])^(a[131] & b[107])^(a[130] & b[108])^(a[129] & b[109])^(a[128] & b[110])^(a[127] & b[111])^(a[126] & b[112])^(a[125] & b[113])^(a[124] & b[114])^(a[123] & b[115])^(a[122] & b[116])^(a[121] & b[117])^(a[120] & b[118])^(a[119] & b[119])^(a[118] & b[120])^(a[117] & b[121])^(a[116] & b[122])^(a[115] & b[123])^(a[114] & b[124])^(a[113] & b[125])^(a[112] & b[126])^(a[111] & b[127])^(a[110] & b[128])^(a[109] & b[129])^(a[108] & b[130])^(a[107] & b[131])^(a[106] & b[132])^(a[105] & b[133])^(a[104] & b[134])^(a[103] & b[135])^(a[102] & b[136])^(a[101] & b[137])^(a[100] & b[138])^(a[99] & b[139])^(a[98] & b[140])^(a[97] & b[141])^(a[96] & b[142])^(a[95] & b[143])^(a[94] & b[144])^(a[93] & b[145])^(a[92] & b[146])^(a[91] & b[147])^(a[90] & b[148])^(a[89] & b[149])^(a[88] & b[150])^(a[87] & b[151])^(a[86] & b[152])^(a[85] & b[153])^(a[84] & b[154])^(a[83] & b[155])^(a[82] & b[156])^(a[81] & b[157])^(a[80] & b[158])^(a[79] & b[159])^(a[78] & b[160])^(a[77] & b[161])^(a[76] & b[162])^(a[75] & b[163])^(a[74] & b[164])^(a[73] & b[165])^(a[72] & b[166])^(a[71] & b[167])^(a[70] & b[168])^(a[69] & b[169])^(a[68] & b[170])^(a[67] & b[171])^(a[66] & b[172])^(a[65] & b[173])^(a[64] & b[174])^(a[63] & b[175])^(a[62] & b[176])^(a[61] & b[177])^(a[60] & b[178])^(a[59] & b[179])^(a[58] & b[180])^(a[57] & b[181])^(a[56] & b[182])^(a[55] & b[183])^(a[54] & b[184])^(a[53] & b[185])^(a[52] & b[186])^(a[51] & b[187])^(a[50] & b[188])^(a[49] & b[189])^(a[48] & b[190])^(a[47] & b[191])^(a[46] & b[192])^(a[45] & b[193])^(a[44] & b[194])^(a[43] & b[195])^(a[42] & b[196])^(a[41] & b[197])^(a[40] & b[198])^(a[39] & b[199])^(a[38] & b[200])^(a[37] & b[201])^(a[36] & b[202])^(a[35] & b[203])^(a[34] & b[204])^(a[33] & b[205])^(a[32] & b[206])^(a[31] & b[207])^(a[30] & b[208])^(a[29] & b[209])^(a[28] & b[210])^(a[27] & b[211])^(a[26] & b[212])^(a[25] & b[213])^(a[24] & b[214])^(a[23] & b[215])^(a[22] & b[216])^(a[21] & b[217])^(a[20] & b[218])^(a[19] & b[219])^(a[18] & b[220])^(a[17] & b[221])^(a[16] & b[222])^(a[15] & b[223])^(a[14] & b[224])^(a[13] & b[225])^(a[12] & b[226])^(a[11] & b[227])^(a[10] & b[228])^(a[9] & b[229])^(a[8] & b[230])^(a[7] & b[231])^(a[6] & b[232]);
assign y[239] = (a[232] & b[7])^(a[231] & b[8])^(a[230] & b[9])^(a[229] & b[10])^(a[228] & b[11])^(a[227] & b[12])^(a[226] & b[13])^(a[225] & b[14])^(a[224] & b[15])^(a[223] & b[16])^(a[222] & b[17])^(a[221] & b[18])^(a[220] & b[19])^(a[219] & b[20])^(a[218] & b[21])^(a[217] & b[22])^(a[216] & b[23])^(a[215] & b[24])^(a[214] & b[25])^(a[213] & b[26])^(a[212] & b[27])^(a[211] & b[28])^(a[210] & b[29])^(a[209] & b[30])^(a[208] & b[31])^(a[207] & b[32])^(a[206] & b[33])^(a[205] & b[34])^(a[204] & b[35])^(a[203] & b[36])^(a[202] & b[37])^(a[201] & b[38])^(a[200] & b[39])^(a[199] & b[40])^(a[198] & b[41])^(a[197] & b[42])^(a[196] & b[43])^(a[195] & b[44])^(a[194] & b[45])^(a[193] & b[46])^(a[192] & b[47])^(a[191] & b[48])^(a[190] & b[49])^(a[189] & b[50])^(a[188] & b[51])^(a[187] & b[52])^(a[186] & b[53])^(a[185] & b[54])^(a[184] & b[55])^(a[183] & b[56])^(a[182] & b[57])^(a[181] & b[58])^(a[180] & b[59])^(a[179] & b[60])^(a[178] & b[61])^(a[177] & b[62])^(a[176] & b[63])^(a[175] & b[64])^(a[174] & b[65])^(a[173] & b[66])^(a[172] & b[67])^(a[171] & b[68])^(a[170] & b[69])^(a[169] & b[70])^(a[168] & b[71])^(a[167] & b[72])^(a[166] & b[73])^(a[165] & b[74])^(a[164] & b[75])^(a[163] & b[76])^(a[162] & b[77])^(a[161] & b[78])^(a[160] & b[79])^(a[159] & b[80])^(a[158] & b[81])^(a[157] & b[82])^(a[156] & b[83])^(a[155] & b[84])^(a[154] & b[85])^(a[153] & b[86])^(a[152] & b[87])^(a[151] & b[88])^(a[150] & b[89])^(a[149] & b[90])^(a[148] & b[91])^(a[147] & b[92])^(a[146] & b[93])^(a[145] & b[94])^(a[144] & b[95])^(a[143] & b[96])^(a[142] & b[97])^(a[141] & b[98])^(a[140] & b[99])^(a[139] & b[100])^(a[138] & b[101])^(a[137] & b[102])^(a[136] & b[103])^(a[135] & b[104])^(a[134] & b[105])^(a[133] & b[106])^(a[132] & b[107])^(a[131] & b[108])^(a[130] & b[109])^(a[129] & b[110])^(a[128] & b[111])^(a[127] & b[112])^(a[126] & b[113])^(a[125] & b[114])^(a[124] & b[115])^(a[123] & b[116])^(a[122] & b[117])^(a[121] & b[118])^(a[120] & b[119])^(a[119] & b[120])^(a[118] & b[121])^(a[117] & b[122])^(a[116] & b[123])^(a[115] & b[124])^(a[114] & b[125])^(a[113] & b[126])^(a[112] & b[127])^(a[111] & b[128])^(a[110] & b[129])^(a[109] & b[130])^(a[108] & b[131])^(a[107] & b[132])^(a[106] & b[133])^(a[105] & b[134])^(a[104] & b[135])^(a[103] & b[136])^(a[102] & b[137])^(a[101] & b[138])^(a[100] & b[139])^(a[99] & b[140])^(a[98] & b[141])^(a[97] & b[142])^(a[96] & b[143])^(a[95] & b[144])^(a[94] & b[145])^(a[93] & b[146])^(a[92] & b[147])^(a[91] & b[148])^(a[90] & b[149])^(a[89] & b[150])^(a[88] & b[151])^(a[87] & b[152])^(a[86] & b[153])^(a[85] & b[154])^(a[84] & b[155])^(a[83] & b[156])^(a[82] & b[157])^(a[81] & b[158])^(a[80] & b[159])^(a[79] & b[160])^(a[78] & b[161])^(a[77] & b[162])^(a[76] & b[163])^(a[75] & b[164])^(a[74] & b[165])^(a[73] & b[166])^(a[72] & b[167])^(a[71] & b[168])^(a[70] & b[169])^(a[69] & b[170])^(a[68] & b[171])^(a[67] & b[172])^(a[66] & b[173])^(a[65] & b[174])^(a[64] & b[175])^(a[63] & b[176])^(a[62] & b[177])^(a[61] & b[178])^(a[60] & b[179])^(a[59] & b[180])^(a[58] & b[181])^(a[57] & b[182])^(a[56] & b[183])^(a[55] & b[184])^(a[54] & b[185])^(a[53] & b[186])^(a[52] & b[187])^(a[51] & b[188])^(a[50] & b[189])^(a[49] & b[190])^(a[48] & b[191])^(a[47] & b[192])^(a[46] & b[193])^(a[45] & b[194])^(a[44] & b[195])^(a[43] & b[196])^(a[42] & b[197])^(a[41] & b[198])^(a[40] & b[199])^(a[39] & b[200])^(a[38] & b[201])^(a[37] & b[202])^(a[36] & b[203])^(a[35] & b[204])^(a[34] & b[205])^(a[33] & b[206])^(a[32] & b[207])^(a[31] & b[208])^(a[30] & b[209])^(a[29] & b[210])^(a[28] & b[211])^(a[27] & b[212])^(a[26] & b[213])^(a[25] & b[214])^(a[24] & b[215])^(a[23] & b[216])^(a[22] & b[217])^(a[21] & b[218])^(a[20] & b[219])^(a[19] & b[220])^(a[18] & b[221])^(a[17] & b[222])^(a[16] & b[223])^(a[15] & b[224])^(a[14] & b[225])^(a[13] & b[226])^(a[12] & b[227])^(a[11] & b[228])^(a[10] & b[229])^(a[9] & b[230])^(a[8] & b[231])^(a[7] & b[232]);
assign y[240] = (a[232] & b[8])^(a[231] & b[9])^(a[230] & b[10])^(a[229] & b[11])^(a[228] & b[12])^(a[227] & b[13])^(a[226] & b[14])^(a[225] & b[15])^(a[224] & b[16])^(a[223] & b[17])^(a[222] & b[18])^(a[221] & b[19])^(a[220] & b[20])^(a[219] & b[21])^(a[218] & b[22])^(a[217] & b[23])^(a[216] & b[24])^(a[215] & b[25])^(a[214] & b[26])^(a[213] & b[27])^(a[212] & b[28])^(a[211] & b[29])^(a[210] & b[30])^(a[209] & b[31])^(a[208] & b[32])^(a[207] & b[33])^(a[206] & b[34])^(a[205] & b[35])^(a[204] & b[36])^(a[203] & b[37])^(a[202] & b[38])^(a[201] & b[39])^(a[200] & b[40])^(a[199] & b[41])^(a[198] & b[42])^(a[197] & b[43])^(a[196] & b[44])^(a[195] & b[45])^(a[194] & b[46])^(a[193] & b[47])^(a[192] & b[48])^(a[191] & b[49])^(a[190] & b[50])^(a[189] & b[51])^(a[188] & b[52])^(a[187] & b[53])^(a[186] & b[54])^(a[185] & b[55])^(a[184] & b[56])^(a[183] & b[57])^(a[182] & b[58])^(a[181] & b[59])^(a[180] & b[60])^(a[179] & b[61])^(a[178] & b[62])^(a[177] & b[63])^(a[176] & b[64])^(a[175] & b[65])^(a[174] & b[66])^(a[173] & b[67])^(a[172] & b[68])^(a[171] & b[69])^(a[170] & b[70])^(a[169] & b[71])^(a[168] & b[72])^(a[167] & b[73])^(a[166] & b[74])^(a[165] & b[75])^(a[164] & b[76])^(a[163] & b[77])^(a[162] & b[78])^(a[161] & b[79])^(a[160] & b[80])^(a[159] & b[81])^(a[158] & b[82])^(a[157] & b[83])^(a[156] & b[84])^(a[155] & b[85])^(a[154] & b[86])^(a[153] & b[87])^(a[152] & b[88])^(a[151] & b[89])^(a[150] & b[90])^(a[149] & b[91])^(a[148] & b[92])^(a[147] & b[93])^(a[146] & b[94])^(a[145] & b[95])^(a[144] & b[96])^(a[143] & b[97])^(a[142] & b[98])^(a[141] & b[99])^(a[140] & b[100])^(a[139] & b[101])^(a[138] & b[102])^(a[137] & b[103])^(a[136] & b[104])^(a[135] & b[105])^(a[134] & b[106])^(a[133] & b[107])^(a[132] & b[108])^(a[131] & b[109])^(a[130] & b[110])^(a[129] & b[111])^(a[128] & b[112])^(a[127] & b[113])^(a[126] & b[114])^(a[125] & b[115])^(a[124] & b[116])^(a[123] & b[117])^(a[122] & b[118])^(a[121] & b[119])^(a[120] & b[120])^(a[119] & b[121])^(a[118] & b[122])^(a[117] & b[123])^(a[116] & b[124])^(a[115] & b[125])^(a[114] & b[126])^(a[113] & b[127])^(a[112] & b[128])^(a[111] & b[129])^(a[110] & b[130])^(a[109] & b[131])^(a[108] & b[132])^(a[107] & b[133])^(a[106] & b[134])^(a[105] & b[135])^(a[104] & b[136])^(a[103] & b[137])^(a[102] & b[138])^(a[101] & b[139])^(a[100] & b[140])^(a[99] & b[141])^(a[98] & b[142])^(a[97] & b[143])^(a[96] & b[144])^(a[95] & b[145])^(a[94] & b[146])^(a[93] & b[147])^(a[92] & b[148])^(a[91] & b[149])^(a[90] & b[150])^(a[89] & b[151])^(a[88] & b[152])^(a[87] & b[153])^(a[86] & b[154])^(a[85] & b[155])^(a[84] & b[156])^(a[83] & b[157])^(a[82] & b[158])^(a[81] & b[159])^(a[80] & b[160])^(a[79] & b[161])^(a[78] & b[162])^(a[77] & b[163])^(a[76] & b[164])^(a[75] & b[165])^(a[74] & b[166])^(a[73] & b[167])^(a[72] & b[168])^(a[71] & b[169])^(a[70] & b[170])^(a[69] & b[171])^(a[68] & b[172])^(a[67] & b[173])^(a[66] & b[174])^(a[65] & b[175])^(a[64] & b[176])^(a[63] & b[177])^(a[62] & b[178])^(a[61] & b[179])^(a[60] & b[180])^(a[59] & b[181])^(a[58] & b[182])^(a[57] & b[183])^(a[56] & b[184])^(a[55] & b[185])^(a[54] & b[186])^(a[53] & b[187])^(a[52] & b[188])^(a[51] & b[189])^(a[50] & b[190])^(a[49] & b[191])^(a[48] & b[192])^(a[47] & b[193])^(a[46] & b[194])^(a[45] & b[195])^(a[44] & b[196])^(a[43] & b[197])^(a[42] & b[198])^(a[41] & b[199])^(a[40] & b[200])^(a[39] & b[201])^(a[38] & b[202])^(a[37] & b[203])^(a[36] & b[204])^(a[35] & b[205])^(a[34] & b[206])^(a[33] & b[207])^(a[32] & b[208])^(a[31] & b[209])^(a[30] & b[210])^(a[29] & b[211])^(a[28] & b[212])^(a[27] & b[213])^(a[26] & b[214])^(a[25] & b[215])^(a[24] & b[216])^(a[23] & b[217])^(a[22] & b[218])^(a[21] & b[219])^(a[20] & b[220])^(a[19] & b[221])^(a[18] & b[222])^(a[17] & b[223])^(a[16] & b[224])^(a[15] & b[225])^(a[14] & b[226])^(a[13] & b[227])^(a[12] & b[228])^(a[11] & b[229])^(a[10] & b[230])^(a[9] & b[231])^(a[8] & b[232]);
assign y[241] = (a[232] & b[9])^(a[231] & b[10])^(a[230] & b[11])^(a[229] & b[12])^(a[228] & b[13])^(a[227] & b[14])^(a[226] & b[15])^(a[225] & b[16])^(a[224] & b[17])^(a[223] & b[18])^(a[222] & b[19])^(a[221] & b[20])^(a[220] & b[21])^(a[219] & b[22])^(a[218] & b[23])^(a[217] & b[24])^(a[216] & b[25])^(a[215] & b[26])^(a[214] & b[27])^(a[213] & b[28])^(a[212] & b[29])^(a[211] & b[30])^(a[210] & b[31])^(a[209] & b[32])^(a[208] & b[33])^(a[207] & b[34])^(a[206] & b[35])^(a[205] & b[36])^(a[204] & b[37])^(a[203] & b[38])^(a[202] & b[39])^(a[201] & b[40])^(a[200] & b[41])^(a[199] & b[42])^(a[198] & b[43])^(a[197] & b[44])^(a[196] & b[45])^(a[195] & b[46])^(a[194] & b[47])^(a[193] & b[48])^(a[192] & b[49])^(a[191] & b[50])^(a[190] & b[51])^(a[189] & b[52])^(a[188] & b[53])^(a[187] & b[54])^(a[186] & b[55])^(a[185] & b[56])^(a[184] & b[57])^(a[183] & b[58])^(a[182] & b[59])^(a[181] & b[60])^(a[180] & b[61])^(a[179] & b[62])^(a[178] & b[63])^(a[177] & b[64])^(a[176] & b[65])^(a[175] & b[66])^(a[174] & b[67])^(a[173] & b[68])^(a[172] & b[69])^(a[171] & b[70])^(a[170] & b[71])^(a[169] & b[72])^(a[168] & b[73])^(a[167] & b[74])^(a[166] & b[75])^(a[165] & b[76])^(a[164] & b[77])^(a[163] & b[78])^(a[162] & b[79])^(a[161] & b[80])^(a[160] & b[81])^(a[159] & b[82])^(a[158] & b[83])^(a[157] & b[84])^(a[156] & b[85])^(a[155] & b[86])^(a[154] & b[87])^(a[153] & b[88])^(a[152] & b[89])^(a[151] & b[90])^(a[150] & b[91])^(a[149] & b[92])^(a[148] & b[93])^(a[147] & b[94])^(a[146] & b[95])^(a[145] & b[96])^(a[144] & b[97])^(a[143] & b[98])^(a[142] & b[99])^(a[141] & b[100])^(a[140] & b[101])^(a[139] & b[102])^(a[138] & b[103])^(a[137] & b[104])^(a[136] & b[105])^(a[135] & b[106])^(a[134] & b[107])^(a[133] & b[108])^(a[132] & b[109])^(a[131] & b[110])^(a[130] & b[111])^(a[129] & b[112])^(a[128] & b[113])^(a[127] & b[114])^(a[126] & b[115])^(a[125] & b[116])^(a[124] & b[117])^(a[123] & b[118])^(a[122] & b[119])^(a[121] & b[120])^(a[120] & b[121])^(a[119] & b[122])^(a[118] & b[123])^(a[117] & b[124])^(a[116] & b[125])^(a[115] & b[126])^(a[114] & b[127])^(a[113] & b[128])^(a[112] & b[129])^(a[111] & b[130])^(a[110] & b[131])^(a[109] & b[132])^(a[108] & b[133])^(a[107] & b[134])^(a[106] & b[135])^(a[105] & b[136])^(a[104] & b[137])^(a[103] & b[138])^(a[102] & b[139])^(a[101] & b[140])^(a[100] & b[141])^(a[99] & b[142])^(a[98] & b[143])^(a[97] & b[144])^(a[96] & b[145])^(a[95] & b[146])^(a[94] & b[147])^(a[93] & b[148])^(a[92] & b[149])^(a[91] & b[150])^(a[90] & b[151])^(a[89] & b[152])^(a[88] & b[153])^(a[87] & b[154])^(a[86] & b[155])^(a[85] & b[156])^(a[84] & b[157])^(a[83] & b[158])^(a[82] & b[159])^(a[81] & b[160])^(a[80] & b[161])^(a[79] & b[162])^(a[78] & b[163])^(a[77] & b[164])^(a[76] & b[165])^(a[75] & b[166])^(a[74] & b[167])^(a[73] & b[168])^(a[72] & b[169])^(a[71] & b[170])^(a[70] & b[171])^(a[69] & b[172])^(a[68] & b[173])^(a[67] & b[174])^(a[66] & b[175])^(a[65] & b[176])^(a[64] & b[177])^(a[63] & b[178])^(a[62] & b[179])^(a[61] & b[180])^(a[60] & b[181])^(a[59] & b[182])^(a[58] & b[183])^(a[57] & b[184])^(a[56] & b[185])^(a[55] & b[186])^(a[54] & b[187])^(a[53] & b[188])^(a[52] & b[189])^(a[51] & b[190])^(a[50] & b[191])^(a[49] & b[192])^(a[48] & b[193])^(a[47] & b[194])^(a[46] & b[195])^(a[45] & b[196])^(a[44] & b[197])^(a[43] & b[198])^(a[42] & b[199])^(a[41] & b[200])^(a[40] & b[201])^(a[39] & b[202])^(a[38] & b[203])^(a[37] & b[204])^(a[36] & b[205])^(a[35] & b[206])^(a[34] & b[207])^(a[33] & b[208])^(a[32] & b[209])^(a[31] & b[210])^(a[30] & b[211])^(a[29] & b[212])^(a[28] & b[213])^(a[27] & b[214])^(a[26] & b[215])^(a[25] & b[216])^(a[24] & b[217])^(a[23] & b[218])^(a[22] & b[219])^(a[21] & b[220])^(a[20] & b[221])^(a[19] & b[222])^(a[18] & b[223])^(a[17] & b[224])^(a[16] & b[225])^(a[15] & b[226])^(a[14] & b[227])^(a[13] & b[228])^(a[12] & b[229])^(a[11] & b[230])^(a[10] & b[231])^(a[9] & b[232]);
assign y[242] = (a[232] & b[10])^(a[231] & b[11])^(a[230] & b[12])^(a[229] & b[13])^(a[228] & b[14])^(a[227] & b[15])^(a[226] & b[16])^(a[225] & b[17])^(a[224] & b[18])^(a[223] & b[19])^(a[222] & b[20])^(a[221] & b[21])^(a[220] & b[22])^(a[219] & b[23])^(a[218] & b[24])^(a[217] & b[25])^(a[216] & b[26])^(a[215] & b[27])^(a[214] & b[28])^(a[213] & b[29])^(a[212] & b[30])^(a[211] & b[31])^(a[210] & b[32])^(a[209] & b[33])^(a[208] & b[34])^(a[207] & b[35])^(a[206] & b[36])^(a[205] & b[37])^(a[204] & b[38])^(a[203] & b[39])^(a[202] & b[40])^(a[201] & b[41])^(a[200] & b[42])^(a[199] & b[43])^(a[198] & b[44])^(a[197] & b[45])^(a[196] & b[46])^(a[195] & b[47])^(a[194] & b[48])^(a[193] & b[49])^(a[192] & b[50])^(a[191] & b[51])^(a[190] & b[52])^(a[189] & b[53])^(a[188] & b[54])^(a[187] & b[55])^(a[186] & b[56])^(a[185] & b[57])^(a[184] & b[58])^(a[183] & b[59])^(a[182] & b[60])^(a[181] & b[61])^(a[180] & b[62])^(a[179] & b[63])^(a[178] & b[64])^(a[177] & b[65])^(a[176] & b[66])^(a[175] & b[67])^(a[174] & b[68])^(a[173] & b[69])^(a[172] & b[70])^(a[171] & b[71])^(a[170] & b[72])^(a[169] & b[73])^(a[168] & b[74])^(a[167] & b[75])^(a[166] & b[76])^(a[165] & b[77])^(a[164] & b[78])^(a[163] & b[79])^(a[162] & b[80])^(a[161] & b[81])^(a[160] & b[82])^(a[159] & b[83])^(a[158] & b[84])^(a[157] & b[85])^(a[156] & b[86])^(a[155] & b[87])^(a[154] & b[88])^(a[153] & b[89])^(a[152] & b[90])^(a[151] & b[91])^(a[150] & b[92])^(a[149] & b[93])^(a[148] & b[94])^(a[147] & b[95])^(a[146] & b[96])^(a[145] & b[97])^(a[144] & b[98])^(a[143] & b[99])^(a[142] & b[100])^(a[141] & b[101])^(a[140] & b[102])^(a[139] & b[103])^(a[138] & b[104])^(a[137] & b[105])^(a[136] & b[106])^(a[135] & b[107])^(a[134] & b[108])^(a[133] & b[109])^(a[132] & b[110])^(a[131] & b[111])^(a[130] & b[112])^(a[129] & b[113])^(a[128] & b[114])^(a[127] & b[115])^(a[126] & b[116])^(a[125] & b[117])^(a[124] & b[118])^(a[123] & b[119])^(a[122] & b[120])^(a[121] & b[121])^(a[120] & b[122])^(a[119] & b[123])^(a[118] & b[124])^(a[117] & b[125])^(a[116] & b[126])^(a[115] & b[127])^(a[114] & b[128])^(a[113] & b[129])^(a[112] & b[130])^(a[111] & b[131])^(a[110] & b[132])^(a[109] & b[133])^(a[108] & b[134])^(a[107] & b[135])^(a[106] & b[136])^(a[105] & b[137])^(a[104] & b[138])^(a[103] & b[139])^(a[102] & b[140])^(a[101] & b[141])^(a[100] & b[142])^(a[99] & b[143])^(a[98] & b[144])^(a[97] & b[145])^(a[96] & b[146])^(a[95] & b[147])^(a[94] & b[148])^(a[93] & b[149])^(a[92] & b[150])^(a[91] & b[151])^(a[90] & b[152])^(a[89] & b[153])^(a[88] & b[154])^(a[87] & b[155])^(a[86] & b[156])^(a[85] & b[157])^(a[84] & b[158])^(a[83] & b[159])^(a[82] & b[160])^(a[81] & b[161])^(a[80] & b[162])^(a[79] & b[163])^(a[78] & b[164])^(a[77] & b[165])^(a[76] & b[166])^(a[75] & b[167])^(a[74] & b[168])^(a[73] & b[169])^(a[72] & b[170])^(a[71] & b[171])^(a[70] & b[172])^(a[69] & b[173])^(a[68] & b[174])^(a[67] & b[175])^(a[66] & b[176])^(a[65] & b[177])^(a[64] & b[178])^(a[63] & b[179])^(a[62] & b[180])^(a[61] & b[181])^(a[60] & b[182])^(a[59] & b[183])^(a[58] & b[184])^(a[57] & b[185])^(a[56] & b[186])^(a[55] & b[187])^(a[54] & b[188])^(a[53] & b[189])^(a[52] & b[190])^(a[51] & b[191])^(a[50] & b[192])^(a[49] & b[193])^(a[48] & b[194])^(a[47] & b[195])^(a[46] & b[196])^(a[45] & b[197])^(a[44] & b[198])^(a[43] & b[199])^(a[42] & b[200])^(a[41] & b[201])^(a[40] & b[202])^(a[39] & b[203])^(a[38] & b[204])^(a[37] & b[205])^(a[36] & b[206])^(a[35] & b[207])^(a[34] & b[208])^(a[33] & b[209])^(a[32] & b[210])^(a[31] & b[211])^(a[30] & b[212])^(a[29] & b[213])^(a[28] & b[214])^(a[27] & b[215])^(a[26] & b[216])^(a[25] & b[217])^(a[24] & b[218])^(a[23] & b[219])^(a[22] & b[220])^(a[21] & b[221])^(a[20] & b[222])^(a[19] & b[223])^(a[18] & b[224])^(a[17] & b[225])^(a[16] & b[226])^(a[15] & b[227])^(a[14] & b[228])^(a[13] & b[229])^(a[12] & b[230])^(a[11] & b[231])^(a[10] & b[232]);
assign y[243] = (a[232] & b[11])^(a[231] & b[12])^(a[230] & b[13])^(a[229] & b[14])^(a[228] & b[15])^(a[227] & b[16])^(a[226] & b[17])^(a[225] & b[18])^(a[224] & b[19])^(a[223] & b[20])^(a[222] & b[21])^(a[221] & b[22])^(a[220] & b[23])^(a[219] & b[24])^(a[218] & b[25])^(a[217] & b[26])^(a[216] & b[27])^(a[215] & b[28])^(a[214] & b[29])^(a[213] & b[30])^(a[212] & b[31])^(a[211] & b[32])^(a[210] & b[33])^(a[209] & b[34])^(a[208] & b[35])^(a[207] & b[36])^(a[206] & b[37])^(a[205] & b[38])^(a[204] & b[39])^(a[203] & b[40])^(a[202] & b[41])^(a[201] & b[42])^(a[200] & b[43])^(a[199] & b[44])^(a[198] & b[45])^(a[197] & b[46])^(a[196] & b[47])^(a[195] & b[48])^(a[194] & b[49])^(a[193] & b[50])^(a[192] & b[51])^(a[191] & b[52])^(a[190] & b[53])^(a[189] & b[54])^(a[188] & b[55])^(a[187] & b[56])^(a[186] & b[57])^(a[185] & b[58])^(a[184] & b[59])^(a[183] & b[60])^(a[182] & b[61])^(a[181] & b[62])^(a[180] & b[63])^(a[179] & b[64])^(a[178] & b[65])^(a[177] & b[66])^(a[176] & b[67])^(a[175] & b[68])^(a[174] & b[69])^(a[173] & b[70])^(a[172] & b[71])^(a[171] & b[72])^(a[170] & b[73])^(a[169] & b[74])^(a[168] & b[75])^(a[167] & b[76])^(a[166] & b[77])^(a[165] & b[78])^(a[164] & b[79])^(a[163] & b[80])^(a[162] & b[81])^(a[161] & b[82])^(a[160] & b[83])^(a[159] & b[84])^(a[158] & b[85])^(a[157] & b[86])^(a[156] & b[87])^(a[155] & b[88])^(a[154] & b[89])^(a[153] & b[90])^(a[152] & b[91])^(a[151] & b[92])^(a[150] & b[93])^(a[149] & b[94])^(a[148] & b[95])^(a[147] & b[96])^(a[146] & b[97])^(a[145] & b[98])^(a[144] & b[99])^(a[143] & b[100])^(a[142] & b[101])^(a[141] & b[102])^(a[140] & b[103])^(a[139] & b[104])^(a[138] & b[105])^(a[137] & b[106])^(a[136] & b[107])^(a[135] & b[108])^(a[134] & b[109])^(a[133] & b[110])^(a[132] & b[111])^(a[131] & b[112])^(a[130] & b[113])^(a[129] & b[114])^(a[128] & b[115])^(a[127] & b[116])^(a[126] & b[117])^(a[125] & b[118])^(a[124] & b[119])^(a[123] & b[120])^(a[122] & b[121])^(a[121] & b[122])^(a[120] & b[123])^(a[119] & b[124])^(a[118] & b[125])^(a[117] & b[126])^(a[116] & b[127])^(a[115] & b[128])^(a[114] & b[129])^(a[113] & b[130])^(a[112] & b[131])^(a[111] & b[132])^(a[110] & b[133])^(a[109] & b[134])^(a[108] & b[135])^(a[107] & b[136])^(a[106] & b[137])^(a[105] & b[138])^(a[104] & b[139])^(a[103] & b[140])^(a[102] & b[141])^(a[101] & b[142])^(a[100] & b[143])^(a[99] & b[144])^(a[98] & b[145])^(a[97] & b[146])^(a[96] & b[147])^(a[95] & b[148])^(a[94] & b[149])^(a[93] & b[150])^(a[92] & b[151])^(a[91] & b[152])^(a[90] & b[153])^(a[89] & b[154])^(a[88] & b[155])^(a[87] & b[156])^(a[86] & b[157])^(a[85] & b[158])^(a[84] & b[159])^(a[83] & b[160])^(a[82] & b[161])^(a[81] & b[162])^(a[80] & b[163])^(a[79] & b[164])^(a[78] & b[165])^(a[77] & b[166])^(a[76] & b[167])^(a[75] & b[168])^(a[74] & b[169])^(a[73] & b[170])^(a[72] & b[171])^(a[71] & b[172])^(a[70] & b[173])^(a[69] & b[174])^(a[68] & b[175])^(a[67] & b[176])^(a[66] & b[177])^(a[65] & b[178])^(a[64] & b[179])^(a[63] & b[180])^(a[62] & b[181])^(a[61] & b[182])^(a[60] & b[183])^(a[59] & b[184])^(a[58] & b[185])^(a[57] & b[186])^(a[56] & b[187])^(a[55] & b[188])^(a[54] & b[189])^(a[53] & b[190])^(a[52] & b[191])^(a[51] & b[192])^(a[50] & b[193])^(a[49] & b[194])^(a[48] & b[195])^(a[47] & b[196])^(a[46] & b[197])^(a[45] & b[198])^(a[44] & b[199])^(a[43] & b[200])^(a[42] & b[201])^(a[41] & b[202])^(a[40] & b[203])^(a[39] & b[204])^(a[38] & b[205])^(a[37] & b[206])^(a[36] & b[207])^(a[35] & b[208])^(a[34] & b[209])^(a[33] & b[210])^(a[32] & b[211])^(a[31] & b[212])^(a[30] & b[213])^(a[29] & b[214])^(a[28] & b[215])^(a[27] & b[216])^(a[26] & b[217])^(a[25] & b[218])^(a[24] & b[219])^(a[23] & b[220])^(a[22] & b[221])^(a[21] & b[222])^(a[20] & b[223])^(a[19] & b[224])^(a[18] & b[225])^(a[17] & b[226])^(a[16] & b[227])^(a[15] & b[228])^(a[14] & b[229])^(a[13] & b[230])^(a[12] & b[231])^(a[11] & b[232]);
assign y[244] = (a[232] & b[12])^(a[231] & b[13])^(a[230] & b[14])^(a[229] & b[15])^(a[228] & b[16])^(a[227] & b[17])^(a[226] & b[18])^(a[225] & b[19])^(a[224] & b[20])^(a[223] & b[21])^(a[222] & b[22])^(a[221] & b[23])^(a[220] & b[24])^(a[219] & b[25])^(a[218] & b[26])^(a[217] & b[27])^(a[216] & b[28])^(a[215] & b[29])^(a[214] & b[30])^(a[213] & b[31])^(a[212] & b[32])^(a[211] & b[33])^(a[210] & b[34])^(a[209] & b[35])^(a[208] & b[36])^(a[207] & b[37])^(a[206] & b[38])^(a[205] & b[39])^(a[204] & b[40])^(a[203] & b[41])^(a[202] & b[42])^(a[201] & b[43])^(a[200] & b[44])^(a[199] & b[45])^(a[198] & b[46])^(a[197] & b[47])^(a[196] & b[48])^(a[195] & b[49])^(a[194] & b[50])^(a[193] & b[51])^(a[192] & b[52])^(a[191] & b[53])^(a[190] & b[54])^(a[189] & b[55])^(a[188] & b[56])^(a[187] & b[57])^(a[186] & b[58])^(a[185] & b[59])^(a[184] & b[60])^(a[183] & b[61])^(a[182] & b[62])^(a[181] & b[63])^(a[180] & b[64])^(a[179] & b[65])^(a[178] & b[66])^(a[177] & b[67])^(a[176] & b[68])^(a[175] & b[69])^(a[174] & b[70])^(a[173] & b[71])^(a[172] & b[72])^(a[171] & b[73])^(a[170] & b[74])^(a[169] & b[75])^(a[168] & b[76])^(a[167] & b[77])^(a[166] & b[78])^(a[165] & b[79])^(a[164] & b[80])^(a[163] & b[81])^(a[162] & b[82])^(a[161] & b[83])^(a[160] & b[84])^(a[159] & b[85])^(a[158] & b[86])^(a[157] & b[87])^(a[156] & b[88])^(a[155] & b[89])^(a[154] & b[90])^(a[153] & b[91])^(a[152] & b[92])^(a[151] & b[93])^(a[150] & b[94])^(a[149] & b[95])^(a[148] & b[96])^(a[147] & b[97])^(a[146] & b[98])^(a[145] & b[99])^(a[144] & b[100])^(a[143] & b[101])^(a[142] & b[102])^(a[141] & b[103])^(a[140] & b[104])^(a[139] & b[105])^(a[138] & b[106])^(a[137] & b[107])^(a[136] & b[108])^(a[135] & b[109])^(a[134] & b[110])^(a[133] & b[111])^(a[132] & b[112])^(a[131] & b[113])^(a[130] & b[114])^(a[129] & b[115])^(a[128] & b[116])^(a[127] & b[117])^(a[126] & b[118])^(a[125] & b[119])^(a[124] & b[120])^(a[123] & b[121])^(a[122] & b[122])^(a[121] & b[123])^(a[120] & b[124])^(a[119] & b[125])^(a[118] & b[126])^(a[117] & b[127])^(a[116] & b[128])^(a[115] & b[129])^(a[114] & b[130])^(a[113] & b[131])^(a[112] & b[132])^(a[111] & b[133])^(a[110] & b[134])^(a[109] & b[135])^(a[108] & b[136])^(a[107] & b[137])^(a[106] & b[138])^(a[105] & b[139])^(a[104] & b[140])^(a[103] & b[141])^(a[102] & b[142])^(a[101] & b[143])^(a[100] & b[144])^(a[99] & b[145])^(a[98] & b[146])^(a[97] & b[147])^(a[96] & b[148])^(a[95] & b[149])^(a[94] & b[150])^(a[93] & b[151])^(a[92] & b[152])^(a[91] & b[153])^(a[90] & b[154])^(a[89] & b[155])^(a[88] & b[156])^(a[87] & b[157])^(a[86] & b[158])^(a[85] & b[159])^(a[84] & b[160])^(a[83] & b[161])^(a[82] & b[162])^(a[81] & b[163])^(a[80] & b[164])^(a[79] & b[165])^(a[78] & b[166])^(a[77] & b[167])^(a[76] & b[168])^(a[75] & b[169])^(a[74] & b[170])^(a[73] & b[171])^(a[72] & b[172])^(a[71] & b[173])^(a[70] & b[174])^(a[69] & b[175])^(a[68] & b[176])^(a[67] & b[177])^(a[66] & b[178])^(a[65] & b[179])^(a[64] & b[180])^(a[63] & b[181])^(a[62] & b[182])^(a[61] & b[183])^(a[60] & b[184])^(a[59] & b[185])^(a[58] & b[186])^(a[57] & b[187])^(a[56] & b[188])^(a[55] & b[189])^(a[54] & b[190])^(a[53] & b[191])^(a[52] & b[192])^(a[51] & b[193])^(a[50] & b[194])^(a[49] & b[195])^(a[48] & b[196])^(a[47] & b[197])^(a[46] & b[198])^(a[45] & b[199])^(a[44] & b[200])^(a[43] & b[201])^(a[42] & b[202])^(a[41] & b[203])^(a[40] & b[204])^(a[39] & b[205])^(a[38] & b[206])^(a[37] & b[207])^(a[36] & b[208])^(a[35] & b[209])^(a[34] & b[210])^(a[33] & b[211])^(a[32] & b[212])^(a[31] & b[213])^(a[30] & b[214])^(a[29] & b[215])^(a[28] & b[216])^(a[27] & b[217])^(a[26] & b[218])^(a[25] & b[219])^(a[24] & b[220])^(a[23] & b[221])^(a[22] & b[222])^(a[21] & b[223])^(a[20] & b[224])^(a[19] & b[225])^(a[18] & b[226])^(a[17] & b[227])^(a[16] & b[228])^(a[15] & b[229])^(a[14] & b[230])^(a[13] & b[231])^(a[12] & b[232]);
assign y[245] = (a[232] & b[13])^(a[231] & b[14])^(a[230] & b[15])^(a[229] & b[16])^(a[228] & b[17])^(a[227] & b[18])^(a[226] & b[19])^(a[225] & b[20])^(a[224] & b[21])^(a[223] & b[22])^(a[222] & b[23])^(a[221] & b[24])^(a[220] & b[25])^(a[219] & b[26])^(a[218] & b[27])^(a[217] & b[28])^(a[216] & b[29])^(a[215] & b[30])^(a[214] & b[31])^(a[213] & b[32])^(a[212] & b[33])^(a[211] & b[34])^(a[210] & b[35])^(a[209] & b[36])^(a[208] & b[37])^(a[207] & b[38])^(a[206] & b[39])^(a[205] & b[40])^(a[204] & b[41])^(a[203] & b[42])^(a[202] & b[43])^(a[201] & b[44])^(a[200] & b[45])^(a[199] & b[46])^(a[198] & b[47])^(a[197] & b[48])^(a[196] & b[49])^(a[195] & b[50])^(a[194] & b[51])^(a[193] & b[52])^(a[192] & b[53])^(a[191] & b[54])^(a[190] & b[55])^(a[189] & b[56])^(a[188] & b[57])^(a[187] & b[58])^(a[186] & b[59])^(a[185] & b[60])^(a[184] & b[61])^(a[183] & b[62])^(a[182] & b[63])^(a[181] & b[64])^(a[180] & b[65])^(a[179] & b[66])^(a[178] & b[67])^(a[177] & b[68])^(a[176] & b[69])^(a[175] & b[70])^(a[174] & b[71])^(a[173] & b[72])^(a[172] & b[73])^(a[171] & b[74])^(a[170] & b[75])^(a[169] & b[76])^(a[168] & b[77])^(a[167] & b[78])^(a[166] & b[79])^(a[165] & b[80])^(a[164] & b[81])^(a[163] & b[82])^(a[162] & b[83])^(a[161] & b[84])^(a[160] & b[85])^(a[159] & b[86])^(a[158] & b[87])^(a[157] & b[88])^(a[156] & b[89])^(a[155] & b[90])^(a[154] & b[91])^(a[153] & b[92])^(a[152] & b[93])^(a[151] & b[94])^(a[150] & b[95])^(a[149] & b[96])^(a[148] & b[97])^(a[147] & b[98])^(a[146] & b[99])^(a[145] & b[100])^(a[144] & b[101])^(a[143] & b[102])^(a[142] & b[103])^(a[141] & b[104])^(a[140] & b[105])^(a[139] & b[106])^(a[138] & b[107])^(a[137] & b[108])^(a[136] & b[109])^(a[135] & b[110])^(a[134] & b[111])^(a[133] & b[112])^(a[132] & b[113])^(a[131] & b[114])^(a[130] & b[115])^(a[129] & b[116])^(a[128] & b[117])^(a[127] & b[118])^(a[126] & b[119])^(a[125] & b[120])^(a[124] & b[121])^(a[123] & b[122])^(a[122] & b[123])^(a[121] & b[124])^(a[120] & b[125])^(a[119] & b[126])^(a[118] & b[127])^(a[117] & b[128])^(a[116] & b[129])^(a[115] & b[130])^(a[114] & b[131])^(a[113] & b[132])^(a[112] & b[133])^(a[111] & b[134])^(a[110] & b[135])^(a[109] & b[136])^(a[108] & b[137])^(a[107] & b[138])^(a[106] & b[139])^(a[105] & b[140])^(a[104] & b[141])^(a[103] & b[142])^(a[102] & b[143])^(a[101] & b[144])^(a[100] & b[145])^(a[99] & b[146])^(a[98] & b[147])^(a[97] & b[148])^(a[96] & b[149])^(a[95] & b[150])^(a[94] & b[151])^(a[93] & b[152])^(a[92] & b[153])^(a[91] & b[154])^(a[90] & b[155])^(a[89] & b[156])^(a[88] & b[157])^(a[87] & b[158])^(a[86] & b[159])^(a[85] & b[160])^(a[84] & b[161])^(a[83] & b[162])^(a[82] & b[163])^(a[81] & b[164])^(a[80] & b[165])^(a[79] & b[166])^(a[78] & b[167])^(a[77] & b[168])^(a[76] & b[169])^(a[75] & b[170])^(a[74] & b[171])^(a[73] & b[172])^(a[72] & b[173])^(a[71] & b[174])^(a[70] & b[175])^(a[69] & b[176])^(a[68] & b[177])^(a[67] & b[178])^(a[66] & b[179])^(a[65] & b[180])^(a[64] & b[181])^(a[63] & b[182])^(a[62] & b[183])^(a[61] & b[184])^(a[60] & b[185])^(a[59] & b[186])^(a[58] & b[187])^(a[57] & b[188])^(a[56] & b[189])^(a[55] & b[190])^(a[54] & b[191])^(a[53] & b[192])^(a[52] & b[193])^(a[51] & b[194])^(a[50] & b[195])^(a[49] & b[196])^(a[48] & b[197])^(a[47] & b[198])^(a[46] & b[199])^(a[45] & b[200])^(a[44] & b[201])^(a[43] & b[202])^(a[42] & b[203])^(a[41] & b[204])^(a[40] & b[205])^(a[39] & b[206])^(a[38] & b[207])^(a[37] & b[208])^(a[36] & b[209])^(a[35] & b[210])^(a[34] & b[211])^(a[33] & b[212])^(a[32] & b[213])^(a[31] & b[214])^(a[30] & b[215])^(a[29] & b[216])^(a[28] & b[217])^(a[27] & b[218])^(a[26] & b[219])^(a[25] & b[220])^(a[24] & b[221])^(a[23] & b[222])^(a[22] & b[223])^(a[21] & b[224])^(a[20] & b[225])^(a[19] & b[226])^(a[18] & b[227])^(a[17] & b[228])^(a[16] & b[229])^(a[15] & b[230])^(a[14] & b[231])^(a[13] & b[232]);
assign y[246] = (a[232] & b[14])^(a[231] & b[15])^(a[230] & b[16])^(a[229] & b[17])^(a[228] & b[18])^(a[227] & b[19])^(a[226] & b[20])^(a[225] & b[21])^(a[224] & b[22])^(a[223] & b[23])^(a[222] & b[24])^(a[221] & b[25])^(a[220] & b[26])^(a[219] & b[27])^(a[218] & b[28])^(a[217] & b[29])^(a[216] & b[30])^(a[215] & b[31])^(a[214] & b[32])^(a[213] & b[33])^(a[212] & b[34])^(a[211] & b[35])^(a[210] & b[36])^(a[209] & b[37])^(a[208] & b[38])^(a[207] & b[39])^(a[206] & b[40])^(a[205] & b[41])^(a[204] & b[42])^(a[203] & b[43])^(a[202] & b[44])^(a[201] & b[45])^(a[200] & b[46])^(a[199] & b[47])^(a[198] & b[48])^(a[197] & b[49])^(a[196] & b[50])^(a[195] & b[51])^(a[194] & b[52])^(a[193] & b[53])^(a[192] & b[54])^(a[191] & b[55])^(a[190] & b[56])^(a[189] & b[57])^(a[188] & b[58])^(a[187] & b[59])^(a[186] & b[60])^(a[185] & b[61])^(a[184] & b[62])^(a[183] & b[63])^(a[182] & b[64])^(a[181] & b[65])^(a[180] & b[66])^(a[179] & b[67])^(a[178] & b[68])^(a[177] & b[69])^(a[176] & b[70])^(a[175] & b[71])^(a[174] & b[72])^(a[173] & b[73])^(a[172] & b[74])^(a[171] & b[75])^(a[170] & b[76])^(a[169] & b[77])^(a[168] & b[78])^(a[167] & b[79])^(a[166] & b[80])^(a[165] & b[81])^(a[164] & b[82])^(a[163] & b[83])^(a[162] & b[84])^(a[161] & b[85])^(a[160] & b[86])^(a[159] & b[87])^(a[158] & b[88])^(a[157] & b[89])^(a[156] & b[90])^(a[155] & b[91])^(a[154] & b[92])^(a[153] & b[93])^(a[152] & b[94])^(a[151] & b[95])^(a[150] & b[96])^(a[149] & b[97])^(a[148] & b[98])^(a[147] & b[99])^(a[146] & b[100])^(a[145] & b[101])^(a[144] & b[102])^(a[143] & b[103])^(a[142] & b[104])^(a[141] & b[105])^(a[140] & b[106])^(a[139] & b[107])^(a[138] & b[108])^(a[137] & b[109])^(a[136] & b[110])^(a[135] & b[111])^(a[134] & b[112])^(a[133] & b[113])^(a[132] & b[114])^(a[131] & b[115])^(a[130] & b[116])^(a[129] & b[117])^(a[128] & b[118])^(a[127] & b[119])^(a[126] & b[120])^(a[125] & b[121])^(a[124] & b[122])^(a[123] & b[123])^(a[122] & b[124])^(a[121] & b[125])^(a[120] & b[126])^(a[119] & b[127])^(a[118] & b[128])^(a[117] & b[129])^(a[116] & b[130])^(a[115] & b[131])^(a[114] & b[132])^(a[113] & b[133])^(a[112] & b[134])^(a[111] & b[135])^(a[110] & b[136])^(a[109] & b[137])^(a[108] & b[138])^(a[107] & b[139])^(a[106] & b[140])^(a[105] & b[141])^(a[104] & b[142])^(a[103] & b[143])^(a[102] & b[144])^(a[101] & b[145])^(a[100] & b[146])^(a[99] & b[147])^(a[98] & b[148])^(a[97] & b[149])^(a[96] & b[150])^(a[95] & b[151])^(a[94] & b[152])^(a[93] & b[153])^(a[92] & b[154])^(a[91] & b[155])^(a[90] & b[156])^(a[89] & b[157])^(a[88] & b[158])^(a[87] & b[159])^(a[86] & b[160])^(a[85] & b[161])^(a[84] & b[162])^(a[83] & b[163])^(a[82] & b[164])^(a[81] & b[165])^(a[80] & b[166])^(a[79] & b[167])^(a[78] & b[168])^(a[77] & b[169])^(a[76] & b[170])^(a[75] & b[171])^(a[74] & b[172])^(a[73] & b[173])^(a[72] & b[174])^(a[71] & b[175])^(a[70] & b[176])^(a[69] & b[177])^(a[68] & b[178])^(a[67] & b[179])^(a[66] & b[180])^(a[65] & b[181])^(a[64] & b[182])^(a[63] & b[183])^(a[62] & b[184])^(a[61] & b[185])^(a[60] & b[186])^(a[59] & b[187])^(a[58] & b[188])^(a[57] & b[189])^(a[56] & b[190])^(a[55] & b[191])^(a[54] & b[192])^(a[53] & b[193])^(a[52] & b[194])^(a[51] & b[195])^(a[50] & b[196])^(a[49] & b[197])^(a[48] & b[198])^(a[47] & b[199])^(a[46] & b[200])^(a[45] & b[201])^(a[44] & b[202])^(a[43] & b[203])^(a[42] & b[204])^(a[41] & b[205])^(a[40] & b[206])^(a[39] & b[207])^(a[38] & b[208])^(a[37] & b[209])^(a[36] & b[210])^(a[35] & b[211])^(a[34] & b[212])^(a[33] & b[213])^(a[32] & b[214])^(a[31] & b[215])^(a[30] & b[216])^(a[29] & b[217])^(a[28] & b[218])^(a[27] & b[219])^(a[26] & b[220])^(a[25] & b[221])^(a[24] & b[222])^(a[23] & b[223])^(a[22] & b[224])^(a[21] & b[225])^(a[20] & b[226])^(a[19] & b[227])^(a[18] & b[228])^(a[17] & b[229])^(a[16] & b[230])^(a[15] & b[231])^(a[14] & b[232]);
assign y[247] = (a[232] & b[15])^(a[231] & b[16])^(a[230] & b[17])^(a[229] & b[18])^(a[228] & b[19])^(a[227] & b[20])^(a[226] & b[21])^(a[225] & b[22])^(a[224] & b[23])^(a[223] & b[24])^(a[222] & b[25])^(a[221] & b[26])^(a[220] & b[27])^(a[219] & b[28])^(a[218] & b[29])^(a[217] & b[30])^(a[216] & b[31])^(a[215] & b[32])^(a[214] & b[33])^(a[213] & b[34])^(a[212] & b[35])^(a[211] & b[36])^(a[210] & b[37])^(a[209] & b[38])^(a[208] & b[39])^(a[207] & b[40])^(a[206] & b[41])^(a[205] & b[42])^(a[204] & b[43])^(a[203] & b[44])^(a[202] & b[45])^(a[201] & b[46])^(a[200] & b[47])^(a[199] & b[48])^(a[198] & b[49])^(a[197] & b[50])^(a[196] & b[51])^(a[195] & b[52])^(a[194] & b[53])^(a[193] & b[54])^(a[192] & b[55])^(a[191] & b[56])^(a[190] & b[57])^(a[189] & b[58])^(a[188] & b[59])^(a[187] & b[60])^(a[186] & b[61])^(a[185] & b[62])^(a[184] & b[63])^(a[183] & b[64])^(a[182] & b[65])^(a[181] & b[66])^(a[180] & b[67])^(a[179] & b[68])^(a[178] & b[69])^(a[177] & b[70])^(a[176] & b[71])^(a[175] & b[72])^(a[174] & b[73])^(a[173] & b[74])^(a[172] & b[75])^(a[171] & b[76])^(a[170] & b[77])^(a[169] & b[78])^(a[168] & b[79])^(a[167] & b[80])^(a[166] & b[81])^(a[165] & b[82])^(a[164] & b[83])^(a[163] & b[84])^(a[162] & b[85])^(a[161] & b[86])^(a[160] & b[87])^(a[159] & b[88])^(a[158] & b[89])^(a[157] & b[90])^(a[156] & b[91])^(a[155] & b[92])^(a[154] & b[93])^(a[153] & b[94])^(a[152] & b[95])^(a[151] & b[96])^(a[150] & b[97])^(a[149] & b[98])^(a[148] & b[99])^(a[147] & b[100])^(a[146] & b[101])^(a[145] & b[102])^(a[144] & b[103])^(a[143] & b[104])^(a[142] & b[105])^(a[141] & b[106])^(a[140] & b[107])^(a[139] & b[108])^(a[138] & b[109])^(a[137] & b[110])^(a[136] & b[111])^(a[135] & b[112])^(a[134] & b[113])^(a[133] & b[114])^(a[132] & b[115])^(a[131] & b[116])^(a[130] & b[117])^(a[129] & b[118])^(a[128] & b[119])^(a[127] & b[120])^(a[126] & b[121])^(a[125] & b[122])^(a[124] & b[123])^(a[123] & b[124])^(a[122] & b[125])^(a[121] & b[126])^(a[120] & b[127])^(a[119] & b[128])^(a[118] & b[129])^(a[117] & b[130])^(a[116] & b[131])^(a[115] & b[132])^(a[114] & b[133])^(a[113] & b[134])^(a[112] & b[135])^(a[111] & b[136])^(a[110] & b[137])^(a[109] & b[138])^(a[108] & b[139])^(a[107] & b[140])^(a[106] & b[141])^(a[105] & b[142])^(a[104] & b[143])^(a[103] & b[144])^(a[102] & b[145])^(a[101] & b[146])^(a[100] & b[147])^(a[99] & b[148])^(a[98] & b[149])^(a[97] & b[150])^(a[96] & b[151])^(a[95] & b[152])^(a[94] & b[153])^(a[93] & b[154])^(a[92] & b[155])^(a[91] & b[156])^(a[90] & b[157])^(a[89] & b[158])^(a[88] & b[159])^(a[87] & b[160])^(a[86] & b[161])^(a[85] & b[162])^(a[84] & b[163])^(a[83] & b[164])^(a[82] & b[165])^(a[81] & b[166])^(a[80] & b[167])^(a[79] & b[168])^(a[78] & b[169])^(a[77] & b[170])^(a[76] & b[171])^(a[75] & b[172])^(a[74] & b[173])^(a[73] & b[174])^(a[72] & b[175])^(a[71] & b[176])^(a[70] & b[177])^(a[69] & b[178])^(a[68] & b[179])^(a[67] & b[180])^(a[66] & b[181])^(a[65] & b[182])^(a[64] & b[183])^(a[63] & b[184])^(a[62] & b[185])^(a[61] & b[186])^(a[60] & b[187])^(a[59] & b[188])^(a[58] & b[189])^(a[57] & b[190])^(a[56] & b[191])^(a[55] & b[192])^(a[54] & b[193])^(a[53] & b[194])^(a[52] & b[195])^(a[51] & b[196])^(a[50] & b[197])^(a[49] & b[198])^(a[48] & b[199])^(a[47] & b[200])^(a[46] & b[201])^(a[45] & b[202])^(a[44] & b[203])^(a[43] & b[204])^(a[42] & b[205])^(a[41] & b[206])^(a[40] & b[207])^(a[39] & b[208])^(a[38] & b[209])^(a[37] & b[210])^(a[36] & b[211])^(a[35] & b[212])^(a[34] & b[213])^(a[33] & b[214])^(a[32] & b[215])^(a[31] & b[216])^(a[30] & b[217])^(a[29] & b[218])^(a[28] & b[219])^(a[27] & b[220])^(a[26] & b[221])^(a[25] & b[222])^(a[24] & b[223])^(a[23] & b[224])^(a[22] & b[225])^(a[21] & b[226])^(a[20] & b[227])^(a[19] & b[228])^(a[18] & b[229])^(a[17] & b[230])^(a[16] & b[231])^(a[15] & b[232]);
assign y[248] = (a[232] & b[16])^(a[231] & b[17])^(a[230] & b[18])^(a[229] & b[19])^(a[228] & b[20])^(a[227] & b[21])^(a[226] & b[22])^(a[225] & b[23])^(a[224] & b[24])^(a[223] & b[25])^(a[222] & b[26])^(a[221] & b[27])^(a[220] & b[28])^(a[219] & b[29])^(a[218] & b[30])^(a[217] & b[31])^(a[216] & b[32])^(a[215] & b[33])^(a[214] & b[34])^(a[213] & b[35])^(a[212] & b[36])^(a[211] & b[37])^(a[210] & b[38])^(a[209] & b[39])^(a[208] & b[40])^(a[207] & b[41])^(a[206] & b[42])^(a[205] & b[43])^(a[204] & b[44])^(a[203] & b[45])^(a[202] & b[46])^(a[201] & b[47])^(a[200] & b[48])^(a[199] & b[49])^(a[198] & b[50])^(a[197] & b[51])^(a[196] & b[52])^(a[195] & b[53])^(a[194] & b[54])^(a[193] & b[55])^(a[192] & b[56])^(a[191] & b[57])^(a[190] & b[58])^(a[189] & b[59])^(a[188] & b[60])^(a[187] & b[61])^(a[186] & b[62])^(a[185] & b[63])^(a[184] & b[64])^(a[183] & b[65])^(a[182] & b[66])^(a[181] & b[67])^(a[180] & b[68])^(a[179] & b[69])^(a[178] & b[70])^(a[177] & b[71])^(a[176] & b[72])^(a[175] & b[73])^(a[174] & b[74])^(a[173] & b[75])^(a[172] & b[76])^(a[171] & b[77])^(a[170] & b[78])^(a[169] & b[79])^(a[168] & b[80])^(a[167] & b[81])^(a[166] & b[82])^(a[165] & b[83])^(a[164] & b[84])^(a[163] & b[85])^(a[162] & b[86])^(a[161] & b[87])^(a[160] & b[88])^(a[159] & b[89])^(a[158] & b[90])^(a[157] & b[91])^(a[156] & b[92])^(a[155] & b[93])^(a[154] & b[94])^(a[153] & b[95])^(a[152] & b[96])^(a[151] & b[97])^(a[150] & b[98])^(a[149] & b[99])^(a[148] & b[100])^(a[147] & b[101])^(a[146] & b[102])^(a[145] & b[103])^(a[144] & b[104])^(a[143] & b[105])^(a[142] & b[106])^(a[141] & b[107])^(a[140] & b[108])^(a[139] & b[109])^(a[138] & b[110])^(a[137] & b[111])^(a[136] & b[112])^(a[135] & b[113])^(a[134] & b[114])^(a[133] & b[115])^(a[132] & b[116])^(a[131] & b[117])^(a[130] & b[118])^(a[129] & b[119])^(a[128] & b[120])^(a[127] & b[121])^(a[126] & b[122])^(a[125] & b[123])^(a[124] & b[124])^(a[123] & b[125])^(a[122] & b[126])^(a[121] & b[127])^(a[120] & b[128])^(a[119] & b[129])^(a[118] & b[130])^(a[117] & b[131])^(a[116] & b[132])^(a[115] & b[133])^(a[114] & b[134])^(a[113] & b[135])^(a[112] & b[136])^(a[111] & b[137])^(a[110] & b[138])^(a[109] & b[139])^(a[108] & b[140])^(a[107] & b[141])^(a[106] & b[142])^(a[105] & b[143])^(a[104] & b[144])^(a[103] & b[145])^(a[102] & b[146])^(a[101] & b[147])^(a[100] & b[148])^(a[99] & b[149])^(a[98] & b[150])^(a[97] & b[151])^(a[96] & b[152])^(a[95] & b[153])^(a[94] & b[154])^(a[93] & b[155])^(a[92] & b[156])^(a[91] & b[157])^(a[90] & b[158])^(a[89] & b[159])^(a[88] & b[160])^(a[87] & b[161])^(a[86] & b[162])^(a[85] & b[163])^(a[84] & b[164])^(a[83] & b[165])^(a[82] & b[166])^(a[81] & b[167])^(a[80] & b[168])^(a[79] & b[169])^(a[78] & b[170])^(a[77] & b[171])^(a[76] & b[172])^(a[75] & b[173])^(a[74] & b[174])^(a[73] & b[175])^(a[72] & b[176])^(a[71] & b[177])^(a[70] & b[178])^(a[69] & b[179])^(a[68] & b[180])^(a[67] & b[181])^(a[66] & b[182])^(a[65] & b[183])^(a[64] & b[184])^(a[63] & b[185])^(a[62] & b[186])^(a[61] & b[187])^(a[60] & b[188])^(a[59] & b[189])^(a[58] & b[190])^(a[57] & b[191])^(a[56] & b[192])^(a[55] & b[193])^(a[54] & b[194])^(a[53] & b[195])^(a[52] & b[196])^(a[51] & b[197])^(a[50] & b[198])^(a[49] & b[199])^(a[48] & b[200])^(a[47] & b[201])^(a[46] & b[202])^(a[45] & b[203])^(a[44] & b[204])^(a[43] & b[205])^(a[42] & b[206])^(a[41] & b[207])^(a[40] & b[208])^(a[39] & b[209])^(a[38] & b[210])^(a[37] & b[211])^(a[36] & b[212])^(a[35] & b[213])^(a[34] & b[214])^(a[33] & b[215])^(a[32] & b[216])^(a[31] & b[217])^(a[30] & b[218])^(a[29] & b[219])^(a[28] & b[220])^(a[27] & b[221])^(a[26] & b[222])^(a[25] & b[223])^(a[24] & b[224])^(a[23] & b[225])^(a[22] & b[226])^(a[21] & b[227])^(a[20] & b[228])^(a[19] & b[229])^(a[18] & b[230])^(a[17] & b[231])^(a[16] & b[232]);
assign y[249] = (a[232] & b[17])^(a[231] & b[18])^(a[230] & b[19])^(a[229] & b[20])^(a[228] & b[21])^(a[227] & b[22])^(a[226] & b[23])^(a[225] & b[24])^(a[224] & b[25])^(a[223] & b[26])^(a[222] & b[27])^(a[221] & b[28])^(a[220] & b[29])^(a[219] & b[30])^(a[218] & b[31])^(a[217] & b[32])^(a[216] & b[33])^(a[215] & b[34])^(a[214] & b[35])^(a[213] & b[36])^(a[212] & b[37])^(a[211] & b[38])^(a[210] & b[39])^(a[209] & b[40])^(a[208] & b[41])^(a[207] & b[42])^(a[206] & b[43])^(a[205] & b[44])^(a[204] & b[45])^(a[203] & b[46])^(a[202] & b[47])^(a[201] & b[48])^(a[200] & b[49])^(a[199] & b[50])^(a[198] & b[51])^(a[197] & b[52])^(a[196] & b[53])^(a[195] & b[54])^(a[194] & b[55])^(a[193] & b[56])^(a[192] & b[57])^(a[191] & b[58])^(a[190] & b[59])^(a[189] & b[60])^(a[188] & b[61])^(a[187] & b[62])^(a[186] & b[63])^(a[185] & b[64])^(a[184] & b[65])^(a[183] & b[66])^(a[182] & b[67])^(a[181] & b[68])^(a[180] & b[69])^(a[179] & b[70])^(a[178] & b[71])^(a[177] & b[72])^(a[176] & b[73])^(a[175] & b[74])^(a[174] & b[75])^(a[173] & b[76])^(a[172] & b[77])^(a[171] & b[78])^(a[170] & b[79])^(a[169] & b[80])^(a[168] & b[81])^(a[167] & b[82])^(a[166] & b[83])^(a[165] & b[84])^(a[164] & b[85])^(a[163] & b[86])^(a[162] & b[87])^(a[161] & b[88])^(a[160] & b[89])^(a[159] & b[90])^(a[158] & b[91])^(a[157] & b[92])^(a[156] & b[93])^(a[155] & b[94])^(a[154] & b[95])^(a[153] & b[96])^(a[152] & b[97])^(a[151] & b[98])^(a[150] & b[99])^(a[149] & b[100])^(a[148] & b[101])^(a[147] & b[102])^(a[146] & b[103])^(a[145] & b[104])^(a[144] & b[105])^(a[143] & b[106])^(a[142] & b[107])^(a[141] & b[108])^(a[140] & b[109])^(a[139] & b[110])^(a[138] & b[111])^(a[137] & b[112])^(a[136] & b[113])^(a[135] & b[114])^(a[134] & b[115])^(a[133] & b[116])^(a[132] & b[117])^(a[131] & b[118])^(a[130] & b[119])^(a[129] & b[120])^(a[128] & b[121])^(a[127] & b[122])^(a[126] & b[123])^(a[125] & b[124])^(a[124] & b[125])^(a[123] & b[126])^(a[122] & b[127])^(a[121] & b[128])^(a[120] & b[129])^(a[119] & b[130])^(a[118] & b[131])^(a[117] & b[132])^(a[116] & b[133])^(a[115] & b[134])^(a[114] & b[135])^(a[113] & b[136])^(a[112] & b[137])^(a[111] & b[138])^(a[110] & b[139])^(a[109] & b[140])^(a[108] & b[141])^(a[107] & b[142])^(a[106] & b[143])^(a[105] & b[144])^(a[104] & b[145])^(a[103] & b[146])^(a[102] & b[147])^(a[101] & b[148])^(a[100] & b[149])^(a[99] & b[150])^(a[98] & b[151])^(a[97] & b[152])^(a[96] & b[153])^(a[95] & b[154])^(a[94] & b[155])^(a[93] & b[156])^(a[92] & b[157])^(a[91] & b[158])^(a[90] & b[159])^(a[89] & b[160])^(a[88] & b[161])^(a[87] & b[162])^(a[86] & b[163])^(a[85] & b[164])^(a[84] & b[165])^(a[83] & b[166])^(a[82] & b[167])^(a[81] & b[168])^(a[80] & b[169])^(a[79] & b[170])^(a[78] & b[171])^(a[77] & b[172])^(a[76] & b[173])^(a[75] & b[174])^(a[74] & b[175])^(a[73] & b[176])^(a[72] & b[177])^(a[71] & b[178])^(a[70] & b[179])^(a[69] & b[180])^(a[68] & b[181])^(a[67] & b[182])^(a[66] & b[183])^(a[65] & b[184])^(a[64] & b[185])^(a[63] & b[186])^(a[62] & b[187])^(a[61] & b[188])^(a[60] & b[189])^(a[59] & b[190])^(a[58] & b[191])^(a[57] & b[192])^(a[56] & b[193])^(a[55] & b[194])^(a[54] & b[195])^(a[53] & b[196])^(a[52] & b[197])^(a[51] & b[198])^(a[50] & b[199])^(a[49] & b[200])^(a[48] & b[201])^(a[47] & b[202])^(a[46] & b[203])^(a[45] & b[204])^(a[44] & b[205])^(a[43] & b[206])^(a[42] & b[207])^(a[41] & b[208])^(a[40] & b[209])^(a[39] & b[210])^(a[38] & b[211])^(a[37] & b[212])^(a[36] & b[213])^(a[35] & b[214])^(a[34] & b[215])^(a[33] & b[216])^(a[32] & b[217])^(a[31] & b[218])^(a[30] & b[219])^(a[29] & b[220])^(a[28] & b[221])^(a[27] & b[222])^(a[26] & b[223])^(a[25] & b[224])^(a[24] & b[225])^(a[23] & b[226])^(a[22] & b[227])^(a[21] & b[228])^(a[20] & b[229])^(a[19] & b[230])^(a[18] & b[231])^(a[17] & b[232]);
assign y[250] = (a[232] & b[18])^(a[231] & b[19])^(a[230] & b[20])^(a[229] & b[21])^(a[228] & b[22])^(a[227] & b[23])^(a[226] & b[24])^(a[225] & b[25])^(a[224] & b[26])^(a[223] & b[27])^(a[222] & b[28])^(a[221] & b[29])^(a[220] & b[30])^(a[219] & b[31])^(a[218] & b[32])^(a[217] & b[33])^(a[216] & b[34])^(a[215] & b[35])^(a[214] & b[36])^(a[213] & b[37])^(a[212] & b[38])^(a[211] & b[39])^(a[210] & b[40])^(a[209] & b[41])^(a[208] & b[42])^(a[207] & b[43])^(a[206] & b[44])^(a[205] & b[45])^(a[204] & b[46])^(a[203] & b[47])^(a[202] & b[48])^(a[201] & b[49])^(a[200] & b[50])^(a[199] & b[51])^(a[198] & b[52])^(a[197] & b[53])^(a[196] & b[54])^(a[195] & b[55])^(a[194] & b[56])^(a[193] & b[57])^(a[192] & b[58])^(a[191] & b[59])^(a[190] & b[60])^(a[189] & b[61])^(a[188] & b[62])^(a[187] & b[63])^(a[186] & b[64])^(a[185] & b[65])^(a[184] & b[66])^(a[183] & b[67])^(a[182] & b[68])^(a[181] & b[69])^(a[180] & b[70])^(a[179] & b[71])^(a[178] & b[72])^(a[177] & b[73])^(a[176] & b[74])^(a[175] & b[75])^(a[174] & b[76])^(a[173] & b[77])^(a[172] & b[78])^(a[171] & b[79])^(a[170] & b[80])^(a[169] & b[81])^(a[168] & b[82])^(a[167] & b[83])^(a[166] & b[84])^(a[165] & b[85])^(a[164] & b[86])^(a[163] & b[87])^(a[162] & b[88])^(a[161] & b[89])^(a[160] & b[90])^(a[159] & b[91])^(a[158] & b[92])^(a[157] & b[93])^(a[156] & b[94])^(a[155] & b[95])^(a[154] & b[96])^(a[153] & b[97])^(a[152] & b[98])^(a[151] & b[99])^(a[150] & b[100])^(a[149] & b[101])^(a[148] & b[102])^(a[147] & b[103])^(a[146] & b[104])^(a[145] & b[105])^(a[144] & b[106])^(a[143] & b[107])^(a[142] & b[108])^(a[141] & b[109])^(a[140] & b[110])^(a[139] & b[111])^(a[138] & b[112])^(a[137] & b[113])^(a[136] & b[114])^(a[135] & b[115])^(a[134] & b[116])^(a[133] & b[117])^(a[132] & b[118])^(a[131] & b[119])^(a[130] & b[120])^(a[129] & b[121])^(a[128] & b[122])^(a[127] & b[123])^(a[126] & b[124])^(a[125] & b[125])^(a[124] & b[126])^(a[123] & b[127])^(a[122] & b[128])^(a[121] & b[129])^(a[120] & b[130])^(a[119] & b[131])^(a[118] & b[132])^(a[117] & b[133])^(a[116] & b[134])^(a[115] & b[135])^(a[114] & b[136])^(a[113] & b[137])^(a[112] & b[138])^(a[111] & b[139])^(a[110] & b[140])^(a[109] & b[141])^(a[108] & b[142])^(a[107] & b[143])^(a[106] & b[144])^(a[105] & b[145])^(a[104] & b[146])^(a[103] & b[147])^(a[102] & b[148])^(a[101] & b[149])^(a[100] & b[150])^(a[99] & b[151])^(a[98] & b[152])^(a[97] & b[153])^(a[96] & b[154])^(a[95] & b[155])^(a[94] & b[156])^(a[93] & b[157])^(a[92] & b[158])^(a[91] & b[159])^(a[90] & b[160])^(a[89] & b[161])^(a[88] & b[162])^(a[87] & b[163])^(a[86] & b[164])^(a[85] & b[165])^(a[84] & b[166])^(a[83] & b[167])^(a[82] & b[168])^(a[81] & b[169])^(a[80] & b[170])^(a[79] & b[171])^(a[78] & b[172])^(a[77] & b[173])^(a[76] & b[174])^(a[75] & b[175])^(a[74] & b[176])^(a[73] & b[177])^(a[72] & b[178])^(a[71] & b[179])^(a[70] & b[180])^(a[69] & b[181])^(a[68] & b[182])^(a[67] & b[183])^(a[66] & b[184])^(a[65] & b[185])^(a[64] & b[186])^(a[63] & b[187])^(a[62] & b[188])^(a[61] & b[189])^(a[60] & b[190])^(a[59] & b[191])^(a[58] & b[192])^(a[57] & b[193])^(a[56] & b[194])^(a[55] & b[195])^(a[54] & b[196])^(a[53] & b[197])^(a[52] & b[198])^(a[51] & b[199])^(a[50] & b[200])^(a[49] & b[201])^(a[48] & b[202])^(a[47] & b[203])^(a[46] & b[204])^(a[45] & b[205])^(a[44] & b[206])^(a[43] & b[207])^(a[42] & b[208])^(a[41] & b[209])^(a[40] & b[210])^(a[39] & b[211])^(a[38] & b[212])^(a[37] & b[213])^(a[36] & b[214])^(a[35] & b[215])^(a[34] & b[216])^(a[33] & b[217])^(a[32] & b[218])^(a[31] & b[219])^(a[30] & b[220])^(a[29] & b[221])^(a[28] & b[222])^(a[27] & b[223])^(a[26] & b[224])^(a[25] & b[225])^(a[24] & b[226])^(a[23] & b[227])^(a[22] & b[228])^(a[21] & b[229])^(a[20] & b[230])^(a[19] & b[231])^(a[18] & b[232]);
assign y[251] = (a[232] & b[19])^(a[231] & b[20])^(a[230] & b[21])^(a[229] & b[22])^(a[228] & b[23])^(a[227] & b[24])^(a[226] & b[25])^(a[225] & b[26])^(a[224] & b[27])^(a[223] & b[28])^(a[222] & b[29])^(a[221] & b[30])^(a[220] & b[31])^(a[219] & b[32])^(a[218] & b[33])^(a[217] & b[34])^(a[216] & b[35])^(a[215] & b[36])^(a[214] & b[37])^(a[213] & b[38])^(a[212] & b[39])^(a[211] & b[40])^(a[210] & b[41])^(a[209] & b[42])^(a[208] & b[43])^(a[207] & b[44])^(a[206] & b[45])^(a[205] & b[46])^(a[204] & b[47])^(a[203] & b[48])^(a[202] & b[49])^(a[201] & b[50])^(a[200] & b[51])^(a[199] & b[52])^(a[198] & b[53])^(a[197] & b[54])^(a[196] & b[55])^(a[195] & b[56])^(a[194] & b[57])^(a[193] & b[58])^(a[192] & b[59])^(a[191] & b[60])^(a[190] & b[61])^(a[189] & b[62])^(a[188] & b[63])^(a[187] & b[64])^(a[186] & b[65])^(a[185] & b[66])^(a[184] & b[67])^(a[183] & b[68])^(a[182] & b[69])^(a[181] & b[70])^(a[180] & b[71])^(a[179] & b[72])^(a[178] & b[73])^(a[177] & b[74])^(a[176] & b[75])^(a[175] & b[76])^(a[174] & b[77])^(a[173] & b[78])^(a[172] & b[79])^(a[171] & b[80])^(a[170] & b[81])^(a[169] & b[82])^(a[168] & b[83])^(a[167] & b[84])^(a[166] & b[85])^(a[165] & b[86])^(a[164] & b[87])^(a[163] & b[88])^(a[162] & b[89])^(a[161] & b[90])^(a[160] & b[91])^(a[159] & b[92])^(a[158] & b[93])^(a[157] & b[94])^(a[156] & b[95])^(a[155] & b[96])^(a[154] & b[97])^(a[153] & b[98])^(a[152] & b[99])^(a[151] & b[100])^(a[150] & b[101])^(a[149] & b[102])^(a[148] & b[103])^(a[147] & b[104])^(a[146] & b[105])^(a[145] & b[106])^(a[144] & b[107])^(a[143] & b[108])^(a[142] & b[109])^(a[141] & b[110])^(a[140] & b[111])^(a[139] & b[112])^(a[138] & b[113])^(a[137] & b[114])^(a[136] & b[115])^(a[135] & b[116])^(a[134] & b[117])^(a[133] & b[118])^(a[132] & b[119])^(a[131] & b[120])^(a[130] & b[121])^(a[129] & b[122])^(a[128] & b[123])^(a[127] & b[124])^(a[126] & b[125])^(a[125] & b[126])^(a[124] & b[127])^(a[123] & b[128])^(a[122] & b[129])^(a[121] & b[130])^(a[120] & b[131])^(a[119] & b[132])^(a[118] & b[133])^(a[117] & b[134])^(a[116] & b[135])^(a[115] & b[136])^(a[114] & b[137])^(a[113] & b[138])^(a[112] & b[139])^(a[111] & b[140])^(a[110] & b[141])^(a[109] & b[142])^(a[108] & b[143])^(a[107] & b[144])^(a[106] & b[145])^(a[105] & b[146])^(a[104] & b[147])^(a[103] & b[148])^(a[102] & b[149])^(a[101] & b[150])^(a[100] & b[151])^(a[99] & b[152])^(a[98] & b[153])^(a[97] & b[154])^(a[96] & b[155])^(a[95] & b[156])^(a[94] & b[157])^(a[93] & b[158])^(a[92] & b[159])^(a[91] & b[160])^(a[90] & b[161])^(a[89] & b[162])^(a[88] & b[163])^(a[87] & b[164])^(a[86] & b[165])^(a[85] & b[166])^(a[84] & b[167])^(a[83] & b[168])^(a[82] & b[169])^(a[81] & b[170])^(a[80] & b[171])^(a[79] & b[172])^(a[78] & b[173])^(a[77] & b[174])^(a[76] & b[175])^(a[75] & b[176])^(a[74] & b[177])^(a[73] & b[178])^(a[72] & b[179])^(a[71] & b[180])^(a[70] & b[181])^(a[69] & b[182])^(a[68] & b[183])^(a[67] & b[184])^(a[66] & b[185])^(a[65] & b[186])^(a[64] & b[187])^(a[63] & b[188])^(a[62] & b[189])^(a[61] & b[190])^(a[60] & b[191])^(a[59] & b[192])^(a[58] & b[193])^(a[57] & b[194])^(a[56] & b[195])^(a[55] & b[196])^(a[54] & b[197])^(a[53] & b[198])^(a[52] & b[199])^(a[51] & b[200])^(a[50] & b[201])^(a[49] & b[202])^(a[48] & b[203])^(a[47] & b[204])^(a[46] & b[205])^(a[45] & b[206])^(a[44] & b[207])^(a[43] & b[208])^(a[42] & b[209])^(a[41] & b[210])^(a[40] & b[211])^(a[39] & b[212])^(a[38] & b[213])^(a[37] & b[214])^(a[36] & b[215])^(a[35] & b[216])^(a[34] & b[217])^(a[33] & b[218])^(a[32] & b[219])^(a[31] & b[220])^(a[30] & b[221])^(a[29] & b[222])^(a[28] & b[223])^(a[27] & b[224])^(a[26] & b[225])^(a[25] & b[226])^(a[24] & b[227])^(a[23] & b[228])^(a[22] & b[229])^(a[21] & b[230])^(a[20] & b[231])^(a[19] & b[232]);
assign y[252] = (a[232] & b[20])^(a[231] & b[21])^(a[230] & b[22])^(a[229] & b[23])^(a[228] & b[24])^(a[227] & b[25])^(a[226] & b[26])^(a[225] & b[27])^(a[224] & b[28])^(a[223] & b[29])^(a[222] & b[30])^(a[221] & b[31])^(a[220] & b[32])^(a[219] & b[33])^(a[218] & b[34])^(a[217] & b[35])^(a[216] & b[36])^(a[215] & b[37])^(a[214] & b[38])^(a[213] & b[39])^(a[212] & b[40])^(a[211] & b[41])^(a[210] & b[42])^(a[209] & b[43])^(a[208] & b[44])^(a[207] & b[45])^(a[206] & b[46])^(a[205] & b[47])^(a[204] & b[48])^(a[203] & b[49])^(a[202] & b[50])^(a[201] & b[51])^(a[200] & b[52])^(a[199] & b[53])^(a[198] & b[54])^(a[197] & b[55])^(a[196] & b[56])^(a[195] & b[57])^(a[194] & b[58])^(a[193] & b[59])^(a[192] & b[60])^(a[191] & b[61])^(a[190] & b[62])^(a[189] & b[63])^(a[188] & b[64])^(a[187] & b[65])^(a[186] & b[66])^(a[185] & b[67])^(a[184] & b[68])^(a[183] & b[69])^(a[182] & b[70])^(a[181] & b[71])^(a[180] & b[72])^(a[179] & b[73])^(a[178] & b[74])^(a[177] & b[75])^(a[176] & b[76])^(a[175] & b[77])^(a[174] & b[78])^(a[173] & b[79])^(a[172] & b[80])^(a[171] & b[81])^(a[170] & b[82])^(a[169] & b[83])^(a[168] & b[84])^(a[167] & b[85])^(a[166] & b[86])^(a[165] & b[87])^(a[164] & b[88])^(a[163] & b[89])^(a[162] & b[90])^(a[161] & b[91])^(a[160] & b[92])^(a[159] & b[93])^(a[158] & b[94])^(a[157] & b[95])^(a[156] & b[96])^(a[155] & b[97])^(a[154] & b[98])^(a[153] & b[99])^(a[152] & b[100])^(a[151] & b[101])^(a[150] & b[102])^(a[149] & b[103])^(a[148] & b[104])^(a[147] & b[105])^(a[146] & b[106])^(a[145] & b[107])^(a[144] & b[108])^(a[143] & b[109])^(a[142] & b[110])^(a[141] & b[111])^(a[140] & b[112])^(a[139] & b[113])^(a[138] & b[114])^(a[137] & b[115])^(a[136] & b[116])^(a[135] & b[117])^(a[134] & b[118])^(a[133] & b[119])^(a[132] & b[120])^(a[131] & b[121])^(a[130] & b[122])^(a[129] & b[123])^(a[128] & b[124])^(a[127] & b[125])^(a[126] & b[126])^(a[125] & b[127])^(a[124] & b[128])^(a[123] & b[129])^(a[122] & b[130])^(a[121] & b[131])^(a[120] & b[132])^(a[119] & b[133])^(a[118] & b[134])^(a[117] & b[135])^(a[116] & b[136])^(a[115] & b[137])^(a[114] & b[138])^(a[113] & b[139])^(a[112] & b[140])^(a[111] & b[141])^(a[110] & b[142])^(a[109] & b[143])^(a[108] & b[144])^(a[107] & b[145])^(a[106] & b[146])^(a[105] & b[147])^(a[104] & b[148])^(a[103] & b[149])^(a[102] & b[150])^(a[101] & b[151])^(a[100] & b[152])^(a[99] & b[153])^(a[98] & b[154])^(a[97] & b[155])^(a[96] & b[156])^(a[95] & b[157])^(a[94] & b[158])^(a[93] & b[159])^(a[92] & b[160])^(a[91] & b[161])^(a[90] & b[162])^(a[89] & b[163])^(a[88] & b[164])^(a[87] & b[165])^(a[86] & b[166])^(a[85] & b[167])^(a[84] & b[168])^(a[83] & b[169])^(a[82] & b[170])^(a[81] & b[171])^(a[80] & b[172])^(a[79] & b[173])^(a[78] & b[174])^(a[77] & b[175])^(a[76] & b[176])^(a[75] & b[177])^(a[74] & b[178])^(a[73] & b[179])^(a[72] & b[180])^(a[71] & b[181])^(a[70] & b[182])^(a[69] & b[183])^(a[68] & b[184])^(a[67] & b[185])^(a[66] & b[186])^(a[65] & b[187])^(a[64] & b[188])^(a[63] & b[189])^(a[62] & b[190])^(a[61] & b[191])^(a[60] & b[192])^(a[59] & b[193])^(a[58] & b[194])^(a[57] & b[195])^(a[56] & b[196])^(a[55] & b[197])^(a[54] & b[198])^(a[53] & b[199])^(a[52] & b[200])^(a[51] & b[201])^(a[50] & b[202])^(a[49] & b[203])^(a[48] & b[204])^(a[47] & b[205])^(a[46] & b[206])^(a[45] & b[207])^(a[44] & b[208])^(a[43] & b[209])^(a[42] & b[210])^(a[41] & b[211])^(a[40] & b[212])^(a[39] & b[213])^(a[38] & b[214])^(a[37] & b[215])^(a[36] & b[216])^(a[35] & b[217])^(a[34] & b[218])^(a[33] & b[219])^(a[32] & b[220])^(a[31] & b[221])^(a[30] & b[222])^(a[29] & b[223])^(a[28] & b[224])^(a[27] & b[225])^(a[26] & b[226])^(a[25] & b[227])^(a[24] & b[228])^(a[23] & b[229])^(a[22] & b[230])^(a[21] & b[231])^(a[20] & b[232]);
assign y[253] = (a[232] & b[21])^(a[231] & b[22])^(a[230] & b[23])^(a[229] & b[24])^(a[228] & b[25])^(a[227] & b[26])^(a[226] & b[27])^(a[225] & b[28])^(a[224] & b[29])^(a[223] & b[30])^(a[222] & b[31])^(a[221] & b[32])^(a[220] & b[33])^(a[219] & b[34])^(a[218] & b[35])^(a[217] & b[36])^(a[216] & b[37])^(a[215] & b[38])^(a[214] & b[39])^(a[213] & b[40])^(a[212] & b[41])^(a[211] & b[42])^(a[210] & b[43])^(a[209] & b[44])^(a[208] & b[45])^(a[207] & b[46])^(a[206] & b[47])^(a[205] & b[48])^(a[204] & b[49])^(a[203] & b[50])^(a[202] & b[51])^(a[201] & b[52])^(a[200] & b[53])^(a[199] & b[54])^(a[198] & b[55])^(a[197] & b[56])^(a[196] & b[57])^(a[195] & b[58])^(a[194] & b[59])^(a[193] & b[60])^(a[192] & b[61])^(a[191] & b[62])^(a[190] & b[63])^(a[189] & b[64])^(a[188] & b[65])^(a[187] & b[66])^(a[186] & b[67])^(a[185] & b[68])^(a[184] & b[69])^(a[183] & b[70])^(a[182] & b[71])^(a[181] & b[72])^(a[180] & b[73])^(a[179] & b[74])^(a[178] & b[75])^(a[177] & b[76])^(a[176] & b[77])^(a[175] & b[78])^(a[174] & b[79])^(a[173] & b[80])^(a[172] & b[81])^(a[171] & b[82])^(a[170] & b[83])^(a[169] & b[84])^(a[168] & b[85])^(a[167] & b[86])^(a[166] & b[87])^(a[165] & b[88])^(a[164] & b[89])^(a[163] & b[90])^(a[162] & b[91])^(a[161] & b[92])^(a[160] & b[93])^(a[159] & b[94])^(a[158] & b[95])^(a[157] & b[96])^(a[156] & b[97])^(a[155] & b[98])^(a[154] & b[99])^(a[153] & b[100])^(a[152] & b[101])^(a[151] & b[102])^(a[150] & b[103])^(a[149] & b[104])^(a[148] & b[105])^(a[147] & b[106])^(a[146] & b[107])^(a[145] & b[108])^(a[144] & b[109])^(a[143] & b[110])^(a[142] & b[111])^(a[141] & b[112])^(a[140] & b[113])^(a[139] & b[114])^(a[138] & b[115])^(a[137] & b[116])^(a[136] & b[117])^(a[135] & b[118])^(a[134] & b[119])^(a[133] & b[120])^(a[132] & b[121])^(a[131] & b[122])^(a[130] & b[123])^(a[129] & b[124])^(a[128] & b[125])^(a[127] & b[126])^(a[126] & b[127])^(a[125] & b[128])^(a[124] & b[129])^(a[123] & b[130])^(a[122] & b[131])^(a[121] & b[132])^(a[120] & b[133])^(a[119] & b[134])^(a[118] & b[135])^(a[117] & b[136])^(a[116] & b[137])^(a[115] & b[138])^(a[114] & b[139])^(a[113] & b[140])^(a[112] & b[141])^(a[111] & b[142])^(a[110] & b[143])^(a[109] & b[144])^(a[108] & b[145])^(a[107] & b[146])^(a[106] & b[147])^(a[105] & b[148])^(a[104] & b[149])^(a[103] & b[150])^(a[102] & b[151])^(a[101] & b[152])^(a[100] & b[153])^(a[99] & b[154])^(a[98] & b[155])^(a[97] & b[156])^(a[96] & b[157])^(a[95] & b[158])^(a[94] & b[159])^(a[93] & b[160])^(a[92] & b[161])^(a[91] & b[162])^(a[90] & b[163])^(a[89] & b[164])^(a[88] & b[165])^(a[87] & b[166])^(a[86] & b[167])^(a[85] & b[168])^(a[84] & b[169])^(a[83] & b[170])^(a[82] & b[171])^(a[81] & b[172])^(a[80] & b[173])^(a[79] & b[174])^(a[78] & b[175])^(a[77] & b[176])^(a[76] & b[177])^(a[75] & b[178])^(a[74] & b[179])^(a[73] & b[180])^(a[72] & b[181])^(a[71] & b[182])^(a[70] & b[183])^(a[69] & b[184])^(a[68] & b[185])^(a[67] & b[186])^(a[66] & b[187])^(a[65] & b[188])^(a[64] & b[189])^(a[63] & b[190])^(a[62] & b[191])^(a[61] & b[192])^(a[60] & b[193])^(a[59] & b[194])^(a[58] & b[195])^(a[57] & b[196])^(a[56] & b[197])^(a[55] & b[198])^(a[54] & b[199])^(a[53] & b[200])^(a[52] & b[201])^(a[51] & b[202])^(a[50] & b[203])^(a[49] & b[204])^(a[48] & b[205])^(a[47] & b[206])^(a[46] & b[207])^(a[45] & b[208])^(a[44] & b[209])^(a[43] & b[210])^(a[42] & b[211])^(a[41] & b[212])^(a[40] & b[213])^(a[39] & b[214])^(a[38] & b[215])^(a[37] & b[216])^(a[36] & b[217])^(a[35] & b[218])^(a[34] & b[219])^(a[33] & b[220])^(a[32] & b[221])^(a[31] & b[222])^(a[30] & b[223])^(a[29] & b[224])^(a[28] & b[225])^(a[27] & b[226])^(a[26] & b[227])^(a[25] & b[228])^(a[24] & b[229])^(a[23] & b[230])^(a[22] & b[231])^(a[21] & b[232]);
assign y[254] = (a[232] & b[22])^(a[231] & b[23])^(a[230] & b[24])^(a[229] & b[25])^(a[228] & b[26])^(a[227] & b[27])^(a[226] & b[28])^(a[225] & b[29])^(a[224] & b[30])^(a[223] & b[31])^(a[222] & b[32])^(a[221] & b[33])^(a[220] & b[34])^(a[219] & b[35])^(a[218] & b[36])^(a[217] & b[37])^(a[216] & b[38])^(a[215] & b[39])^(a[214] & b[40])^(a[213] & b[41])^(a[212] & b[42])^(a[211] & b[43])^(a[210] & b[44])^(a[209] & b[45])^(a[208] & b[46])^(a[207] & b[47])^(a[206] & b[48])^(a[205] & b[49])^(a[204] & b[50])^(a[203] & b[51])^(a[202] & b[52])^(a[201] & b[53])^(a[200] & b[54])^(a[199] & b[55])^(a[198] & b[56])^(a[197] & b[57])^(a[196] & b[58])^(a[195] & b[59])^(a[194] & b[60])^(a[193] & b[61])^(a[192] & b[62])^(a[191] & b[63])^(a[190] & b[64])^(a[189] & b[65])^(a[188] & b[66])^(a[187] & b[67])^(a[186] & b[68])^(a[185] & b[69])^(a[184] & b[70])^(a[183] & b[71])^(a[182] & b[72])^(a[181] & b[73])^(a[180] & b[74])^(a[179] & b[75])^(a[178] & b[76])^(a[177] & b[77])^(a[176] & b[78])^(a[175] & b[79])^(a[174] & b[80])^(a[173] & b[81])^(a[172] & b[82])^(a[171] & b[83])^(a[170] & b[84])^(a[169] & b[85])^(a[168] & b[86])^(a[167] & b[87])^(a[166] & b[88])^(a[165] & b[89])^(a[164] & b[90])^(a[163] & b[91])^(a[162] & b[92])^(a[161] & b[93])^(a[160] & b[94])^(a[159] & b[95])^(a[158] & b[96])^(a[157] & b[97])^(a[156] & b[98])^(a[155] & b[99])^(a[154] & b[100])^(a[153] & b[101])^(a[152] & b[102])^(a[151] & b[103])^(a[150] & b[104])^(a[149] & b[105])^(a[148] & b[106])^(a[147] & b[107])^(a[146] & b[108])^(a[145] & b[109])^(a[144] & b[110])^(a[143] & b[111])^(a[142] & b[112])^(a[141] & b[113])^(a[140] & b[114])^(a[139] & b[115])^(a[138] & b[116])^(a[137] & b[117])^(a[136] & b[118])^(a[135] & b[119])^(a[134] & b[120])^(a[133] & b[121])^(a[132] & b[122])^(a[131] & b[123])^(a[130] & b[124])^(a[129] & b[125])^(a[128] & b[126])^(a[127] & b[127])^(a[126] & b[128])^(a[125] & b[129])^(a[124] & b[130])^(a[123] & b[131])^(a[122] & b[132])^(a[121] & b[133])^(a[120] & b[134])^(a[119] & b[135])^(a[118] & b[136])^(a[117] & b[137])^(a[116] & b[138])^(a[115] & b[139])^(a[114] & b[140])^(a[113] & b[141])^(a[112] & b[142])^(a[111] & b[143])^(a[110] & b[144])^(a[109] & b[145])^(a[108] & b[146])^(a[107] & b[147])^(a[106] & b[148])^(a[105] & b[149])^(a[104] & b[150])^(a[103] & b[151])^(a[102] & b[152])^(a[101] & b[153])^(a[100] & b[154])^(a[99] & b[155])^(a[98] & b[156])^(a[97] & b[157])^(a[96] & b[158])^(a[95] & b[159])^(a[94] & b[160])^(a[93] & b[161])^(a[92] & b[162])^(a[91] & b[163])^(a[90] & b[164])^(a[89] & b[165])^(a[88] & b[166])^(a[87] & b[167])^(a[86] & b[168])^(a[85] & b[169])^(a[84] & b[170])^(a[83] & b[171])^(a[82] & b[172])^(a[81] & b[173])^(a[80] & b[174])^(a[79] & b[175])^(a[78] & b[176])^(a[77] & b[177])^(a[76] & b[178])^(a[75] & b[179])^(a[74] & b[180])^(a[73] & b[181])^(a[72] & b[182])^(a[71] & b[183])^(a[70] & b[184])^(a[69] & b[185])^(a[68] & b[186])^(a[67] & b[187])^(a[66] & b[188])^(a[65] & b[189])^(a[64] & b[190])^(a[63] & b[191])^(a[62] & b[192])^(a[61] & b[193])^(a[60] & b[194])^(a[59] & b[195])^(a[58] & b[196])^(a[57] & b[197])^(a[56] & b[198])^(a[55] & b[199])^(a[54] & b[200])^(a[53] & b[201])^(a[52] & b[202])^(a[51] & b[203])^(a[50] & b[204])^(a[49] & b[205])^(a[48] & b[206])^(a[47] & b[207])^(a[46] & b[208])^(a[45] & b[209])^(a[44] & b[210])^(a[43] & b[211])^(a[42] & b[212])^(a[41] & b[213])^(a[40] & b[214])^(a[39] & b[215])^(a[38] & b[216])^(a[37] & b[217])^(a[36] & b[218])^(a[35] & b[219])^(a[34] & b[220])^(a[33] & b[221])^(a[32] & b[222])^(a[31] & b[223])^(a[30] & b[224])^(a[29] & b[225])^(a[28] & b[226])^(a[27] & b[227])^(a[26] & b[228])^(a[25] & b[229])^(a[24] & b[230])^(a[23] & b[231])^(a[22] & b[232]);
assign y[255] = (a[232] & b[23])^(a[231] & b[24])^(a[230] & b[25])^(a[229] & b[26])^(a[228] & b[27])^(a[227] & b[28])^(a[226] & b[29])^(a[225] & b[30])^(a[224] & b[31])^(a[223] & b[32])^(a[222] & b[33])^(a[221] & b[34])^(a[220] & b[35])^(a[219] & b[36])^(a[218] & b[37])^(a[217] & b[38])^(a[216] & b[39])^(a[215] & b[40])^(a[214] & b[41])^(a[213] & b[42])^(a[212] & b[43])^(a[211] & b[44])^(a[210] & b[45])^(a[209] & b[46])^(a[208] & b[47])^(a[207] & b[48])^(a[206] & b[49])^(a[205] & b[50])^(a[204] & b[51])^(a[203] & b[52])^(a[202] & b[53])^(a[201] & b[54])^(a[200] & b[55])^(a[199] & b[56])^(a[198] & b[57])^(a[197] & b[58])^(a[196] & b[59])^(a[195] & b[60])^(a[194] & b[61])^(a[193] & b[62])^(a[192] & b[63])^(a[191] & b[64])^(a[190] & b[65])^(a[189] & b[66])^(a[188] & b[67])^(a[187] & b[68])^(a[186] & b[69])^(a[185] & b[70])^(a[184] & b[71])^(a[183] & b[72])^(a[182] & b[73])^(a[181] & b[74])^(a[180] & b[75])^(a[179] & b[76])^(a[178] & b[77])^(a[177] & b[78])^(a[176] & b[79])^(a[175] & b[80])^(a[174] & b[81])^(a[173] & b[82])^(a[172] & b[83])^(a[171] & b[84])^(a[170] & b[85])^(a[169] & b[86])^(a[168] & b[87])^(a[167] & b[88])^(a[166] & b[89])^(a[165] & b[90])^(a[164] & b[91])^(a[163] & b[92])^(a[162] & b[93])^(a[161] & b[94])^(a[160] & b[95])^(a[159] & b[96])^(a[158] & b[97])^(a[157] & b[98])^(a[156] & b[99])^(a[155] & b[100])^(a[154] & b[101])^(a[153] & b[102])^(a[152] & b[103])^(a[151] & b[104])^(a[150] & b[105])^(a[149] & b[106])^(a[148] & b[107])^(a[147] & b[108])^(a[146] & b[109])^(a[145] & b[110])^(a[144] & b[111])^(a[143] & b[112])^(a[142] & b[113])^(a[141] & b[114])^(a[140] & b[115])^(a[139] & b[116])^(a[138] & b[117])^(a[137] & b[118])^(a[136] & b[119])^(a[135] & b[120])^(a[134] & b[121])^(a[133] & b[122])^(a[132] & b[123])^(a[131] & b[124])^(a[130] & b[125])^(a[129] & b[126])^(a[128] & b[127])^(a[127] & b[128])^(a[126] & b[129])^(a[125] & b[130])^(a[124] & b[131])^(a[123] & b[132])^(a[122] & b[133])^(a[121] & b[134])^(a[120] & b[135])^(a[119] & b[136])^(a[118] & b[137])^(a[117] & b[138])^(a[116] & b[139])^(a[115] & b[140])^(a[114] & b[141])^(a[113] & b[142])^(a[112] & b[143])^(a[111] & b[144])^(a[110] & b[145])^(a[109] & b[146])^(a[108] & b[147])^(a[107] & b[148])^(a[106] & b[149])^(a[105] & b[150])^(a[104] & b[151])^(a[103] & b[152])^(a[102] & b[153])^(a[101] & b[154])^(a[100] & b[155])^(a[99] & b[156])^(a[98] & b[157])^(a[97] & b[158])^(a[96] & b[159])^(a[95] & b[160])^(a[94] & b[161])^(a[93] & b[162])^(a[92] & b[163])^(a[91] & b[164])^(a[90] & b[165])^(a[89] & b[166])^(a[88] & b[167])^(a[87] & b[168])^(a[86] & b[169])^(a[85] & b[170])^(a[84] & b[171])^(a[83] & b[172])^(a[82] & b[173])^(a[81] & b[174])^(a[80] & b[175])^(a[79] & b[176])^(a[78] & b[177])^(a[77] & b[178])^(a[76] & b[179])^(a[75] & b[180])^(a[74] & b[181])^(a[73] & b[182])^(a[72] & b[183])^(a[71] & b[184])^(a[70] & b[185])^(a[69] & b[186])^(a[68] & b[187])^(a[67] & b[188])^(a[66] & b[189])^(a[65] & b[190])^(a[64] & b[191])^(a[63] & b[192])^(a[62] & b[193])^(a[61] & b[194])^(a[60] & b[195])^(a[59] & b[196])^(a[58] & b[197])^(a[57] & b[198])^(a[56] & b[199])^(a[55] & b[200])^(a[54] & b[201])^(a[53] & b[202])^(a[52] & b[203])^(a[51] & b[204])^(a[50] & b[205])^(a[49] & b[206])^(a[48] & b[207])^(a[47] & b[208])^(a[46] & b[209])^(a[45] & b[210])^(a[44] & b[211])^(a[43] & b[212])^(a[42] & b[213])^(a[41] & b[214])^(a[40] & b[215])^(a[39] & b[216])^(a[38] & b[217])^(a[37] & b[218])^(a[36] & b[219])^(a[35] & b[220])^(a[34] & b[221])^(a[33] & b[222])^(a[32] & b[223])^(a[31] & b[224])^(a[30] & b[225])^(a[29] & b[226])^(a[28] & b[227])^(a[27] & b[228])^(a[26] & b[229])^(a[25] & b[230])^(a[24] & b[231])^(a[23] & b[232]);
assign y[256] = (a[232] & b[24])^(a[231] & b[25])^(a[230] & b[26])^(a[229] & b[27])^(a[228] & b[28])^(a[227] & b[29])^(a[226] & b[30])^(a[225] & b[31])^(a[224] & b[32])^(a[223] & b[33])^(a[222] & b[34])^(a[221] & b[35])^(a[220] & b[36])^(a[219] & b[37])^(a[218] & b[38])^(a[217] & b[39])^(a[216] & b[40])^(a[215] & b[41])^(a[214] & b[42])^(a[213] & b[43])^(a[212] & b[44])^(a[211] & b[45])^(a[210] & b[46])^(a[209] & b[47])^(a[208] & b[48])^(a[207] & b[49])^(a[206] & b[50])^(a[205] & b[51])^(a[204] & b[52])^(a[203] & b[53])^(a[202] & b[54])^(a[201] & b[55])^(a[200] & b[56])^(a[199] & b[57])^(a[198] & b[58])^(a[197] & b[59])^(a[196] & b[60])^(a[195] & b[61])^(a[194] & b[62])^(a[193] & b[63])^(a[192] & b[64])^(a[191] & b[65])^(a[190] & b[66])^(a[189] & b[67])^(a[188] & b[68])^(a[187] & b[69])^(a[186] & b[70])^(a[185] & b[71])^(a[184] & b[72])^(a[183] & b[73])^(a[182] & b[74])^(a[181] & b[75])^(a[180] & b[76])^(a[179] & b[77])^(a[178] & b[78])^(a[177] & b[79])^(a[176] & b[80])^(a[175] & b[81])^(a[174] & b[82])^(a[173] & b[83])^(a[172] & b[84])^(a[171] & b[85])^(a[170] & b[86])^(a[169] & b[87])^(a[168] & b[88])^(a[167] & b[89])^(a[166] & b[90])^(a[165] & b[91])^(a[164] & b[92])^(a[163] & b[93])^(a[162] & b[94])^(a[161] & b[95])^(a[160] & b[96])^(a[159] & b[97])^(a[158] & b[98])^(a[157] & b[99])^(a[156] & b[100])^(a[155] & b[101])^(a[154] & b[102])^(a[153] & b[103])^(a[152] & b[104])^(a[151] & b[105])^(a[150] & b[106])^(a[149] & b[107])^(a[148] & b[108])^(a[147] & b[109])^(a[146] & b[110])^(a[145] & b[111])^(a[144] & b[112])^(a[143] & b[113])^(a[142] & b[114])^(a[141] & b[115])^(a[140] & b[116])^(a[139] & b[117])^(a[138] & b[118])^(a[137] & b[119])^(a[136] & b[120])^(a[135] & b[121])^(a[134] & b[122])^(a[133] & b[123])^(a[132] & b[124])^(a[131] & b[125])^(a[130] & b[126])^(a[129] & b[127])^(a[128] & b[128])^(a[127] & b[129])^(a[126] & b[130])^(a[125] & b[131])^(a[124] & b[132])^(a[123] & b[133])^(a[122] & b[134])^(a[121] & b[135])^(a[120] & b[136])^(a[119] & b[137])^(a[118] & b[138])^(a[117] & b[139])^(a[116] & b[140])^(a[115] & b[141])^(a[114] & b[142])^(a[113] & b[143])^(a[112] & b[144])^(a[111] & b[145])^(a[110] & b[146])^(a[109] & b[147])^(a[108] & b[148])^(a[107] & b[149])^(a[106] & b[150])^(a[105] & b[151])^(a[104] & b[152])^(a[103] & b[153])^(a[102] & b[154])^(a[101] & b[155])^(a[100] & b[156])^(a[99] & b[157])^(a[98] & b[158])^(a[97] & b[159])^(a[96] & b[160])^(a[95] & b[161])^(a[94] & b[162])^(a[93] & b[163])^(a[92] & b[164])^(a[91] & b[165])^(a[90] & b[166])^(a[89] & b[167])^(a[88] & b[168])^(a[87] & b[169])^(a[86] & b[170])^(a[85] & b[171])^(a[84] & b[172])^(a[83] & b[173])^(a[82] & b[174])^(a[81] & b[175])^(a[80] & b[176])^(a[79] & b[177])^(a[78] & b[178])^(a[77] & b[179])^(a[76] & b[180])^(a[75] & b[181])^(a[74] & b[182])^(a[73] & b[183])^(a[72] & b[184])^(a[71] & b[185])^(a[70] & b[186])^(a[69] & b[187])^(a[68] & b[188])^(a[67] & b[189])^(a[66] & b[190])^(a[65] & b[191])^(a[64] & b[192])^(a[63] & b[193])^(a[62] & b[194])^(a[61] & b[195])^(a[60] & b[196])^(a[59] & b[197])^(a[58] & b[198])^(a[57] & b[199])^(a[56] & b[200])^(a[55] & b[201])^(a[54] & b[202])^(a[53] & b[203])^(a[52] & b[204])^(a[51] & b[205])^(a[50] & b[206])^(a[49] & b[207])^(a[48] & b[208])^(a[47] & b[209])^(a[46] & b[210])^(a[45] & b[211])^(a[44] & b[212])^(a[43] & b[213])^(a[42] & b[214])^(a[41] & b[215])^(a[40] & b[216])^(a[39] & b[217])^(a[38] & b[218])^(a[37] & b[219])^(a[36] & b[220])^(a[35] & b[221])^(a[34] & b[222])^(a[33] & b[223])^(a[32] & b[224])^(a[31] & b[225])^(a[30] & b[226])^(a[29] & b[227])^(a[28] & b[228])^(a[27] & b[229])^(a[26] & b[230])^(a[25] & b[231])^(a[24] & b[232]);
assign y[257] = (a[232] & b[25])^(a[231] & b[26])^(a[230] & b[27])^(a[229] & b[28])^(a[228] & b[29])^(a[227] & b[30])^(a[226] & b[31])^(a[225] & b[32])^(a[224] & b[33])^(a[223] & b[34])^(a[222] & b[35])^(a[221] & b[36])^(a[220] & b[37])^(a[219] & b[38])^(a[218] & b[39])^(a[217] & b[40])^(a[216] & b[41])^(a[215] & b[42])^(a[214] & b[43])^(a[213] & b[44])^(a[212] & b[45])^(a[211] & b[46])^(a[210] & b[47])^(a[209] & b[48])^(a[208] & b[49])^(a[207] & b[50])^(a[206] & b[51])^(a[205] & b[52])^(a[204] & b[53])^(a[203] & b[54])^(a[202] & b[55])^(a[201] & b[56])^(a[200] & b[57])^(a[199] & b[58])^(a[198] & b[59])^(a[197] & b[60])^(a[196] & b[61])^(a[195] & b[62])^(a[194] & b[63])^(a[193] & b[64])^(a[192] & b[65])^(a[191] & b[66])^(a[190] & b[67])^(a[189] & b[68])^(a[188] & b[69])^(a[187] & b[70])^(a[186] & b[71])^(a[185] & b[72])^(a[184] & b[73])^(a[183] & b[74])^(a[182] & b[75])^(a[181] & b[76])^(a[180] & b[77])^(a[179] & b[78])^(a[178] & b[79])^(a[177] & b[80])^(a[176] & b[81])^(a[175] & b[82])^(a[174] & b[83])^(a[173] & b[84])^(a[172] & b[85])^(a[171] & b[86])^(a[170] & b[87])^(a[169] & b[88])^(a[168] & b[89])^(a[167] & b[90])^(a[166] & b[91])^(a[165] & b[92])^(a[164] & b[93])^(a[163] & b[94])^(a[162] & b[95])^(a[161] & b[96])^(a[160] & b[97])^(a[159] & b[98])^(a[158] & b[99])^(a[157] & b[100])^(a[156] & b[101])^(a[155] & b[102])^(a[154] & b[103])^(a[153] & b[104])^(a[152] & b[105])^(a[151] & b[106])^(a[150] & b[107])^(a[149] & b[108])^(a[148] & b[109])^(a[147] & b[110])^(a[146] & b[111])^(a[145] & b[112])^(a[144] & b[113])^(a[143] & b[114])^(a[142] & b[115])^(a[141] & b[116])^(a[140] & b[117])^(a[139] & b[118])^(a[138] & b[119])^(a[137] & b[120])^(a[136] & b[121])^(a[135] & b[122])^(a[134] & b[123])^(a[133] & b[124])^(a[132] & b[125])^(a[131] & b[126])^(a[130] & b[127])^(a[129] & b[128])^(a[128] & b[129])^(a[127] & b[130])^(a[126] & b[131])^(a[125] & b[132])^(a[124] & b[133])^(a[123] & b[134])^(a[122] & b[135])^(a[121] & b[136])^(a[120] & b[137])^(a[119] & b[138])^(a[118] & b[139])^(a[117] & b[140])^(a[116] & b[141])^(a[115] & b[142])^(a[114] & b[143])^(a[113] & b[144])^(a[112] & b[145])^(a[111] & b[146])^(a[110] & b[147])^(a[109] & b[148])^(a[108] & b[149])^(a[107] & b[150])^(a[106] & b[151])^(a[105] & b[152])^(a[104] & b[153])^(a[103] & b[154])^(a[102] & b[155])^(a[101] & b[156])^(a[100] & b[157])^(a[99] & b[158])^(a[98] & b[159])^(a[97] & b[160])^(a[96] & b[161])^(a[95] & b[162])^(a[94] & b[163])^(a[93] & b[164])^(a[92] & b[165])^(a[91] & b[166])^(a[90] & b[167])^(a[89] & b[168])^(a[88] & b[169])^(a[87] & b[170])^(a[86] & b[171])^(a[85] & b[172])^(a[84] & b[173])^(a[83] & b[174])^(a[82] & b[175])^(a[81] & b[176])^(a[80] & b[177])^(a[79] & b[178])^(a[78] & b[179])^(a[77] & b[180])^(a[76] & b[181])^(a[75] & b[182])^(a[74] & b[183])^(a[73] & b[184])^(a[72] & b[185])^(a[71] & b[186])^(a[70] & b[187])^(a[69] & b[188])^(a[68] & b[189])^(a[67] & b[190])^(a[66] & b[191])^(a[65] & b[192])^(a[64] & b[193])^(a[63] & b[194])^(a[62] & b[195])^(a[61] & b[196])^(a[60] & b[197])^(a[59] & b[198])^(a[58] & b[199])^(a[57] & b[200])^(a[56] & b[201])^(a[55] & b[202])^(a[54] & b[203])^(a[53] & b[204])^(a[52] & b[205])^(a[51] & b[206])^(a[50] & b[207])^(a[49] & b[208])^(a[48] & b[209])^(a[47] & b[210])^(a[46] & b[211])^(a[45] & b[212])^(a[44] & b[213])^(a[43] & b[214])^(a[42] & b[215])^(a[41] & b[216])^(a[40] & b[217])^(a[39] & b[218])^(a[38] & b[219])^(a[37] & b[220])^(a[36] & b[221])^(a[35] & b[222])^(a[34] & b[223])^(a[33] & b[224])^(a[32] & b[225])^(a[31] & b[226])^(a[30] & b[227])^(a[29] & b[228])^(a[28] & b[229])^(a[27] & b[230])^(a[26] & b[231])^(a[25] & b[232]);
assign y[258] = (a[232] & b[26])^(a[231] & b[27])^(a[230] & b[28])^(a[229] & b[29])^(a[228] & b[30])^(a[227] & b[31])^(a[226] & b[32])^(a[225] & b[33])^(a[224] & b[34])^(a[223] & b[35])^(a[222] & b[36])^(a[221] & b[37])^(a[220] & b[38])^(a[219] & b[39])^(a[218] & b[40])^(a[217] & b[41])^(a[216] & b[42])^(a[215] & b[43])^(a[214] & b[44])^(a[213] & b[45])^(a[212] & b[46])^(a[211] & b[47])^(a[210] & b[48])^(a[209] & b[49])^(a[208] & b[50])^(a[207] & b[51])^(a[206] & b[52])^(a[205] & b[53])^(a[204] & b[54])^(a[203] & b[55])^(a[202] & b[56])^(a[201] & b[57])^(a[200] & b[58])^(a[199] & b[59])^(a[198] & b[60])^(a[197] & b[61])^(a[196] & b[62])^(a[195] & b[63])^(a[194] & b[64])^(a[193] & b[65])^(a[192] & b[66])^(a[191] & b[67])^(a[190] & b[68])^(a[189] & b[69])^(a[188] & b[70])^(a[187] & b[71])^(a[186] & b[72])^(a[185] & b[73])^(a[184] & b[74])^(a[183] & b[75])^(a[182] & b[76])^(a[181] & b[77])^(a[180] & b[78])^(a[179] & b[79])^(a[178] & b[80])^(a[177] & b[81])^(a[176] & b[82])^(a[175] & b[83])^(a[174] & b[84])^(a[173] & b[85])^(a[172] & b[86])^(a[171] & b[87])^(a[170] & b[88])^(a[169] & b[89])^(a[168] & b[90])^(a[167] & b[91])^(a[166] & b[92])^(a[165] & b[93])^(a[164] & b[94])^(a[163] & b[95])^(a[162] & b[96])^(a[161] & b[97])^(a[160] & b[98])^(a[159] & b[99])^(a[158] & b[100])^(a[157] & b[101])^(a[156] & b[102])^(a[155] & b[103])^(a[154] & b[104])^(a[153] & b[105])^(a[152] & b[106])^(a[151] & b[107])^(a[150] & b[108])^(a[149] & b[109])^(a[148] & b[110])^(a[147] & b[111])^(a[146] & b[112])^(a[145] & b[113])^(a[144] & b[114])^(a[143] & b[115])^(a[142] & b[116])^(a[141] & b[117])^(a[140] & b[118])^(a[139] & b[119])^(a[138] & b[120])^(a[137] & b[121])^(a[136] & b[122])^(a[135] & b[123])^(a[134] & b[124])^(a[133] & b[125])^(a[132] & b[126])^(a[131] & b[127])^(a[130] & b[128])^(a[129] & b[129])^(a[128] & b[130])^(a[127] & b[131])^(a[126] & b[132])^(a[125] & b[133])^(a[124] & b[134])^(a[123] & b[135])^(a[122] & b[136])^(a[121] & b[137])^(a[120] & b[138])^(a[119] & b[139])^(a[118] & b[140])^(a[117] & b[141])^(a[116] & b[142])^(a[115] & b[143])^(a[114] & b[144])^(a[113] & b[145])^(a[112] & b[146])^(a[111] & b[147])^(a[110] & b[148])^(a[109] & b[149])^(a[108] & b[150])^(a[107] & b[151])^(a[106] & b[152])^(a[105] & b[153])^(a[104] & b[154])^(a[103] & b[155])^(a[102] & b[156])^(a[101] & b[157])^(a[100] & b[158])^(a[99] & b[159])^(a[98] & b[160])^(a[97] & b[161])^(a[96] & b[162])^(a[95] & b[163])^(a[94] & b[164])^(a[93] & b[165])^(a[92] & b[166])^(a[91] & b[167])^(a[90] & b[168])^(a[89] & b[169])^(a[88] & b[170])^(a[87] & b[171])^(a[86] & b[172])^(a[85] & b[173])^(a[84] & b[174])^(a[83] & b[175])^(a[82] & b[176])^(a[81] & b[177])^(a[80] & b[178])^(a[79] & b[179])^(a[78] & b[180])^(a[77] & b[181])^(a[76] & b[182])^(a[75] & b[183])^(a[74] & b[184])^(a[73] & b[185])^(a[72] & b[186])^(a[71] & b[187])^(a[70] & b[188])^(a[69] & b[189])^(a[68] & b[190])^(a[67] & b[191])^(a[66] & b[192])^(a[65] & b[193])^(a[64] & b[194])^(a[63] & b[195])^(a[62] & b[196])^(a[61] & b[197])^(a[60] & b[198])^(a[59] & b[199])^(a[58] & b[200])^(a[57] & b[201])^(a[56] & b[202])^(a[55] & b[203])^(a[54] & b[204])^(a[53] & b[205])^(a[52] & b[206])^(a[51] & b[207])^(a[50] & b[208])^(a[49] & b[209])^(a[48] & b[210])^(a[47] & b[211])^(a[46] & b[212])^(a[45] & b[213])^(a[44] & b[214])^(a[43] & b[215])^(a[42] & b[216])^(a[41] & b[217])^(a[40] & b[218])^(a[39] & b[219])^(a[38] & b[220])^(a[37] & b[221])^(a[36] & b[222])^(a[35] & b[223])^(a[34] & b[224])^(a[33] & b[225])^(a[32] & b[226])^(a[31] & b[227])^(a[30] & b[228])^(a[29] & b[229])^(a[28] & b[230])^(a[27] & b[231])^(a[26] & b[232]);
assign y[259] = (a[232] & b[27])^(a[231] & b[28])^(a[230] & b[29])^(a[229] & b[30])^(a[228] & b[31])^(a[227] & b[32])^(a[226] & b[33])^(a[225] & b[34])^(a[224] & b[35])^(a[223] & b[36])^(a[222] & b[37])^(a[221] & b[38])^(a[220] & b[39])^(a[219] & b[40])^(a[218] & b[41])^(a[217] & b[42])^(a[216] & b[43])^(a[215] & b[44])^(a[214] & b[45])^(a[213] & b[46])^(a[212] & b[47])^(a[211] & b[48])^(a[210] & b[49])^(a[209] & b[50])^(a[208] & b[51])^(a[207] & b[52])^(a[206] & b[53])^(a[205] & b[54])^(a[204] & b[55])^(a[203] & b[56])^(a[202] & b[57])^(a[201] & b[58])^(a[200] & b[59])^(a[199] & b[60])^(a[198] & b[61])^(a[197] & b[62])^(a[196] & b[63])^(a[195] & b[64])^(a[194] & b[65])^(a[193] & b[66])^(a[192] & b[67])^(a[191] & b[68])^(a[190] & b[69])^(a[189] & b[70])^(a[188] & b[71])^(a[187] & b[72])^(a[186] & b[73])^(a[185] & b[74])^(a[184] & b[75])^(a[183] & b[76])^(a[182] & b[77])^(a[181] & b[78])^(a[180] & b[79])^(a[179] & b[80])^(a[178] & b[81])^(a[177] & b[82])^(a[176] & b[83])^(a[175] & b[84])^(a[174] & b[85])^(a[173] & b[86])^(a[172] & b[87])^(a[171] & b[88])^(a[170] & b[89])^(a[169] & b[90])^(a[168] & b[91])^(a[167] & b[92])^(a[166] & b[93])^(a[165] & b[94])^(a[164] & b[95])^(a[163] & b[96])^(a[162] & b[97])^(a[161] & b[98])^(a[160] & b[99])^(a[159] & b[100])^(a[158] & b[101])^(a[157] & b[102])^(a[156] & b[103])^(a[155] & b[104])^(a[154] & b[105])^(a[153] & b[106])^(a[152] & b[107])^(a[151] & b[108])^(a[150] & b[109])^(a[149] & b[110])^(a[148] & b[111])^(a[147] & b[112])^(a[146] & b[113])^(a[145] & b[114])^(a[144] & b[115])^(a[143] & b[116])^(a[142] & b[117])^(a[141] & b[118])^(a[140] & b[119])^(a[139] & b[120])^(a[138] & b[121])^(a[137] & b[122])^(a[136] & b[123])^(a[135] & b[124])^(a[134] & b[125])^(a[133] & b[126])^(a[132] & b[127])^(a[131] & b[128])^(a[130] & b[129])^(a[129] & b[130])^(a[128] & b[131])^(a[127] & b[132])^(a[126] & b[133])^(a[125] & b[134])^(a[124] & b[135])^(a[123] & b[136])^(a[122] & b[137])^(a[121] & b[138])^(a[120] & b[139])^(a[119] & b[140])^(a[118] & b[141])^(a[117] & b[142])^(a[116] & b[143])^(a[115] & b[144])^(a[114] & b[145])^(a[113] & b[146])^(a[112] & b[147])^(a[111] & b[148])^(a[110] & b[149])^(a[109] & b[150])^(a[108] & b[151])^(a[107] & b[152])^(a[106] & b[153])^(a[105] & b[154])^(a[104] & b[155])^(a[103] & b[156])^(a[102] & b[157])^(a[101] & b[158])^(a[100] & b[159])^(a[99] & b[160])^(a[98] & b[161])^(a[97] & b[162])^(a[96] & b[163])^(a[95] & b[164])^(a[94] & b[165])^(a[93] & b[166])^(a[92] & b[167])^(a[91] & b[168])^(a[90] & b[169])^(a[89] & b[170])^(a[88] & b[171])^(a[87] & b[172])^(a[86] & b[173])^(a[85] & b[174])^(a[84] & b[175])^(a[83] & b[176])^(a[82] & b[177])^(a[81] & b[178])^(a[80] & b[179])^(a[79] & b[180])^(a[78] & b[181])^(a[77] & b[182])^(a[76] & b[183])^(a[75] & b[184])^(a[74] & b[185])^(a[73] & b[186])^(a[72] & b[187])^(a[71] & b[188])^(a[70] & b[189])^(a[69] & b[190])^(a[68] & b[191])^(a[67] & b[192])^(a[66] & b[193])^(a[65] & b[194])^(a[64] & b[195])^(a[63] & b[196])^(a[62] & b[197])^(a[61] & b[198])^(a[60] & b[199])^(a[59] & b[200])^(a[58] & b[201])^(a[57] & b[202])^(a[56] & b[203])^(a[55] & b[204])^(a[54] & b[205])^(a[53] & b[206])^(a[52] & b[207])^(a[51] & b[208])^(a[50] & b[209])^(a[49] & b[210])^(a[48] & b[211])^(a[47] & b[212])^(a[46] & b[213])^(a[45] & b[214])^(a[44] & b[215])^(a[43] & b[216])^(a[42] & b[217])^(a[41] & b[218])^(a[40] & b[219])^(a[39] & b[220])^(a[38] & b[221])^(a[37] & b[222])^(a[36] & b[223])^(a[35] & b[224])^(a[34] & b[225])^(a[33] & b[226])^(a[32] & b[227])^(a[31] & b[228])^(a[30] & b[229])^(a[29] & b[230])^(a[28] & b[231])^(a[27] & b[232]);
assign y[260] = (a[232] & b[28])^(a[231] & b[29])^(a[230] & b[30])^(a[229] & b[31])^(a[228] & b[32])^(a[227] & b[33])^(a[226] & b[34])^(a[225] & b[35])^(a[224] & b[36])^(a[223] & b[37])^(a[222] & b[38])^(a[221] & b[39])^(a[220] & b[40])^(a[219] & b[41])^(a[218] & b[42])^(a[217] & b[43])^(a[216] & b[44])^(a[215] & b[45])^(a[214] & b[46])^(a[213] & b[47])^(a[212] & b[48])^(a[211] & b[49])^(a[210] & b[50])^(a[209] & b[51])^(a[208] & b[52])^(a[207] & b[53])^(a[206] & b[54])^(a[205] & b[55])^(a[204] & b[56])^(a[203] & b[57])^(a[202] & b[58])^(a[201] & b[59])^(a[200] & b[60])^(a[199] & b[61])^(a[198] & b[62])^(a[197] & b[63])^(a[196] & b[64])^(a[195] & b[65])^(a[194] & b[66])^(a[193] & b[67])^(a[192] & b[68])^(a[191] & b[69])^(a[190] & b[70])^(a[189] & b[71])^(a[188] & b[72])^(a[187] & b[73])^(a[186] & b[74])^(a[185] & b[75])^(a[184] & b[76])^(a[183] & b[77])^(a[182] & b[78])^(a[181] & b[79])^(a[180] & b[80])^(a[179] & b[81])^(a[178] & b[82])^(a[177] & b[83])^(a[176] & b[84])^(a[175] & b[85])^(a[174] & b[86])^(a[173] & b[87])^(a[172] & b[88])^(a[171] & b[89])^(a[170] & b[90])^(a[169] & b[91])^(a[168] & b[92])^(a[167] & b[93])^(a[166] & b[94])^(a[165] & b[95])^(a[164] & b[96])^(a[163] & b[97])^(a[162] & b[98])^(a[161] & b[99])^(a[160] & b[100])^(a[159] & b[101])^(a[158] & b[102])^(a[157] & b[103])^(a[156] & b[104])^(a[155] & b[105])^(a[154] & b[106])^(a[153] & b[107])^(a[152] & b[108])^(a[151] & b[109])^(a[150] & b[110])^(a[149] & b[111])^(a[148] & b[112])^(a[147] & b[113])^(a[146] & b[114])^(a[145] & b[115])^(a[144] & b[116])^(a[143] & b[117])^(a[142] & b[118])^(a[141] & b[119])^(a[140] & b[120])^(a[139] & b[121])^(a[138] & b[122])^(a[137] & b[123])^(a[136] & b[124])^(a[135] & b[125])^(a[134] & b[126])^(a[133] & b[127])^(a[132] & b[128])^(a[131] & b[129])^(a[130] & b[130])^(a[129] & b[131])^(a[128] & b[132])^(a[127] & b[133])^(a[126] & b[134])^(a[125] & b[135])^(a[124] & b[136])^(a[123] & b[137])^(a[122] & b[138])^(a[121] & b[139])^(a[120] & b[140])^(a[119] & b[141])^(a[118] & b[142])^(a[117] & b[143])^(a[116] & b[144])^(a[115] & b[145])^(a[114] & b[146])^(a[113] & b[147])^(a[112] & b[148])^(a[111] & b[149])^(a[110] & b[150])^(a[109] & b[151])^(a[108] & b[152])^(a[107] & b[153])^(a[106] & b[154])^(a[105] & b[155])^(a[104] & b[156])^(a[103] & b[157])^(a[102] & b[158])^(a[101] & b[159])^(a[100] & b[160])^(a[99] & b[161])^(a[98] & b[162])^(a[97] & b[163])^(a[96] & b[164])^(a[95] & b[165])^(a[94] & b[166])^(a[93] & b[167])^(a[92] & b[168])^(a[91] & b[169])^(a[90] & b[170])^(a[89] & b[171])^(a[88] & b[172])^(a[87] & b[173])^(a[86] & b[174])^(a[85] & b[175])^(a[84] & b[176])^(a[83] & b[177])^(a[82] & b[178])^(a[81] & b[179])^(a[80] & b[180])^(a[79] & b[181])^(a[78] & b[182])^(a[77] & b[183])^(a[76] & b[184])^(a[75] & b[185])^(a[74] & b[186])^(a[73] & b[187])^(a[72] & b[188])^(a[71] & b[189])^(a[70] & b[190])^(a[69] & b[191])^(a[68] & b[192])^(a[67] & b[193])^(a[66] & b[194])^(a[65] & b[195])^(a[64] & b[196])^(a[63] & b[197])^(a[62] & b[198])^(a[61] & b[199])^(a[60] & b[200])^(a[59] & b[201])^(a[58] & b[202])^(a[57] & b[203])^(a[56] & b[204])^(a[55] & b[205])^(a[54] & b[206])^(a[53] & b[207])^(a[52] & b[208])^(a[51] & b[209])^(a[50] & b[210])^(a[49] & b[211])^(a[48] & b[212])^(a[47] & b[213])^(a[46] & b[214])^(a[45] & b[215])^(a[44] & b[216])^(a[43] & b[217])^(a[42] & b[218])^(a[41] & b[219])^(a[40] & b[220])^(a[39] & b[221])^(a[38] & b[222])^(a[37] & b[223])^(a[36] & b[224])^(a[35] & b[225])^(a[34] & b[226])^(a[33] & b[227])^(a[32] & b[228])^(a[31] & b[229])^(a[30] & b[230])^(a[29] & b[231])^(a[28] & b[232]);
assign y[261] = (a[232] & b[29])^(a[231] & b[30])^(a[230] & b[31])^(a[229] & b[32])^(a[228] & b[33])^(a[227] & b[34])^(a[226] & b[35])^(a[225] & b[36])^(a[224] & b[37])^(a[223] & b[38])^(a[222] & b[39])^(a[221] & b[40])^(a[220] & b[41])^(a[219] & b[42])^(a[218] & b[43])^(a[217] & b[44])^(a[216] & b[45])^(a[215] & b[46])^(a[214] & b[47])^(a[213] & b[48])^(a[212] & b[49])^(a[211] & b[50])^(a[210] & b[51])^(a[209] & b[52])^(a[208] & b[53])^(a[207] & b[54])^(a[206] & b[55])^(a[205] & b[56])^(a[204] & b[57])^(a[203] & b[58])^(a[202] & b[59])^(a[201] & b[60])^(a[200] & b[61])^(a[199] & b[62])^(a[198] & b[63])^(a[197] & b[64])^(a[196] & b[65])^(a[195] & b[66])^(a[194] & b[67])^(a[193] & b[68])^(a[192] & b[69])^(a[191] & b[70])^(a[190] & b[71])^(a[189] & b[72])^(a[188] & b[73])^(a[187] & b[74])^(a[186] & b[75])^(a[185] & b[76])^(a[184] & b[77])^(a[183] & b[78])^(a[182] & b[79])^(a[181] & b[80])^(a[180] & b[81])^(a[179] & b[82])^(a[178] & b[83])^(a[177] & b[84])^(a[176] & b[85])^(a[175] & b[86])^(a[174] & b[87])^(a[173] & b[88])^(a[172] & b[89])^(a[171] & b[90])^(a[170] & b[91])^(a[169] & b[92])^(a[168] & b[93])^(a[167] & b[94])^(a[166] & b[95])^(a[165] & b[96])^(a[164] & b[97])^(a[163] & b[98])^(a[162] & b[99])^(a[161] & b[100])^(a[160] & b[101])^(a[159] & b[102])^(a[158] & b[103])^(a[157] & b[104])^(a[156] & b[105])^(a[155] & b[106])^(a[154] & b[107])^(a[153] & b[108])^(a[152] & b[109])^(a[151] & b[110])^(a[150] & b[111])^(a[149] & b[112])^(a[148] & b[113])^(a[147] & b[114])^(a[146] & b[115])^(a[145] & b[116])^(a[144] & b[117])^(a[143] & b[118])^(a[142] & b[119])^(a[141] & b[120])^(a[140] & b[121])^(a[139] & b[122])^(a[138] & b[123])^(a[137] & b[124])^(a[136] & b[125])^(a[135] & b[126])^(a[134] & b[127])^(a[133] & b[128])^(a[132] & b[129])^(a[131] & b[130])^(a[130] & b[131])^(a[129] & b[132])^(a[128] & b[133])^(a[127] & b[134])^(a[126] & b[135])^(a[125] & b[136])^(a[124] & b[137])^(a[123] & b[138])^(a[122] & b[139])^(a[121] & b[140])^(a[120] & b[141])^(a[119] & b[142])^(a[118] & b[143])^(a[117] & b[144])^(a[116] & b[145])^(a[115] & b[146])^(a[114] & b[147])^(a[113] & b[148])^(a[112] & b[149])^(a[111] & b[150])^(a[110] & b[151])^(a[109] & b[152])^(a[108] & b[153])^(a[107] & b[154])^(a[106] & b[155])^(a[105] & b[156])^(a[104] & b[157])^(a[103] & b[158])^(a[102] & b[159])^(a[101] & b[160])^(a[100] & b[161])^(a[99] & b[162])^(a[98] & b[163])^(a[97] & b[164])^(a[96] & b[165])^(a[95] & b[166])^(a[94] & b[167])^(a[93] & b[168])^(a[92] & b[169])^(a[91] & b[170])^(a[90] & b[171])^(a[89] & b[172])^(a[88] & b[173])^(a[87] & b[174])^(a[86] & b[175])^(a[85] & b[176])^(a[84] & b[177])^(a[83] & b[178])^(a[82] & b[179])^(a[81] & b[180])^(a[80] & b[181])^(a[79] & b[182])^(a[78] & b[183])^(a[77] & b[184])^(a[76] & b[185])^(a[75] & b[186])^(a[74] & b[187])^(a[73] & b[188])^(a[72] & b[189])^(a[71] & b[190])^(a[70] & b[191])^(a[69] & b[192])^(a[68] & b[193])^(a[67] & b[194])^(a[66] & b[195])^(a[65] & b[196])^(a[64] & b[197])^(a[63] & b[198])^(a[62] & b[199])^(a[61] & b[200])^(a[60] & b[201])^(a[59] & b[202])^(a[58] & b[203])^(a[57] & b[204])^(a[56] & b[205])^(a[55] & b[206])^(a[54] & b[207])^(a[53] & b[208])^(a[52] & b[209])^(a[51] & b[210])^(a[50] & b[211])^(a[49] & b[212])^(a[48] & b[213])^(a[47] & b[214])^(a[46] & b[215])^(a[45] & b[216])^(a[44] & b[217])^(a[43] & b[218])^(a[42] & b[219])^(a[41] & b[220])^(a[40] & b[221])^(a[39] & b[222])^(a[38] & b[223])^(a[37] & b[224])^(a[36] & b[225])^(a[35] & b[226])^(a[34] & b[227])^(a[33] & b[228])^(a[32] & b[229])^(a[31] & b[230])^(a[30] & b[231])^(a[29] & b[232]);
assign y[262] = (a[232] & b[30])^(a[231] & b[31])^(a[230] & b[32])^(a[229] & b[33])^(a[228] & b[34])^(a[227] & b[35])^(a[226] & b[36])^(a[225] & b[37])^(a[224] & b[38])^(a[223] & b[39])^(a[222] & b[40])^(a[221] & b[41])^(a[220] & b[42])^(a[219] & b[43])^(a[218] & b[44])^(a[217] & b[45])^(a[216] & b[46])^(a[215] & b[47])^(a[214] & b[48])^(a[213] & b[49])^(a[212] & b[50])^(a[211] & b[51])^(a[210] & b[52])^(a[209] & b[53])^(a[208] & b[54])^(a[207] & b[55])^(a[206] & b[56])^(a[205] & b[57])^(a[204] & b[58])^(a[203] & b[59])^(a[202] & b[60])^(a[201] & b[61])^(a[200] & b[62])^(a[199] & b[63])^(a[198] & b[64])^(a[197] & b[65])^(a[196] & b[66])^(a[195] & b[67])^(a[194] & b[68])^(a[193] & b[69])^(a[192] & b[70])^(a[191] & b[71])^(a[190] & b[72])^(a[189] & b[73])^(a[188] & b[74])^(a[187] & b[75])^(a[186] & b[76])^(a[185] & b[77])^(a[184] & b[78])^(a[183] & b[79])^(a[182] & b[80])^(a[181] & b[81])^(a[180] & b[82])^(a[179] & b[83])^(a[178] & b[84])^(a[177] & b[85])^(a[176] & b[86])^(a[175] & b[87])^(a[174] & b[88])^(a[173] & b[89])^(a[172] & b[90])^(a[171] & b[91])^(a[170] & b[92])^(a[169] & b[93])^(a[168] & b[94])^(a[167] & b[95])^(a[166] & b[96])^(a[165] & b[97])^(a[164] & b[98])^(a[163] & b[99])^(a[162] & b[100])^(a[161] & b[101])^(a[160] & b[102])^(a[159] & b[103])^(a[158] & b[104])^(a[157] & b[105])^(a[156] & b[106])^(a[155] & b[107])^(a[154] & b[108])^(a[153] & b[109])^(a[152] & b[110])^(a[151] & b[111])^(a[150] & b[112])^(a[149] & b[113])^(a[148] & b[114])^(a[147] & b[115])^(a[146] & b[116])^(a[145] & b[117])^(a[144] & b[118])^(a[143] & b[119])^(a[142] & b[120])^(a[141] & b[121])^(a[140] & b[122])^(a[139] & b[123])^(a[138] & b[124])^(a[137] & b[125])^(a[136] & b[126])^(a[135] & b[127])^(a[134] & b[128])^(a[133] & b[129])^(a[132] & b[130])^(a[131] & b[131])^(a[130] & b[132])^(a[129] & b[133])^(a[128] & b[134])^(a[127] & b[135])^(a[126] & b[136])^(a[125] & b[137])^(a[124] & b[138])^(a[123] & b[139])^(a[122] & b[140])^(a[121] & b[141])^(a[120] & b[142])^(a[119] & b[143])^(a[118] & b[144])^(a[117] & b[145])^(a[116] & b[146])^(a[115] & b[147])^(a[114] & b[148])^(a[113] & b[149])^(a[112] & b[150])^(a[111] & b[151])^(a[110] & b[152])^(a[109] & b[153])^(a[108] & b[154])^(a[107] & b[155])^(a[106] & b[156])^(a[105] & b[157])^(a[104] & b[158])^(a[103] & b[159])^(a[102] & b[160])^(a[101] & b[161])^(a[100] & b[162])^(a[99] & b[163])^(a[98] & b[164])^(a[97] & b[165])^(a[96] & b[166])^(a[95] & b[167])^(a[94] & b[168])^(a[93] & b[169])^(a[92] & b[170])^(a[91] & b[171])^(a[90] & b[172])^(a[89] & b[173])^(a[88] & b[174])^(a[87] & b[175])^(a[86] & b[176])^(a[85] & b[177])^(a[84] & b[178])^(a[83] & b[179])^(a[82] & b[180])^(a[81] & b[181])^(a[80] & b[182])^(a[79] & b[183])^(a[78] & b[184])^(a[77] & b[185])^(a[76] & b[186])^(a[75] & b[187])^(a[74] & b[188])^(a[73] & b[189])^(a[72] & b[190])^(a[71] & b[191])^(a[70] & b[192])^(a[69] & b[193])^(a[68] & b[194])^(a[67] & b[195])^(a[66] & b[196])^(a[65] & b[197])^(a[64] & b[198])^(a[63] & b[199])^(a[62] & b[200])^(a[61] & b[201])^(a[60] & b[202])^(a[59] & b[203])^(a[58] & b[204])^(a[57] & b[205])^(a[56] & b[206])^(a[55] & b[207])^(a[54] & b[208])^(a[53] & b[209])^(a[52] & b[210])^(a[51] & b[211])^(a[50] & b[212])^(a[49] & b[213])^(a[48] & b[214])^(a[47] & b[215])^(a[46] & b[216])^(a[45] & b[217])^(a[44] & b[218])^(a[43] & b[219])^(a[42] & b[220])^(a[41] & b[221])^(a[40] & b[222])^(a[39] & b[223])^(a[38] & b[224])^(a[37] & b[225])^(a[36] & b[226])^(a[35] & b[227])^(a[34] & b[228])^(a[33] & b[229])^(a[32] & b[230])^(a[31] & b[231])^(a[30] & b[232]);
assign y[263] = (a[232] & b[31])^(a[231] & b[32])^(a[230] & b[33])^(a[229] & b[34])^(a[228] & b[35])^(a[227] & b[36])^(a[226] & b[37])^(a[225] & b[38])^(a[224] & b[39])^(a[223] & b[40])^(a[222] & b[41])^(a[221] & b[42])^(a[220] & b[43])^(a[219] & b[44])^(a[218] & b[45])^(a[217] & b[46])^(a[216] & b[47])^(a[215] & b[48])^(a[214] & b[49])^(a[213] & b[50])^(a[212] & b[51])^(a[211] & b[52])^(a[210] & b[53])^(a[209] & b[54])^(a[208] & b[55])^(a[207] & b[56])^(a[206] & b[57])^(a[205] & b[58])^(a[204] & b[59])^(a[203] & b[60])^(a[202] & b[61])^(a[201] & b[62])^(a[200] & b[63])^(a[199] & b[64])^(a[198] & b[65])^(a[197] & b[66])^(a[196] & b[67])^(a[195] & b[68])^(a[194] & b[69])^(a[193] & b[70])^(a[192] & b[71])^(a[191] & b[72])^(a[190] & b[73])^(a[189] & b[74])^(a[188] & b[75])^(a[187] & b[76])^(a[186] & b[77])^(a[185] & b[78])^(a[184] & b[79])^(a[183] & b[80])^(a[182] & b[81])^(a[181] & b[82])^(a[180] & b[83])^(a[179] & b[84])^(a[178] & b[85])^(a[177] & b[86])^(a[176] & b[87])^(a[175] & b[88])^(a[174] & b[89])^(a[173] & b[90])^(a[172] & b[91])^(a[171] & b[92])^(a[170] & b[93])^(a[169] & b[94])^(a[168] & b[95])^(a[167] & b[96])^(a[166] & b[97])^(a[165] & b[98])^(a[164] & b[99])^(a[163] & b[100])^(a[162] & b[101])^(a[161] & b[102])^(a[160] & b[103])^(a[159] & b[104])^(a[158] & b[105])^(a[157] & b[106])^(a[156] & b[107])^(a[155] & b[108])^(a[154] & b[109])^(a[153] & b[110])^(a[152] & b[111])^(a[151] & b[112])^(a[150] & b[113])^(a[149] & b[114])^(a[148] & b[115])^(a[147] & b[116])^(a[146] & b[117])^(a[145] & b[118])^(a[144] & b[119])^(a[143] & b[120])^(a[142] & b[121])^(a[141] & b[122])^(a[140] & b[123])^(a[139] & b[124])^(a[138] & b[125])^(a[137] & b[126])^(a[136] & b[127])^(a[135] & b[128])^(a[134] & b[129])^(a[133] & b[130])^(a[132] & b[131])^(a[131] & b[132])^(a[130] & b[133])^(a[129] & b[134])^(a[128] & b[135])^(a[127] & b[136])^(a[126] & b[137])^(a[125] & b[138])^(a[124] & b[139])^(a[123] & b[140])^(a[122] & b[141])^(a[121] & b[142])^(a[120] & b[143])^(a[119] & b[144])^(a[118] & b[145])^(a[117] & b[146])^(a[116] & b[147])^(a[115] & b[148])^(a[114] & b[149])^(a[113] & b[150])^(a[112] & b[151])^(a[111] & b[152])^(a[110] & b[153])^(a[109] & b[154])^(a[108] & b[155])^(a[107] & b[156])^(a[106] & b[157])^(a[105] & b[158])^(a[104] & b[159])^(a[103] & b[160])^(a[102] & b[161])^(a[101] & b[162])^(a[100] & b[163])^(a[99] & b[164])^(a[98] & b[165])^(a[97] & b[166])^(a[96] & b[167])^(a[95] & b[168])^(a[94] & b[169])^(a[93] & b[170])^(a[92] & b[171])^(a[91] & b[172])^(a[90] & b[173])^(a[89] & b[174])^(a[88] & b[175])^(a[87] & b[176])^(a[86] & b[177])^(a[85] & b[178])^(a[84] & b[179])^(a[83] & b[180])^(a[82] & b[181])^(a[81] & b[182])^(a[80] & b[183])^(a[79] & b[184])^(a[78] & b[185])^(a[77] & b[186])^(a[76] & b[187])^(a[75] & b[188])^(a[74] & b[189])^(a[73] & b[190])^(a[72] & b[191])^(a[71] & b[192])^(a[70] & b[193])^(a[69] & b[194])^(a[68] & b[195])^(a[67] & b[196])^(a[66] & b[197])^(a[65] & b[198])^(a[64] & b[199])^(a[63] & b[200])^(a[62] & b[201])^(a[61] & b[202])^(a[60] & b[203])^(a[59] & b[204])^(a[58] & b[205])^(a[57] & b[206])^(a[56] & b[207])^(a[55] & b[208])^(a[54] & b[209])^(a[53] & b[210])^(a[52] & b[211])^(a[51] & b[212])^(a[50] & b[213])^(a[49] & b[214])^(a[48] & b[215])^(a[47] & b[216])^(a[46] & b[217])^(a[45] & b[218])^(a[44] & b[219])^(a[43] & b[220])^(a[42] & b[221])^(a[41] & b[222])^(a[40] & b[223])^(a[39] & b[224])^(a[38] & b[225])^(a[37] & b[226])^(a[36] & b[227])^(a[35] & b[228])^(a[34] & b[229])^(a[33] & b[230])^(a[32] & b[231])^(a[31] & b[232]);
assign y[264] = (a[232] & b[32])^(a[231] & b[33])^(a[230] & b[34])^(a[229] & b[35])^(a[228] & b[36])^(a[227] & b[37])^(a[226] & b[38])^(a[225] & b[39])^(a[224] & b[40])^(a[223] & b[41])^(a[222] & b[42])^(a[221] & b[43])^(a[220] & b[44])^(a[219] & b[45])^(a[218] & b[46])^(a[217] & b[47])^(a[216] & b[48])^(a[215] & b[49])^(a[214] & b[50])^(a[213] & b[51])^(a[212] & b[52])^(a[211] & b[53])^(a[210] & b[54])^(a[209] & b[55])^(a[208] & b[56])^(a[207] & b[57])^(a[206] & b[58])^(a[205] & b[59])^(a[204] & b[60])^(a[203] & b[61])^(a[202] & b[62])^(a[201] & b[63])^(a[200] & b[64])^(a[199] & b[65])^(a[198] & b[66])^(a[197] & b[67])^(a[196] & b[68])^(a[195] & b[69])^(a[194] & b[70])^(a[193] & b[71])^(a[192] & b[72])^(a[191] & b[73])^(a[190] & b[74])^(a[189] & b[75])^(a[188] & b[76])^(a[187] & b[77])^(a[186] & b[78])^(a[185] & b[79])^(a[184] & b[80])^(a[183] & b[81])^(a[182] & b[82])^(a[181] & b[83])^(a[180] & b[84])^(a[179] & b[85])^(a[178] & b[86])^(a[177] & b[87])^(a[176] & b[88])^(a[175] & b[89])^(a[174] & b[90])^(a[173] & b[91])^(a[172] & b[92])^(a[171] & b[93])^(a[170] & b[94])^(a[169] & b[95])^(a[168] & b[96])^(a[167] & b[97])^(a[166] & b[98])^(a[165] & b[99])^(a[164] & b[100])^(a[163] & b[101])^(a[162] & b[102])^(a[161] & b[103])^(a[160] & b[104])^(a[159] & b[105])^(a[158] & b[106])^(a[157] & b[107])^(a[156] & b[108])^(a[155] & b[109])^(a[154] & b[110])^(a[153] & b[111])^(a[152] & b[112])^(a[151] & b[113])^(a[150] & b[114])^(a[149] & b[115])^(a[148] & b[116])^(a[147] & b[117])^(a[146] & b[118])^(a[145] & b[119])^(a[144] & b[120])^(a[143] & b[121])^(a[142] & b[122])^(a[141] & b[123])^(a[140] & b[124])^(a[139] & b[125])^(a[138] & b[126])^(a[137] & b[127])^(a[136] & b[128])^(a[135] & b[129])^(a[134] & b[130])^(a[133] & b[131])^(a[132] & b[132])^(a[131] & b[133])^(a[130] & b[134])^(a[129] & b[135])^(a[128] & b[136])^(a[127] & b[137])^(a[126] & b[138])^(a[125] & b[139])^(a[124] & b[140])^(a[123] & b[141])^(a[122] & b[142])^(a[121] & b[143])^(a[120] & b[144])^(a[119] & b[145])^(a[118] & b[146])^(a[117] & b[147])^(a[116] & b[148])^(a[115] & b[149])^(a[114] & b[150])^(a[113] & b[151])^(a[112] & b[152])^(a[111] & b[153])^(a[110] & b[154])^(a[109] & b[155])^(a[108] & b[156])^(a[107] & b[157])^(a[106] & b[158])^(a[105] & b[159])^(a[104] & b[160])^(a[103] & b[161])^(a[102] & b[162])^(a[101] & b[163])^(a[100] & b[164])^(a[99] & b[165])^(a[98] & b[166])^(a[97] & b[167])^(a[96] & b[168])^(a[95] & b[169])^(a[94] & b[170])^(a[93] & b[171])^(a[92] & b[172])^(a[91] & b[173])^(a[90] & b[174])^(a[89] & b[175])^(a[88] & b[176])^(a[87] & b[177])^(a[86] & b[178])^(a[85] & b[179])^(a[84] & b[180])^(a[83] & b[181])^(a[82] & b[182])^(a[81] & b[183])^(a[80] & b[184])^(a[79] & b[185])^(a[78] & b[186])^(a[77] & b[187])^(a[76] & b[188])^(a[75] & b[189])^(a[74] & b[190])^(a[73] & b[191])^(a[72] & b[192])^(a[71] & b[193])^(a[70] & b[194])^(a[69] & b[195])^(a[68] & b[196])^(a[67] & b[197])^(a[66] & b[198])^(a[65] & b[199])^(a[64] & b[200])^(a[63] & b[201])^(a[62] & b[202])^(a[61] & b[203])^(a[60] & b[204])^(a[59] & b[205])^(a[58] & b[206])^(a[57] & b[207])^(a[56] & b[208])^(a[55] & b[209])^(a[54] & b[210])^(a[53] & b[211])^(a[52] & b[212])^(a[51] & b[213])^(a[50] & b[214])^(a[49] & b[215])^(a[48] & b[216])^(a[47] & b[217])^(a[46] & b[218])^(a[45] & b[219])^(a[44] & b[220])^(a[43] & b[221])^(a[42] & b[222])^(a[41] & b[223])^(a[40] & b[224])^(a[39] & b[225])^(a[38] & b[226])^(a[37] & b[227])^(a[36] & b[228])^(a[35] & b[229])^(a[34] & b[230])^(a[33] & b[231])^(a[32] & b[232]);
assign y[265] = (a[232] & b[33])^(a[231] & b[34])^(a[230] & b[35])^(a[229] & b[36])^(a[228] & b[37])^(a[227] & b[38])^(a[226] & b[39])^(a[225] & b[40])^(a[224] & b[41])^(a[223] & b[42])^(a[222] & b[43])^(a[221] & b[44])^(a[220] & b[45])^(a[219] & b[46])^(a[218] & b[47])^(a[217] & b[48])^(a[216] & b[49])^(a[215] & b[50])^(a[214] & b[51])^(a[213] & b[52])^(a[212] & b[53])^(a[211] & b[54])^(a[210] & b[55])^(a[209] & b[56])^(a[208] & b[57])^(a[207] & b[58])^(a[206] & b[59])^(a[205] & b[60])^(a[204] & b[61])^(a[203] & b[62])^(a[202] & b[63])^(a[201] & b[64])^(a[200] & b[65])^(a[199] & b[66])^(a[198] & b[67])^(a[197] & b[68])^(a[196] & b[69])^(a[195] & b[70])^(a[194] & b[71])^(a[193] & b[72])^(a[192] & b[73])^(a[191] & b[74])^(a[190] & b[75])^(a[189] & b[76])^(a[188] & b[77])^(a[187] & b[78])^(a[186] & b[79])^(a[185] & b[80])^(a[184] & b[81])^(a[183] & b[82])^(a[182] & b[83])^(a[181] & b[84])^(a[180] & b[85])^(a[179] & b[86])^(a[178] & b[87])^(a[177] & b[88])^(a[176] & b[89])^(a[175] & b[90])^(a[174] & b[91])^(a[173] & b[92])^(a[172] & b[93])^(a[171] & b[94])^(a[170] & b[95])^(a[169] & b[96])^(a[168] & b[97])^(a[167] & b[98])^(a[166] & b[99])^(a[165] & b[100])^(a[164] & b[101])^(a[163] & b[102])^(a[162] & b[103])^(a[161] & b[104])^(a[160] & b[105])^(a[159] & b[106])^(a[158] & b[107])^(a[157] & b[108])^(a[156] & b[109])^(a[155] & b[110])^(a[154] & b[111])^(a[153] & b[112])^(a[152] & b[113])^(a[151] & b[114])^(a[150] & b[115])^(a[149] & b[116])^(a[148] & b[117])^(a[147] & b[118])^(a[146] & b[119])^(a[145] & b[120])^(a[144] & b[121])^(a[143] & b[122])^(a[142] & b[123])^(a[141] & b[124])^(a[140] & b[125])^(a[139] & b[126])^(a[138] & b[127])^(a[137] & b[128])^(a[136] & b[129])^(a[135] & b[130])^(a[134] & b[131])^(a[133] & b[132])^(a[132] & b[133])^(a[131] & b[134])^(a[130] & b[135])^(a[129] & b[136])^(a[128] & b[137])^(a[127] & b[138])^(a[126] & b[139])^(a[125] & b[140])^(a[124] & b[141])^(a[123] & b[142])^(a[122] & b[143])^(a[121] & b[144])^(a[120] & b[145])^(a[119] & b[146])^(a[118] & b[147])^(a[117] & b[148])^(a[116] & b[149])^(a[115] & b[150])^(a[114] & b[151])^(a[113] & b[152])^(a[112] & b[153])^(a[111] & b[154])^(a[110] & b[155])^(a[109] & b[156])^(a[108] & b[157])^(a[107] & b[158])^(a[106] & b[159])^(a[105] & b[160])^(a[104] & b[161])^(a[103] & b[162])^(a[102] & b[163])^(a[101] & b[164])^(a[100] & b[165])^(a[99] & b[166])^(a[98] & b[167])^(a[97] & b[168])^(a[96] & b[169])^(a[95] & b[170])^(a[94] & b[171])^(a[93] & b[172])^(a[92] & b[173])^(a[91] & b[174])^(a[90] & b[175])^(a[89] & b[176])^(a[88] & b[177])^(a[87] & b[178])^(a[86] & b[179])^(a[85] & b[180])^(a[84] & b[181])^(a[83] & b[182])^(a[82] & b[183])^(a[81] & b[184])^(a[80] & b[185])^(a[79] & b[186])^(a[78] & b[187])^(a[77] & b[188])^(a[76] & b[189])^(a[75] & b[190])^(a[74] & b[191])^(a[73] & b[192])^(a[72] & b[193])^(a[71] & b[194])^(a[70] & b[195])^(a[69] & b[196])^(a[68] & b[197])^(a[67] & b[198])^(a[66] & b[199])^(a[65] & b[200])^(a[64] & b[201])^(a[63] & b[202])^(a[62] & b[203])^(a[61] & b[204])^(a[60] & b[205])^(a[59] & b[206])^(a[58] & b[207])^(a[57] & b[208])^(a[56] & b[209])^(a[55] & b[210])^(a[54] & b[211])^(a[53] & b[212])^(a[52] & b[213])^(a[51] & b[214])^(a[50] & b[215])^(a[49] & b[216])^(a[48] & b[217])^(a[47] & b[218])^(a[46] & b[219])^(a[45] & b[220])^(a[44] & b[221])^(a[43] & b[222])^(a[42] & b[223])^(a[41] & b[224])^(a[40] & b[225])^(a[39] & b[226])^(a[38] & b[227])^(a[37] & b[228])^(a[36] & b[229])^(a[35] & b[230])^(a[34] & b[231])^(a[33] & b[232]);
assign y[266] = (a[232] & b[34])^(a[231] & b[35])^(a[230] & b[36])^(a[229] & b[37])^(a[228] & b[38])^(a[227] & b[39])^(a[226] & b[40])^(a[225] & b[41])^(a[224] & b[42])^(a[223] & b[43])^(a[222] & b[44])^(a[221] & b[45])^(a[220] & b[46])^(a[219] & b[47])^(a[218] & b[48])^(a[217] & b[49])^(a[216] & b[50])^(a[215] & b[51])^(a[214] & b[52])^(a[213] & b[53])^(a[212] & b[54])^(a[211] & b[55])^(a[210] & b[56])^(a[209] & b[57])^(a[208] & b[58])^(a[207] & b[59])^(a[206] & b[60])^(a[205] & b[61])^(a[204] & b[62])^(a[203] & b[63])^(a[202] & b[64])^(a[201] & b[65])^(a[200] & b[66])^(a[199] & b[67])^(a[198] & b[68])^(a[197] & b[69])^(a[196] & b[70])^(a[195] & b[71])^(a[194] & b[72])^(a[193] & b[73])^(a[192] & b[74])^(a[191] & b[75])^(a[190] & b[76])^(a[189] & b[77])^(a[188] & b[78])^(a[187] & b[79])^(a[186] & b[80])^(a[185] & b[81])^(a[184] & b[82])^(a[183] & b[83])^(a[182] & b[84])^(a[181] & b[85])^(a[180] & b[86])^(a[179] & b[87])^(a[178] & b[88])^(a[177] & b[89])^(a[176] & b[90])^(a[175] & b[91])^(a[174] & b[92])^(a[173] & b[93])^(a[172] & b[94])^(a[171] & b[95])^(a[170] & b[96])^(a[169] & b[97])^(a[168] & b[98])^(a[167] & b[99])^(a[166] & b[100])^(a[165] & b[101])^(a[164] & b[102])^(a[163] & b[103])^(a[162] & b[104])^(a[161] & b[105])^(a[160] & b[106])^(a[159] & b[107])^(a[158] & b[108])^(a[157] & b[109])^(a[156] & b[110])^(a[155] & b[111])^(a[154] & b[112])^(a[153] & b[113])^(a[152] & b[114])^(a[151] & b[115])^(a[150] & b[116])^(a[149] & b[117])^(a[148] & b[118])^(a[147] & b[119])^(a[146] & b[120])^(a[145] & b[121])^(a[144] & b[122])^(a[143] & b[123])^(a[142] & b[124])^(a[141] & b[125])^(a[140] & b[126])^(a[139] & b[127])^(a[138] & b[128])^(a[137] & b[129])^(a[136] & b[130])^(a[135] & b[131])^(a[134] & b[132])^(a[133] & b[133])^(a[132] & b[134])^(a[131] & b[135])^(a[130] & b[136])^(a[129] & b[137])^(a[128] & b[138])^(a[127] & b[139])^(a[126] & b[140])^(a[125] & b[141])^(a[124] & b[142])^(a[123] & b[143])^(a[122] & b[144])^(a[121] & b[145])^(a[120] & b[146])^(a[119] & b[147])^(a[118] & b[148])^(a[117] & b[149])^(a[116] & b[150])^(a[115] & b[151])^(a[114] & b[152])^(a[113] & b[153])^(a[112] & b[154])^(a[111] & b[155])^(a[110] & b[156])^(a[109] & b[157])^(a[108] & b[158])^(a[107] & b[159])^(a[106] & b[160])^(a[105] & b[161])^(a[104] & b[162])^(a[103] & b[163])^(a[102] & b[164])^(a[101] & b[165])^(a[100] & b[166])^(a[99] & b[167])^(a[98] & b[168])^(a[97] & b[169])^(a[96] & b[170])^(a[95] & b[171])^(a[94] & b[172])^(a[93] & b[173])^(a[92] & b[174])^(a[91] & b[175])^(a[90] & b[176])^(a[89] & b[177])^(a[88] & b[178])^(a[87] & b[179])^(a[86] & b[180])^(a[85] & b[181])^(a[84] & b[182])^(a[83] & b[183])^(a[82] & b[184])^(a[81] & b[185])^(a[80] & b[186])^(a[79] & b[187])^(a[78] & b[188])^(a[77] & b[189])^(a[76] & b[190])^(a[75] & b[191])^(a[74] & b[192])^(a[73] & b[193])^(a[72] & b[194])^(a[71] & b[195])^(a[70] & b[196])^(a[69] & b[197])^(a[68] & b[198])^(a[67] & b[199])^(a[66] & b[200])^(a[65] & b[201])^(a[64] & b[202])^(a[63] & b[203])^(a[62] & b[204])^(a[61] & b[205])^(a[60] & b[206])^(a[59] & b[207])^(a[58] & b[208])^(a[57] & b[209])^(a[56] & b[210])^(a[55] & b[211])^(a[54] & b[212])^(a[53] & b[213])^(a[52] & b[214])^(a[51] & b[215])^(a[50] & b[216])^(a[49] & b[217])^(a[48] & b[218])^(a[47] & b[219])^(a[46] & b[220])^(a[45] & b[221])^(a[44] & b[222])^(a[43] & b[223])^(a[42] & b[224])^(a[41] & b[225])^(a[40] & b[226])^(a[39] & b[227])^(a[38] & b[228])^(a[37] & b[229])^(a[36] & b[230])^(a[35] & b[231])^(a[34] & b[232]);
assign y[267] = (a[232] & b[35])^(a[231] & b[36])^(a[230] & b[37])^(a[229] & b[38])^(a[228] & b[39])^(a[227] & b[40])^(a[226] & b[41])^(a[225] & b[42])^(a[224] & b[43])^(a[223] & b[44])^(a[222] & b[45])^(a[221] & b[46])^(a[220] & b[47])^(a[219] & b[48])^(a[218] & b[49])^(a[217] & b[50])^(a[216] & b[51])^(a[215] & b[52])^(a[214] & b[53])^(a[213] & b[54])^(a[212] & b[55])^(a[211] & b[56])^(a[210] & b[57])^(a[209] & b[58])^(a[208] & b[59])^(a[207] & b[60])^(a[206] & b[61])^(a[205] & b[62])^(a[204] & b[63])^(a[203] & b[64])^(a[202] & b[65])^(a[201] & b[66])^(a[200] & b[67])^(a[199] & b[68])^(a[198] & b[69])^(a[197] & b[70])^(a[196] & b[71])^(a[195] & b[72])^(a[194] & b[73])^(a[193] & b[74])^(a[192] & b[75])^(a[191] & b[76])^(a[190] & b[77])^(a[189] & b[78])^(a[188] & b[79])^(a[187] & b[80])^(a[186] & b[81])^(a[185] & b[82])^(a[184] & b[83])^(a[183] & b[84])^(a[182] & b[85])^(a[181] & b[86])^(a[180] & b[87])^(a[179] & b[88])^(a[178] & b[89])^(a[177] & b[90])^(a[176] & b[91])^(a[175] & b[92])^(a[174] & b[93])^(a[173] & b[94])^(a[172] & b[95])^(a[171] & b[96])^(a[170] & b[97])^(a[169] & b[98])^(a[168] & b[99])^(a[167] & b[100])^(a[166] & b[101])^(a[165] & b[102])^(a[164] & b[103])^(a[163] & b[104])^(a[162] & b[105])^(a[161] & b[106])^(a[160] & b[107])^(a[159] & b[108])^(a[158] & b[109])^(a[157] & b[110])^(a[156] & b[111])^(a[155] & b[112])^(a[154] & b[113])^(a[153] & b[114])^(a[152] & b[115])^(a[151] & b[116])^(a[150] & b[117])^(a[149] & b[118])^(a[148] & b[119])^(a[147] & b[120])^(a[146] & b[121])^(a[145] & b[122])^(a[144] & b[123])^(a[143] & b[124])^(a[142] & b[125])^(a[141] & b[126])^(a[140] & b[127])^(a[139] & b[128])^(a[138] & b[129])^(a[137] & b[130])^(a[136] & b[131])^(a[135] & b[132])^(a[134] & b[133])^(a[133] & b[134])^(a[132] & b[135])^(a[131] & b[136])^(a[130] & b[137])^(a[129] & b[138])^(a[128] & b[139])^(a[127] & b[140])^(a[126] & b[141])^(a[125] & b[142])^(a[124] & b[143])^(a[123] & b[144])^(a[122] & b[145])^(a[121] & b[146])^(a[120] & b[147])^(a[119] & b[148])^(a[118] & b[149])^(a[117] & b[150])^(a[116] & b[151])^(a[115] & b[152])^(a[114] & b[153])^(a[113] & b[154])^(a[112] & b[155])^(a[111] & b[156])^(a[110] & b[157])^(a[109] & b[158])^(a[108] & b[159])^(a[107] & b[160])^(a[106] & b[161])^(a[105] & b[162])^(a[104] & b[163])^(a[103] & b[164])^(a[102] & b[165])^(a[101] & b[166])^(a[100] & b[167])^(a[99] & b[168])^(a[98] & b[169])^(a[97] & b[170])^(a[96] & b[171])^(a[95] & b[172])^(a[94] & b[173])^(a[93] & b[174])^(a[92] & b[175])^(a[91] & b[176])^(a[90] & b[177])^(a[89] & b[178])^(a[88] & b[179])^(a[87] & b[180])^(a[86] & b[181])^(a[85] & b[182])^(a[84] & b[183])^(a[83] & b[184])^(a[82] & b[185])^(a[81] & b[186])^(a[80] & b[187])^(a[79] & b[188])^(a[78] & b[189])^(a[77] & b[190])^(a[76] & b[191])^(a[75] & b[192])^(a[74] & b[193])^(a[73] & b[194])^(a[72] & b[195])^(a[71] & b[196])^(a[70] & b[197])^(a[69] & b[198])^(a[68] & b[199])^(a[67] & b[200])^(a[66] & b[201])^(a[65] & b[202])^(a[64] & b[203])^(a[63] & b[204])^(a[62] & b[205])^(a[61] & b[206])^(a[60] & b[207])^(a[59] & b[208])^(a[58] & b[209])^(a[57] & b[210])^(a[56] & b[211])^(a[55] & b[212])^(a[54] & b[213])^(a[53] & b[214])^(a[52] & b[215])^(a[51] & b[216])^(a[50] & b[217])^(a[49] & b[218])^(a[48] & b[219])^(a[47] & b[220])^(a[46] & b[221])^(a[45] & b[222])^(a[44] & b[223])^(a[43] & b[224])^(a[42] & b[225])^(a[41] & b[226])^(a[40] & b[227])^(a[39] & b[228])^(a[38] & b[229])^(a[37] & b[230])^(a[36] & b[231])^(a[35] & b[232]);
assign y[268] = (a[232] & b[36])^(a[231] & b[37])^(a[230] & b[38])^(a[229] & b[39])^(a[228] & b[40])^(a[227] & b[41])^(a[226] & b[42])^(a[225] & b[43])^(a[224] & b[44])^(a[223] & b[45])^(a[222] & b[46])^(a[221] & b[47])^(a[220] & b[48])^(a[219] & b[49])^(a[218] & b[50])^(a[217] & b[51])^(a[216] & b[52])^(a[215] & b[53])^(a[214] & b[54])^(a[213] & b[55])^(a[212] & b[56])^(a[211] & b[57])^(a[210] & b[58])^(a[209] & b[59])^(a[208] & b[60])^(a[207] & b[61])^(a[206] & b[62])^(a[205] & b[63])^(a[204] & b[64])^(a[203] & b[65])^(a[202] & b[66])^(a[201] & b[67])^(a[200] & b[68])^(a[199] & b[69])^(a[198] & b[70])^(a[197] & b[71])^(a[196] & b[72])^(a[195] & b[73])^(a[194] & b[74])^(a[193] & b[75])^(a[192] & b[76])^(a[191] & b[77])^(a[190] & b[78])^(a[189] & b[79])^(a[188] & b[80])^(a[187] & b[81])^(a[186] & b[82])^(a[185] & b[83])^(a[184] & b[84])^(a[183] & b[85])^(a[182] & b[86])^(a[181] & b[87])^(a[180] & b[88])^(a[179] & b[89])^(a[178] & b[90])^(a[177] & b[91])^(a[176] & b[92])^(a[175] & b[93])^(a[174] & b[94])^(a[173] & b[95])^(a[172] & b[96])^(a[171] & b[97])^(a[170] & b[98])^(a[169] & b[99])^(a[168] & b[100])^(a[167] & b[101])^(a[166] & b[102])^(a[165] & b[103])^(a[164] & b[104])^(a[163] & b[105])^(a[162] & b[106])^(a[161] & b[107])^(a[160] & b[108])^(a[159] & b[109])^(a[158] & b[110])^(a[157] & b[111])^(a[156] & b[112])^(a[155] & b[113])^(a[154] & b[114])^(a[153] & b[115])^(a[152] & b[116])^(a[151] & b[117])^(a[150] & b[118])^(a[149] & b[119])^(a[148] & b[120])^(a[147] & b[121])^(a[146] & b[122])^(a[145] & b[123])^(a[144] & b[124])^(a[143] & b[125])^(a[142] & b[126])^(a[141] & b[127])^(a[140] & b[128])^(a[139] & b[129])^(a[138] & b[130])^(a[137] & b[131])^(a[136] & b[132])^(a[135] & b[133])^(a[134] & b[134])^(a[133] & b[135])^(a[132] & b[136])^(a[131] & b[137])^(a[130] & b[138])^(a[129] & b[139])^(a[128] & b[140])^(a[127] & b[141])^(a[126] & b[142])^(a[125] & b[143])^(a[124] & b[144])^(a[123] & b[145])^(a[122] & b[146])^(a[121] & b[147])^(a[120] & b[148])^(a[119] & b[149])^(a[118] & b[150])^(a[117] & b[151])^(a[116] & b[152])^(a[115] & b[153])^(a[114] & b[154])^(a[113] & b[155])^(a[112] & b[156])^(a[111] & b[157])^(a[110] & b[158])^(a[109] & b[159])^(a[108] & b[160])^(a[107] & b[161])^(a[106] & b[162])^(a[105] & b[163])^(a[104] & b[164])^(a[103] & b[165])^(a[102] & b[166])^(a[101] & b[167])^(a[100] & b[168])^(a[99] & b[169])^(a[98] & b[170])^(a[97] & b[171])^(a[96] & b[172])^(a[95] & b[173])^(a[94] & b[174])^(a[93] & b[175])^(a[92] & b[176])^(a[91] & b[177])^(a[90] & b[178])^(a[89] & b[179])^(a[88] & b[180])^(a[87] & b[181])^(a[86] & b[182])^(a[85] & b[183])^(a[84] & b[184])^(a[83] & b[185])^(a[82] & b[186])^(a[81] & b[187])^(a[80] & b[188])^(a[79] & b[189])^(a[78] & b[190])^(a[77] & b[191])^(a[76] & b[192])^(a[75] & b[193])^(a[74] & b[194])^(a[73] & b[195])^(a[72] & b[196])^(a[71] & b[197])^(a[70] & b[198])^(a[69] & b[199])^(a[68] & b[200])^(a[67] & b[201])^(a[66] & b[202])^(a[65] & b[203])^(a[64] & b[204])^(a[63] & b[205])^(a[62] & b[206])^(a[61] & b[207])^(a[60] & b[208])^(a[59] & b[209])^(a[58] & b[210])^(a[57] & b[211])^(a[56] & b[212])^(a[55] & b[213])^(a[54] & b[214])^(a[53] & b[215])^(a[52] & b[216])^(a[51] & b[217])^(a[50] & b[218])^(a[49] & b[219])^(a[48] & b[220])^(a[47] & b[221])^(a[46] & b[222])^(a[45] & b[223])^(a[44] & b[224])^(a[43] & b[225])^(a[42] & b[226])^(a[41] & b[227])^(a[40] & b[228])^(a[39] & b[229])^(a[38] & b[230])^(a[37] & b[231])^(a[36] & b[232]);
assign y[269] = (a[232] & b[37])^(a[231] & b[38])^(a[230] & b[39])^(a[229] & b[40])^(a[228] & b[41])^(a[227] & b[42])^(a[226] & b[43])^(a[225] & b[44])^(a[224] & b[45])^(a[223] & b[46])^(a[222] & b[47])^(a[221] & b[48])^(a[220] & b[49])^(a[219] & b[50])^(a[218] & b[51])^(a[217] & b[52])^(a[216] & b[53])^(a[215] & b[54])^(a[214] & b[55])^(a[213] & b[56])^(a[212] & b[57])^(a[211] & b[58])^(a[210] & b[59])^(a[209] & b[60])^(a[208] & b[61])^(a[207] & b[62])^(a[206] & b[63])^(a[205] & b[64])^(a[204] & b[65])^(a[203] & b[66])^(a[202] & b[67])^(a[201] & b[68])^(a[200] & b[69])^(a[199] & b[70])^(a[198] & b[71])^(a[197] & b[72])^(a[196] & b[73])^(a[195] & b[74])^(a[194] & b[75])^(a[193] & b[76])^(a[192] & b[77])^(a[191] & b[78])^(a[190] & b[79])^(a[189] & b[80])^(a[188] & b[81])^(a[187] & b[82])^(a[186] & b[83])^(a[185] & b[84])^(a[184] & b[85])^(a[183] & b[86])^(a[182] & b[87])^(a[181] & b[88])^(a[180] & b[89])^(a[179] & b[90])^(a[178] & b[91])^(a[177] & b[92])^(a[176] & b[93])^(a[175] & b[94])^(a[174] & b[95])^(a[173] & b[96])^(a[172] & b[97])^(a[171] & b[98])^(a[170] & b[99])^(a[169] & b[100])^(a[168] & b[101])^(a[167] & b[102])^(a[166] & b[103])^(a[165] & b[104])^(a[164] & b[105])^(a[163] & b[106])^(a[162] & b[107])^(a[161] & b[108])^(a[160] & b[109])^(a[159] & b[110])^(a[158] & b[111])^(a[157] & b[112])^(a[156] & b[113])^(a[155] & b[114])^(a[154] & b[115])^(a[153] & b[116])^(a[152] & b[117])^(a[151] & b[118])^(a[150] & b[119])^(a[149] & b[120])^(a[148] & b[121])^(a[147] & b[122])^(a[146] & b[123])^(a[145] & b[124])^(a[144] & b[125])^(a[143] & b[126])^(a[142] & b[127])^(a[141] & b[128])^(a[140] & b[129])^(a[139] & b[130])^(a[138] & b[131])^(a[137] & b[132])^(a[136] & b[133])^(a[135] & b[134])^(a[134] & b[135])^(a[133] & b[136])^(a[132] & b[137])^(a[131] & b[138])^(a[130] & b[139])^(a[129] & b[140])^(a[128] & b[141])^(a[127] & b[142])^(a[126] & b[143])^(a[125] & b[144])^(a[124] & b[145])^(a[123] & b[146])^(a[122] & b[147])^(a[121] & b[148])^(a[120] & b[149])^(a[119] & b[150])^(a[118] & b[151])^(a[117] & b[152])^(a[116] & b[153])^(a[115] & b[154])^(a[114] & b[155])^(a[113] & b[156])^(a[112] & b[157])^(a[111] & b[158])^(a[110] & b[159])^(a[109] & b[160])^(a[108] & b[161])^(a[107] & b[162])^(a[106] & b[163])^(a[105] & b[164])^(a[104] & b[165])^(a[103] & b[166])^(a[102] & b[167])^(a[101] & b[168])^(a[100] & b[169])^(a[99] & b[170])^(a[98] & b[171])^(a[97] & b[172])^(a[96] & b[173])^(a[95] & b[174])^(a[94] & b[175])^(a[93] & b[176])^(a[92] & b[177])^(a[91] & b[178])^(a[90] & b[179])^(a[89] & b[180])^(a[88] & b[181])^(a[87] & b[182])^(a[86] & b[183])^(a[85] & b[184])^(a[84] & b[185])^(a[83] & b[186])^(a[82] & b[187])^(a[81] & b[188])^(a[80] & b[189])^(a[79] & b[190])^(a[78] & b[191])^(a[77] & b[192])^(a[76] & b[193])^(a[75] & b[194])^(a[74] & b[195])^(a[73] & b[196])^(a[72] & b[197])^(a[71] & b[198])^(a[70] & b[199])^(a[69] & b[200])^(a[68] & b[201])^(a[67] & b[202])^(a[66] & b[203])^(a[65] & b[204])^(a[64] & b[205])^(a[63] & b[206])^(a[62] & b[207])^(a[61] & b[208])^(a[60] & b[209])^(a[59] & b[210])^(a[58] & b[211])^(a[57] & b[212])^(a[56] & b[213])^(a[55] & b[214])^(a[54] & b[215])^(a[53] & b[216])^(a[52] & b[217])^(a[51] & b[218])^(a[50] & b[219])^(a[49] & b[220])^(a[48] & b[221])^(a[47] & b[222])^(a[46] & b[223])^(a[45] & b[224])^(a[44] & b[225])^(a[43] & b[226])^(a[42] & b[227])^(a[41] & b[228])^(a[40] & b[229])^(a[39] & b[230])^(a[38] & b[231])^(a[37] & b[232]);
assign y[270] = (a[232] & b[38])^(a[231] & b[39])^(a[230] & b[40])^(a[229] & b[41])^(a[228] & b[42])^(a[227] & b[43])^(a[226] & b[44])^(a[225] & b[45])^(a[224] & b[46])^(a[223] & b[47])^(a[222] & b[48])^(a[221] & b[49])^(a[220] & b[50])^(a[219] & b[51])^(a[218] & b[52])^(a[217] & b[53])^(a[216] & b[54])^(a[215] & b[55])^(a[214] & b[56])^(a[213] & b[57])^(a[212] & b[58])^(a[211] & b[59])^(a[210] & b[60])^(a[209] & b[61])^(a[208] & b[62])^(a[207] & b[63])^(a[206] & b[64])^(a[205] & b[65])^(a[204] & b[66])^(a[203] & b[67])^(a[202] & b[68])^(a[201] & b[69])^(a[200] & b[70])^(a[199] & b[71])^(a[198] & b[72])^(a[197] & b[73])^(a[196] & b[74])^(a[195] & b[75])^(a[194] & b[76])^(a[193] & b[77])^(a[192] & b[78])^(a[191] & b[79])^(a[190] & b[80])^(a[189] & b[81])^(a[188] & b[82])^(a[187] & b[83])^(a[186] & b[84])^(a[185] & b[85])^(a[184] & b[86])^(a[183] & b[87])^(a[182] & b[88])^(a[181] & b[89])^(a[180] & b[90])^(a[179] & b[91])^(a[178] & b[92])^(a[177] & b[93])^(a[176] & b[94])^(a[175] & b[95])^(a[174] & b[96])^(a[173] & b[97])^(a[172] & b[98])^(a[171] & b[99])^(a[170] & b[100])^(a[169] & b[101])^(a[168] & b[102])^(a[167] & b[103])^(a[166] & b[104])^(a[165] & b[105])^(a[164] & b[106])^(a[163] & b[107])^(a[162] & b[108])^(a[161] & b[109])^(a[160] & b[110])^(a[159] & b[111])^(a[158] & b[112])^(a[157] & b[113])^(a[156] & b[114])^(a[155] & b[115])^(a[154] & b[116])^(a[153] & b[117])^(a[152] & b[118])^(a[151] & b[119])^(a[150] & b[120])^(a[149] & b[121])^(a[148] & b[122])^(a[147] & b[123])^(a[146] & b[124])^(a[145] & b[125])^(a[144] & b[126])^(a[143] & b[127])^(a[142] & b[128])^(a[141] & b[129])^(a[140] & b[130])^(a[139] & b[131])^(a[138] & b[132])^(a[137] & b[133])^(a[136] & b[134])^(a[135] & b[135])^(a[134] & b[136])^(a[133] & b[137])^(a[132] & b[138])^(a[131] & b[139])^(a[130] & b[140])^(a[129] & b[141])^(a[128] & b[142])^(a[127] & b[143])^(a[126] & b[144])^(a[125] & b[145])^(a[124] & b[146])^(a[123] & b[147])^(a[122] & b[148])^(a[121] & b[149])^(a[120] & b[150])^(a[119] & b[151])^(a[118] & b[152])^(a[117] & b[153])^(a[116] & b[154])^(a[115] & b[155])^(a[114] & b[156])^(a[113] & b[157])^(a[112] & b[158])^(a[111] & b[159])^(a[110] & b[160])^(a[109] & b[161])^(a[108] & b[162])^(a[107] & b[163])^(a[106] & b[164])^(a[105] & b[165])^(a[104] & b[166])^(a[103] & b[167])^(a[102] & b[168])^(a[101] & b[169])^(a[100] & b[170])^(a[99] & b[171])^(a[98] & b[172])^(a[97] & b[173])^(a[96] & b[174])^(a[95] & b[175])^(a[94] & b[176])^(a[93] & b[177])^(a[92] & b[178])^(a[91] & b[179])^(a[90] & b[180])^(a[89] & b[181])^(a[88] & b[182])^(a[87] & b[183])^(a[86] & b[184])^(a[85] & b[185])^(a[84] & b[186])^(a[83] & b[187])^(a[82] & b[188])^(a[81] & b[189])^(a[80] & b[190])^(a[79] & b[191])^(a[78] & b[192])^(a[77] & b[193])^(a[76] & b[194])^(a[75] & b[195])^(a[74] & b[196])^(a[73] & b[197])^(a[72] & b[198])^(a[71] & b[199])^(a[70] & b[200])^(a[69] & b[201])^(a[68] & b[202])^(a[67] & b[203])^(a[66] & b[204])^(a[65] & b[205])^(a[64] & b[206])^(a[63] & b[207])^(a[62] & b[208])^(a[61] & b[209])^(a[60] & b[210])^(a[59] & b[211])^(a[58] & b[212])^(a[57] & b[213])^(a[56] & b[214])^(a[55] & b[215])^(a[54] & b[216])^(a[53] & b[217])^(a[52] & b[218])^(a[51] & b[219])^(a[50] & b[220])^(a[49] & b[221])^(a[48] & b[222])^(a[47] & b[223])^(a[46] & b[224])^(a[45] & b[225])^(a[44] & b[226])^(a[43] & b[227])^(a[42] & b[228])^(a[41] & b[229])^(a[40] & b[230])^(a[39] & b[231])^(a[38] & b[232]);
assign y[271] = (a[232] & b[39])^(a[231] & b[40])^(a[230] & b[41])^(a[229] & b[42])^(a[228] & b[43])^(a[227] & b[44])^(a[226] & b[45])^(a[225] & b[46])^(a[224] & b[47])^(a[223] & b[48])^(a[222] & b[49])^(a[221] & b[50])^(a[220] & b[51])^(a[219] & b[52])^(a[218] & b[53])^(a[217] & b[54])^(a[216] & b[55])^(a[215] & b[56])^(a[214] & b[57])^(a[213] & b[58])^(a[212] & b[59])^(a[211] & b[60])^(a[210] & b[61])^(a[209] & b[62])^(a[208] & b[63])^(a[207] & b[64])^(a[206] & b[65])^(a[205] & b[66])^(a[204] & b[67])^(a[203] & b[68])^(a[202] & b[69])^(a[201] & b[70])^(a[200] & b[71])^(a[199] & b[72])^(a[198] & b[73])^(a[197] & b[74])^(a[196] & b[75])^(a[195] & b[76])^(a[194] & b[77])^(a[193] & b[78])^(a[192] & b[79])^(a[191] & b[80])^(a[190] & b[81])^(a[189] & b[82])^(a[188] & b[83])^(a[187] & b[84])^(a[186] & b[85])^(a[185] & b[86])^(a[184] & b[87])^(a[183] & b[88])^(a[182] & b[89])^(a[181] & b[90])^(a[180] & b[91])^(a[179] & b[92])^(a[178] & b[93])^(a[177] & b[94])^(a[176] & b[95])^(a[175] & b[96])^(a[174] & b[97])^(a[173] & b[98])^(a[172] & b[99])^(a[171] & b[100])^(a[170] & b[101])^(a[169] & b[102])^(a[168] & b[103])^(a[167] & b[104])^(a[166] & b[105])^(a[165] & b[106])^(a[164] & b[107])^(a[163] & b[108])^(a[162] & b[109])^(a[161] & b[110])^(a[160] & b[111])^(a[159] & b[112])^(a[158] & b[113])^(a[157] & b[114])^(a[156] & b[115])^(a[155] & b[116])^(a[154] & b[117])^(a[153] & b[118])^(a[152] & b[119])^(a[151] & b[120])^(a[150] & b[121])^(a[149] & b[122])^(a[148] & b[123])^(a[147] & b[124])^(a[146] & b[125])^(a[145] & b[126])^(a[144] & b[127])^(a[143] & b[128])^(a[142] & b[129])^(a[141] & b[130])^(a[140] & b[131])^(a[139] & b[132])^(a[138] & b[133])^(a[137] & b[134])^(a[136] & b[135])^(a[135] & b[136])^(a[134] & b[137])^(a[133] & b[138])^(a[132] & b[139])^(a[131] & b[140])^(a[130] & b[141])^(a[129] & b[142])^(a[128] & b[143])^(a[127] & b[144])^(a[126] & b[145])^(a[125] & b[146])^(a[124] & b[147])^(a[123] & b[148])^(a[122] & b[149])^(a[121] & b[150])^(a[120] & b[151])^(a[119] & b[152])^(a[118] & b[153])^(a[117] & b[154])^(a[116] & b[155])^(a[115] & b[156])^(a[114] & b[157])^(a[113] & b[158])^(a[112] & b[159])^(a[111] & b[160])^(a[110] & b[161])^(a[109] & b[162])^(a[108] & b[163])^(a[107] & b[164])^(a[106] & b[165])^(a[105] & b[166])^(a[104] & b[167])^(a[103] & b[168])^(a[102] & b[169])^(a[101] & b[170])^(a[100] & b[171])^(a[99] & b[172])^(a[98] & b[173])^(a[97] & b[174])^(a[96] & b[175])^(a[95] & b[176])^(a[94] & b[177])^(a[93] & b[178])^(a[92] & b[179])^(a[91] & b[180])^(a[90] & b[181])^(a[89] & b[182])^(a[88] & b[183])^(a[87] & b[184])^(a[86] & b[185])^(a[85] & b[186])^(a[84] & b[187])^(a[83] & b[188])^(a[82] & b[189])^(a[81] & b[190])^(a[80] & b[191])^(a[79] & b[192])^(a[78] & b[193])^(a[77] & b[194])^(a[76] & b[195])^(a[75] & b[196])^(a[74] & b[197])^(a[73] & b[198])^(a[72] & b[199])^(a[71] & b[200])^(a[70] & b[201])^(a[69] & b[202])^(a[68] & b[203])^(a[67] & b[204])^(a[66] & b[205])^(a[65] & b[206])^(a[64] & b[207])^(a[63] & b[208])^(a[62] & b[209])^(a[61] & b[210])^(a[60] & b[211])^(a[59] & b[212])^(a[58] & b[213])^(a[57] & b[214])^(a[56] & b[215])^(a[55] & b[216])^(a[54] & b[217])^(a[53] & b[218])^(a[52] & b[219])^(a[51] & b[220])^(a[50] & b[221])^(a[49] & b[222])^(a[48] & b[223])^(a[47] & b[224])^(a[46] & b[225])^(a[45] & b[226])^(a[44] & b[227])^(a[43] & b[228])^(a[42] & b[229])^(a[41] & b[230])^(a[40] & b[231])^(a[39] & b[232]);
assign y[272] = (a[232] & b[40])^(a[231] & b[41])^(a[230] & b[42])^(a[229] & b[43])^(a[228] & b[44])^(a[227] & b[45])^(a[226] & b[46])^(a[225] & b[47])^(a[224] & b[48])^(a[223] & b[49])^(a[222] & b[50])^(a[221] & b[51])^(a[220] & b[52])^(a[219] & b[53])^(a[218] & b[54])^(a[217] & b[55])^(a[216] & b[56])^(a[215] & b[57])^(a[214] & b[58])^(a[213] & b[59])^(a[212] & b[60])^(a[211] & b[61])^(a[210] & b[62])^(a[209] & b[63])^(a[208] & b[64])^(a[207] & b[65])^(a[206] & b[66])^(a[205] & b[67])^(a[204] & b[68])^(a[203] & b[69])^(a[202] & b[70])^(a[201] & b[71])^(a[200] & b[72])^(a[199] & b[73])^(a[198] & b[74])^(a[197] & b[75])^(a[196] & b[76])^(a[195] & b[77])^(a[194] & b[78])^(a[193] & b[79])^(a[192] & b[80])^(a[191] & b[81])^(a[190] & b[82])^(a[189] & b[83])^(a[188] & b[84])^(a[187] & b[85])^(a[186] & b[86])^(a[185] & b[87])^(a[184] & b[88])^(a[183] & b[89])^(a[182] & b[90])^(a[181] & b[91])^(a[180] & b[92])^(a[179] & b[93])^(a[178] & b[94])^(a[177] & b[95])^(a[176] & b[96])^(a[175] & b[97])^(a[174] & b[98])^(a[173] & b[99])^(a[172] & b[100])^(a[171] & b[101])^(a[170] & b[102])^(a[169] & b[103])^(a[168] & b[104])^(a[167] & b[105])^(a[166] & b[106])^(a[165] & b[107])^(a[164] & b[108])^(a[163] & b[109])^(a[162] & b[110])^(a[161] & b[111])^(a[160] & b[112])^(a[159] & b[113])^(a[158] & b[114])^(a[157] & b[115])^(a[156] & b[116])^(a[155] & b[117])^(a[154] & b[118])^(a[153] & b[119])^(a[152] & b[120])^(a[151] & b[121])^(a[150] & b[122])^(a[149] & b[123])^(a[148] & b[124])^(a[147] & b[125])^(a[146] & b[126])^(a[145] & b[127])^(a[144] & b[128])^(a[143] & b[129])^(a[142] & b[130])^(a[141] & b[131])^(a[140] & b[132])^(a[139] & b[133])^(a[138] & b[134])^(a[137] & b[135])^(a[136] & b[136])^(a[135] & b[137])^(a[134] & b[138])^(a[133] & b[139])^(a[132] & b[140])^(a[131] & b[141])^(a[130] & b[142])^(a[129] & b[143])^(a[128] & b[144])^(a[127] & b[145])^(a[126] & b[146])^(a[125] & b[147])^(a[124] & b[148])^(a[123] & b[149])^(a[122] & b[150])^(a[121] & b[151])^(a[120] & b[152])^(a[119] & b[153])^(a[118] & b[154])^(a[117] & b[155])^(a[116] & b[156])^(a[115] & b[157])^(a[114] & b[158])^(a[113] & b[159])^(a[112] & b[160])^(a[111] & b[161])^(a[110] & b[162])^(a[109] & b[163])^(a[108] & b[164])^(a[107] & b[165])^(a[106] & b[166])^(a[105] & b[167])^(a[104] & b[168])^(a[103] & b[169])^(a[102] & b[170])^(a[101] & b[171])^(a[100] & b[172])^(a[99] & b[173])^(a[98] & b[174])^(a[97] & b[175])^(a[96] & b[176])^(a[95] & b[177])^(a[94] & b[178])^(a[93] & b[179])^(a[92] & b[180])^(a[91] & b[181])^(a[90] & b[182])^(a[89] & b[183])^(a[88] & b[184])^(a[87] & b[185])^(a[86] & b[186])^(a[85] & b[187])^(a[84] & b[188])^(a[83] & b[189])^(a[82] & b[190])^(a[81] & b[191])^(a[80] & b[192])^(a[79] & b[193])^(a[78] & b[194])^(a[77] & b[195])^(a[76] & b[196])^(a[75] & b[197])^(a[74] & b[198])^(a[73] & b[199])^(a[72] & b[200])^(a[71] & b[201])^(a[70] & b[202])^(a[69] & b[203])^(a[68] & b[204])^(a[67] & b[205])^(a[66] & b[206])^(a[65] & b[207])^(a[64] & b[208])^(a[63] & b[209])^(a[62] & b[210])^(a[61] & b[211])^(a[60] & b[212])^(a[59] & b[213])^(a[58] & b[214])^(a[57] & b[215])^(a[56] & b[216])^(a[55] & b[217])^(a[54] & b[218])^(a[53] & b[219])^(a[52] & b[220])^(a[51] & b[221])^(a[50] & b[222])^(a[49] & b[223])^(a[48] & b[224])^(a[47] & b[225])^(a[46] & b[226])^(a[45] & b[227])^(a[44] & b[228])^(a[43] & b[229])^(a[42] & b[230])^(a[41] & b[231])^(a[40] & b[232]);
assign y[273] = (a[232] & b[41])^(a[231] & b[42])^(a[230] & b[43])^(a[229] & b[44])^(a[228] & b[45])^(a[227] & b[46])^(a[226] & b[47])^(a[225] & b[48])^(a[224] & b[49])^(a[223] & b[50])^(a[222] & b[51])^(a[221] & b[52])^(a[220] & b[53])^(a[219] & b[54])^(a[218] & b[55])^(a[217] & b[56])^(a[216] & b[57])^(a[215] & b[58])^(a[214] & b[59])^(a[213] & b[60])^(a[212] & b[61])^(a[211] & b[62])^(a[210] & b[63])^(a[209] & b[64])^(a[208] & b[65])^(a[207] & b[66])^(a[206] & b[67])^(a[205] & b[68])^(a[204] & b[69])^(a[203] & b[70])^(a[202] & b[71])^(a[201] & b[72])^(a[200] & b[73])^(a[199] & b[74])^(a[198] & b[75])^(a[197] & b[76])^(a[196] & b[77])^(a[195] & b[78])^(a[194] & b[79])^(a[193] & b[80])^(a[192] & b[81])^(a[191] & b[82])^(a[190] & b[83])^(a[189] & b[84])^(a[188] & b[85])^(a[187] & b[86])^(a[186] & b[87])^(a[185] & b[88])^(a[184] & b[89])^(a[183] & b[90])^(a[182] & b[91])^(a[181] & b[92])^(a[180] & b[93])^(a[179] & b[94])^(a[178] & b[95])^(a[177] & b[96])^(a[176] & b[97])^(a[175] & b[98])^(a[174] & b[99])^(a[173] & b[100])^(a[172] & b[101])^(a[171] & b[102])^(a[170] & b[103])^(a[169] & b[104])^(a[168] & b[105])^(a[167] & b[106])^(a[166] & b[107])^(a[165] & b[108])^(a[164] & b[109])^(a[163] & b[110])^(a[162] & b[111])^(a[161] & b[112])^(a[160] & b[113])^(a[159] & b[114])^(a[158] & b[115])^(a[157] & b[116])^(a[156] & b[117])^(a[155] & b[118])^(a[154] & b[119])^(a[153] & b[120])^(a[152] & b[121])^(a[151] & b[122])^(a[150] & b[123])^(a[149] & b[124])^(a[148] & b[125])^(a[147] & b[126])^(a[146] & b[127])^(a[145] & b[128])^(a[144] & b[129])^(a[143] & b[130])^(a[142] & b[131])^(a[141] & b[132])^(a[140] & b[133])^(a[139] & b[134])^(a[138] & b[135])^(a[137] & b[136])^(a[136] & b[137])^(a[135] & b[138])^(a[134] & b[139])^(a[133] & b[140])^(a[132] & b[141])^(a[131] & b[142])^(a[130] & b[143])^(a[129] & b[144])^(a[128] & b[145])^(a[127] & b[146])^(a[126] & b[147])^(a[125] & b[148])^(a[124] & b[149])^(a[123] & b[150])^(a[122] & b[151])^(a[121] & b[152])^(a[120] & b[153])^(a[119] & b[154])^(a[118] & b[155])^(a[117] & b[156])^(a[116] & b[157])^(a[115] & b[158])^(a[114] & b[159])^(a[113] & b[160])^(a[112] & b[161])^(a[111] & b[162])^(a[110] & b[163])^(a[109] & b[164])^(a[108] & b[165])^(a[107] & b[166])^(a[106] & b[167])^(a[105] & b[168])^(a[104] & b[169])^(a[103] & b[170])^(a[102] & b[171])^(a[101] & b[172])^(a[100] & b[173])^(a[99] & b[174])^(a[98] & b[175])^(a[97] & b[176])^(a[96] & b[177])^(a[95] & b[178])^(a[94] & b[179])^(a[93] & b[180])^(a[92] & b[181])^(a[91] & b[182])^(a[90] & b[183])^(a[89] & b[184])^(a[88] & b[185])^(a[87] & b[186])^(a[86] & b[187])^(a[85] & b[188])^(a[84] & b[189])^(a[83] & b[190])^(a[82] & b[191])^(a[81] & b[192])^(a[80] & b[193])^(a[79] & b[194])^(a[78] & b[195])^(a[77] & b[196])^(a[76] & b[197])^(a[75] & b[198])^(a[74] & b[199])^(a[73] & b[200])^(a[72] & b[201])^(a[71] & b[202])^(a[70] & b[203])^(a[69] & b[204])^(a[68] & b[205])^(a[67] & b[206])^(a[66] & b[207])^(a[65] & b[208])^(a[64] & b[209])^(a[63] & b[210])^(a[62] & b[211])^(a[61] & b[212])^(a[60] & b[213])^(a[59] & b[214])^(a[58] & b[215])^(a[57] & b[216])^(a[56] & b[217])^(a[55] & b[218])^(a[54] & b[219])^(a[53] & b[220])^(a[52] & b[221])^(a[51] & b[222])^(a[50] & b[223])^(a[49] & b[224])^(a[48] & b[225])^(a[47] & b[226])^(a[46] & b[227])^(a[45] & b[228])^(a[44] & b[229])^(a[43] & b[230])^(a[42] & b[231])^(a[41] & b[232]);
assign y[274] = (a[232] & b[42])^(a[231] & b[43])^(a[230] & b[44])^(a[229] & b[45])^(a[228] & b[46])^(a[227] & b[47])^(a[226] & b[48])^(a[225] & b[49])^(a[224] & b[50])^(a[223] & b[51])^(a[222] & b[52])^(a[221] & b[53])^(a[220] & b[54])^(a[219] & b[55])^(a[218] & b[56])^(a[217] & b[57])^(a[216] & b[58])^(a[215] & b[59])^(a[214] & b[60])^(a[213] & b[61])^(a[212] & b[62])^(a[211] & b[63])^(a[210] & b[64])^(a[209] & b[65])^(a[208] & b[66])^(a[207] & b[67])^(a[206] & b[68])^(a[205] & b[69])^(a[204] & b[70])^(a[203] & b[71])^(a[202] & b[72])^(a[201] & b[73])^(a[200] & b[74])^(a[199] & b[75])^(a[198] & b[76])^(a[197] & b[77])^(a[196] & b[78])^(a[195] & b[79])^(a[194] & b[80])^(a[193] & b[81])^(a[192] & b[82])^(a[191] & b[83])^(a[190] & b[84])^(a[189] & b[85])^(a[188] & b[86])^(a[187] & b[87])^(a[186] & b[88])^(a[185] & b[89])^(a[184] & b[90])^(a[183] & b[91])^(a[182] & b[92])^(a[181] & b[93])^(a[180] & b[94])^(a[179] & b[95])^(a[178] & b[96])^(a[177] & b[97])^(a[176] & b[98])^(a[175] & b[99])^(a[174] & b[100])^(a[173] & b[101])^(a[172] & b[102])^(a[171] & b[103])^(a[170] & b[104])^(a[169] & b[105])^(a[168] & b[106])^(a[167] & b[107])^(a[166] & b[108])^(a[165] & b[109])^(a[164] & b[110])^(a[163] & b[111])^(a[162] & b[112])^(a[161] & b[113])^(a[160] & b[114])^(a[159] & b[115])^(a[158] & b[116])^(a[157] & b[117])^(a[156] & b[118])^(a[155] & b[119])^(a[154] & b[120])^(a[153] & b[121])^(a[152] & b[122])^(a[151] & b[123])^(a[150] & b[124])^(a[149] & b[125])^(a[148] & b[126])^(a[147] & b[127])^(a[146] & b[128])^(a[145] & b[129])^(a[144] & b[130])^(a[143] & b[131])^(a[142] & b[132])^(a[141] & b[133])^(a[140] & b[134])^(a[139] & b[135])^(a[138] & b[136])^(a[137] & b[137])^(a[136] & b[138])^(a[135] & b[139])^(a[134] & b[140])^(a[133] & b[141])^(a[132] & b[142])^(a[131] & b[143])^(a[130] & b[144])^(a[129] & b[145])^(a[128] & b[146])^(a[127] & b[147])^(a[126] & b[148])^(a[125] & b[149])^(a[124] & b[150])^(a[123] & b[151])^(a[122] & b[152])^(a[121] & b[153])^(a[120] & b[154])^(a[119] & b[155])^(a[118] & b[156])^(a[117] & b[157])^(a[116] & b[158])^(a[115] & b[159])^(a[114] & b[160])^(a[113] & b[161])^(a[112] & b[162])^(a[111] & b[163])^(a[110] & b[164])^(a[109] & b[165])^(a[108] & b[166])^(a[107] & b[167])^(a[106] & b[168])^(a[105] & b[169])^(a[104] & b[170])^(a[103] & b[171])^(a[102] & b[172])^(a[101] & b[173])^(a[100] & b[174])^(a[99] & b[175])^(a[98] & b[176])^(a[97] & b[177])^(a[96] & b[178])^(a[95] & b[179])^(a[94] & b[180])^(a[93] & b[181])^(a[92] & b[182])^(a[91] & b[183])^(a[90] & b[184])^(a[89] & b[185])^(a[88] & b[186])^(a[87] & b[187])^(a[86] & b[188])^(a[85] & b[189])^(a[84] & b[190])^(a[83] & b[191])^(a[82] & b[192])^(a[81] & b[193])^(a[80] & b[194])^(a[79] & b[195])^(a[78] & b[196])^(a[77] & b[197])^(a[76] & b[198])^(a[75] & b[199])^(a[74] & b[200])^(a[73] & b[201])^(a[72] & b[202])^(a[71] & b[203])^(a[70] & b[204])^(a[69] & b[205])^(a[68] & b[206])^(a[67] & b[207])^(a[66] & b[208])^(a[65] & b[209])^(a[64] & b[210])^(a[63] & b[211])^(a[62] & b[212])^(a[61] & b[213])^(a[60] & b[214])^(a[59] & b[215])^(a[58] & b[216])^(a[57] & b[217])^(a[56] & b[218])^(a[55] & b[219])^(a[54] & b[220])^(a[53] & b[221])^(a[52] & b[222])^(a[51] & b[223])^(a[50] & b[224])^(a[49] & b[225])^(a[48] & b[226])^(a[47] & b[227])^(a[46] & b[228])^(a[45] & b[229])^(a[44] & b[230])^(a[43] & b[231])^(a[42] & b[232]);
assign y[275] = (a[232] & b[43])^(a[231] & b[44])^(a[230] & b[45])^(a[229] & b[46])^(a[228] & b[47])^(a[227] & b[48])^(a[226] & b[49])^(a[225] & b[50])^(a[224] & b[51])^(a[223] & b[52])^(a[222] & b[53])^(a[221] & b[54])^(a[220] & b[55])^(a[219] & b[56])^(a[218] & b[57])^(a[217] & b[58])^(a[216] & b[59])^(a[215] & b[60])^(a[214] & b[61])^(a[213] & b[62])^(a[212] & b[63])^(a[211] & b[64])^(a[210] & b[65])^(a[209] & b[66])^(a[208] & b[67])^(a[207] & b[68])^(a[206] & b[69])^(a[205] & b[70])^(a[204] & b[71])^(a[203] & b[72])^(a[202] & b[73])^(a[201] & b[74])^(a[200] & b[75])^(a[199] & b[76])^(a[198] & b[77])^(a[197] & b[78])^(a[196] & b[79])^(a[195] & b[80])^(a[194] & b[81])^(a[193] & b[82])^(a[192] & b[83])^(a[191] & b[84])^(a[190] & b[85])^(a[189] & b[86])^(a[188] & b[87])^(a[187] & b[88])^(a[186] & b[89])^(a[185] & b[90])^(a[184] & b[91])^(a[183] & b[92])^(a[182] & b[93])^(a[181] & b[94])^(a[180] & b[95])^(a[179] & b[96])^(a[178] & b[97])^(a[177] & b[98])^(a[176] & b[99])^(a[175] & b[100])^(a[174] & b[101])^(a[173] & b[102])^(a[172] & b[103])^(a[171] & b[104])^(a[170] & b[105])^(a[169] & b[106])^(a[168] & b[107])^(a[167] & b[108])^(a[166] & b[109])^(a[165] & b[110])^(a[164] & b[111])^(a[163] & b[112])^(a[162] & b[113])^(a[161] & b[114])^(a[160] & b[115])^(a[159] & b[116])^(a[158] & b[117])^(a[157] & b[118])^(a[156] & b[119])^(a[155] & b[120])^(a[154] & b[121])^(a[153] & b[122])^(a[152] & b[123])^(a[151] & b[124])^(a[150] & b[125])^(a[149] & b[126])^(a[148] & b[127])^(a[147] & b[128])^(a[146] & b[129])^(a[145] & b[130])^(a[144] & b[131])^(a[143] & b[132])^(a[142] & b[133])^(a[141] & b[134])^(a[140] & b[135])^(a[139] & b[136])^(a[138] & b[137])^(a[137] & b[138])^(a[136] & b[139])^(a[135] & b[140])^(a[134] & b[141])^(a[133] & b[142])^(a[132] & b[143])^(a[131] & b[144])^(a[130] & b[145])^(a[129] & b[146])^(a[128] & b[147])^(a[127] & b[148])^(a[126] & b[149])^(a[125] & b[150])^(a[124] & b[151])^(a[123] & b[152])^(a[122] & b[153])^(a[121] & b[154])^(a[120] & b[155])^(a[119] & b[156])^(a[118] & b[157])^(a[117] & b[158])^(a[116] & b[159])^(a[115] & b[160])^(a[114] & b[161])^(a[113] & b[162])^(a[112] & b[163])^(a[111] & b[164])^(a[110] & b[165])^(a[109] & b[166])^(a[108] & b[167])^(a[107] & b[168])^(a[106] & b[169])^(a[105] & b[170])^(a[104] & b[171])^(a[103] & b[172])^(a[102] & b[173])^(a[101] & b[174])^(a[100] & b[175])^(a[99] & b[176])^(a[98] & b[177])^(a[97] & b[178])^(a[96] & b[179])^(a[95] & b[180])^(a[94] & b[181])^(a[93] & b[182])^(a[92] & b[183])^(a[91] & b[184])^(a[90] & b[185])^(a[89] & b[186])^(a[88] & b[187])^(a[87] & b[188])^(a[86] & b[189])^(a[85] & b[190])^(a[84] & b[191])^(a[83] & b[192])^(a[82] & b[193])^(a[81] & b[194])^(a[80] & b[195])^(a[79] & b[196])^(a[78] & b[197])^(a[77] & b[198])^(a[76] & b[199])^(a[75] & b[200])^(a[74] & b[201])^(a[73] & b[202])^(a[72] & b[203])^(a[71] & b[204])^(a[70] & b[205])^(a[69] & b[206])^(a[68] & b[207])^(a[67] & b[208])^(a[66] & b[209])^(a[65] & b[210])^(a[64] & b[211])^(a[63] & b[212])^(a[62] & b[213])^(a[61] & b[214])^(a[60] & b[215])^(a[59] & b[216])^(a[58] & b[217])^(a[57] & b[218])^(a[56] & b[219])^(a[55] & b[220])^(a[54] & b[221])^(a[53] & b[222])^(a[52] & b[223])^(a[51] & b[224])^(a[50] & b[225])^(a[49] & b[226])^(a[48] & b[227])^(a[47] & b[228])^(a[46] & b[229])^(a[45] & b[230])^(a[44] & b[231])^(a[43] & b[232]);
assign y[276] = (a[232] & b[44])^(a[231] & b[45])^(a[230] & b[46])^(a[229] & b[47])^(a[228] & b[48])^(a[227] & b[49])^(a[226] & b[50])^(a[225] & b[51])^(a[224] & b[52])^(a[223] & b[53])^(a[222] & b[54])^(a[221] & b[55])^(a[220] & b[56])^(a[219] & b[57])^(a[218] & b[58])^(a[217] & b[59])^(a[216] & b[60])^(a[215] & b[61])^(a[214] & b[62])^(a[213] & b[63])^(a[212] & b[64])^(a[211] & b[65])^(a[210] & b[66])^(a[209] & b[67])^(a[208] & b[68])^(a[207] & b[69])^(a[206] & b[70])^(a[205] & b[71])^(a[204] & b[72])^(a[203] & b[73])^(a[202] & b[74])^(a[201] & b[75])^(a[200] & b[76])^(a[199] & b[77])^(a[198] & b[78])^(a[197] & b[79])^(a[196] & b[80])^(a[195] & b[81])^(a[194] & b[82])^(a[193] & b[83])^(a[192] & b[84])^(a[191] & b[85])^(a[190] & b[86])^(a[189] & b[87])^(a[188] & b[88])^(a[187] & b[89])^(a[186] & b[90])^(a[185] & b[91])^(a[184] & b[92])^(a[183] & b[93])^(a[182] & b[94])^(a[181] & b[95])^(a[180] & b[96])^(a[179] & b[97])^(a[178] & b[98])^(a[177] & b[99])^(a[176] & b[100])^(a[175] & b[101])^(a[174] & b[102])^(a[173] & b[103])^(a[172] & b[104])^(a[171] & b[105])^(a[170] & b[106])^(a[169] & b[107])^(a[168] & b[108])^(a[167] & b[109])^(a[166] & b[110])^(a[165] & b[111])^(a[164] & b[112])^(a[163] & b[113])^(a[162] & b[114])^(a[161] & b[115])^(a[160] & b[116])^(a[159] & b[117])^(a[158] & b[118])^(a[157] & b[119])^(a[156] & b[120])^(a[155] & b[121])^(a[154] & b[122])^(a[153] & b[123])^(a[152] & b[124])^(a[151] & b[125])^(a[150] & b[126])^(a[149] & b[127])^(a[148] & b[128])^(a[147] & b[129])^(a[146] & b[130])^(a[145] & b[131])^(a[144] & b[132])^(a[143] & b[133])^(a[142] & b[134])^(a[141] & b[135])^(a[140] & b[136])^(a[139] & b[137])^(a[138] & b[138])^(a[137] & b[139])^(a[136] & b[140])^(a[135] & b[141])^(a[134] & b[142])^(a[133] & b[143])^(a[132] & b[144])^(a[131] & b[145])^(a[130] & b[146])^(a[129] & b[147])^(a[128] & b[148])^(a[127] & b[149])^(a[126] & b[150])^(a[125] & b[151])^(a[124] & b[152])^(a[123] & b[153])^(a[122] & b[154])^(a[121] & b[155])^(a[120] & b[156])^(a[119] & b[157])^(a[118] & b[158])^(a[117] & b[159])^(a[116] & b[160])^(a[115] & b[161])^(a[114] & b[162])^(a[113] & b[163])^(a[112] & b[164])^(a[111] & b[165])^(a[110] & b[166])^(a[109] & b[167])^(a[108] & b[168])^(a[107] & b[169])^(a[106] & b[170])^(a[105] & b[171])^(a[104] & b[172])^(a[103] & b[173])^(a[102] & b[174])^(a[101] & b[175])^(a[100] & b[176])^(a[99] & b[177])^(a[98] & b[178])^(a[97] & b[179])^(a[96] & b[180])^(a[95] & b[181])^(a[94] & b[182])^(a[93] & b[183])^(a[92] & b[184])^(a[91] & b[185])^(a[90] & b[186])^(a[89] & b[187])^(a[88] & b[188])^(a[87] & b[189])^(a[86] & b[190])^(a[85] & b[191])^(a[84] & b[192])^(a[83] & b[193])^(a[82] & b[194])^(a[81] & b[195])^(a[80] & b[196])^(a[79] & b[197])^(a[78] & b[198])^(a[77] & b[199])^(a[76] & b[200])^(a[75] & b[201])^(a[74] & b[202])^(a[73] & b[203])^(a[72] & b[204])^(a[71] & b[205])^(a[70] & b[206])^(a[69] & b[207])^(a[68] & b[208])^(a[67] & b[209])^(a[66] & b[210])^(a[65] & b[211])^(a[64] & b[212])^(a[63] & b[213])^(a[62] & b[214])^(a[61] & b[215])^(a[60] & b[216])^(a[59] & b[217])^(a[58] & b[218])^(a[57] & b[219])^(a[56] & b[220])^(a[55] & b[221])^(a[54] & b[222])^(a[53] & b[223])^(a[52] & b[224])^(a[51] & b[225])^(a[50] & b[226])^(a[49] & b[227])^(a[48] & b[228])^(a[47] & b[229])^(a[46] & b[230])^(a[45] & b[231])^(a[44] & b[232]);
assign y[277] = (a[232] & b[45])^(a[231] & b[46])^(a[230] & b[47])^(a[229] & b[48])^(a[228] & b[49])^(a[227] & b[50])^(a[226] & b[51])^(a[225] & b[52])^(a[224] & b[53])^(a[223] & b[54])^(a[222] & b[55])^(a[221] & b[56])^(a[220] & b[57])^(a[219] & b[58])^(a[218] & b[59])^(a[217] & b[60])^(a[216] & b[61])^(a[215] & b[62])^(a[214] & b[63])^(a[213] & b[64])^(a[212] & b[65])^(a[211] & b[66])^(a[210] & b[67])^(a[209] & b[68])^(a[208] & b[69])^(a[207] & b[70])^(a[206] & b[71])^(a[205] & b[72])^(a[204] & b[73])^(a[203] & b[74])^(a[202] & b[75])^(a[201] & b[76])^(a[200] & b[77])^(a[199] & b[78])^(a[198] & b[79])^(a[197] & b[80])^(a[196] & b[81])^(a[195] & b[82])^(a[194] & b[83])^(a[193] & b[84])^(a[192] & b[85])^(a[191] & b[86])^(a[190] & b[87])^(a[189] & b[88])^(a[188] & b[89])^(a[187] & b[90])^(a[186] & b[91])^(a[185] & b[92])^(a[184] & b[93])^(a[183] & b[94])^(a[182] & b[95])^(a[181] & b[96])^(a[180] & b[97])^(a[179] & b[98])^(a[178] & b[99])^(a[177] & b[100])^(a[176] & b[101])^(a[175] & b[102])^(a[174] & b[103])^(a[173] & b[104])^(a[172] & b[105])^(a[171] & b[106])^(a[170] & b[107])^(a[169] & b[108])^(a[168] & b[109])^(a[167] & b[110])^(a[166] & b[111])^(a[165] & b[112])^(a[164] & b[113])^(a[163] & b[114])^(a[162] & b[115])^(a[161] & b[116])^(a[160] & b[117])^(a[159] & b[118])^(a[158] & b[119])^(a[157] & b[120])^(a[156] & b[121])^(a[155] & b[122])^(a[154] & b[123])^(a[153] & b[124])^(a[152] & b[125])^(a[151] & b[126])^(a[150] & b[127])^(a[149] & b[128])^(a[148] & b[129])^(a[147] & b[130])^(a[146] & b[131])^(a[145] & b[132])^(a[144] & b[133])^(a[143] & b[134])^(a[142] & b[135])^(a[141] & b[136])^(a[140] & b[137])^(a[139] & b[138])^(a[138] & b[139])^(a[137] & b[140])^(a[136] & b[141])^(a[135] & b[142])^(a[134] & b[143])^(a[133] & b[144])^(a[132] & b[145])^(a[131] & b[146])^(a[130] & b[147])^(a[129] & b[148])^(a[128] & b[149])^(a[127] & b[150])^(a[126] & b[151])^(a[125] & b[152])^(a[124] & b[153])^(a[123] & b[154])^(a[122] & b[155])^(a[121] & b[156])^(a[120] & b[157])^(a[119] & b[158])^(a[118] & b[159])^(a[117] & b[160])^(a[116] & b[161])^(a[115] & b[162])^(a[114] & b[163])^(a[113] & b[164])^(a[112] & b[165])^(a[111] & b[166])^(a[110] & b[167])^(a[109] & b[168])^(a[108] & b[169])^(a[107] & b[170])^(a[106] & b[171])^(a[105] & b[172])^(a[104] & b[173])^(a[103] & b[174])^(a[102] & b[175])^(a[101] & b[176])^(a[100] & b[177])^(a[99] & b[178])^(a[98] & b[179])^(a[97] & b[180])^(a[96] & b[181])^(a[95] & b[182])^(a[94] & b[183])^(a[93] & b[184])^(a[92] & b[185])^(a[91] & b[186])^(a[90] & b[187])^(a[89] & b[188])^(a[88] & b[189])^(a[87] & b[190])^(a[86] & b[191])^(a[85] & b[192])^(a[84] & b[193])^(a[83] & b[194])^(a[82] & b[195])^(a[81] & b[196])^(a[80] & b[197])^(a[79] & b[198])^(a[78] & b[199])^(a[77] & b[200])^(a[76] & b[201])^(a[75] & b[202])^(a[74] & b[203])^(a[73] & b[204])^(a[72] & b[205])^(a[71] & b[206])^(a[70] & b[207])^(a[69] & b[208])^(a[68] & b[209])^(a[67] & b[210])^(a[66] & b[211])^(a[65] & b[212])^(a[64] & b[213])^(a[63] & b[214])^(a[62] & b[215])^(a[61] & b[216])^(a[60] & b[217])^(a[59] & b[218])^(a[58] & b[219])^(a[57] & b[220])^(a[56] & b[221])^(a[55] & b[222])^(a[54] & b[223])^(a[53] & b[224])^(a[52] & b[225])^(a[51] & b[226])^(a[50] & b[227])^(a[49] & b[228])^(a[48] & b[229])^(a[47] & b[230])^(a[46] & b[231])^(a[45] & b[232]);
assign y[278] = (a[232] & b[46])^(a[231] & b[47])^(a[230] & b[48])^(a[229] & b[49])^(a[228] & b[50])^(a[227] & b[51])^(a[226] & b[52])^(a[225] & b[53])^(a[224] & b[54])^(a[223] & b[55])^(a[222] & b[56])^(a[221] & b[57])^(a[220] & b[58])^(a[219] & b[59])^(a[218] & b[60])^(a[217] & b[61])^(a[216] & b[62])^(a[215] & b[63])^(a[214] & b[64])^(a[213] & b[65])^(a[212] & b[66])^(a[211] & b[67])^(a[210] & b[68])^(a[209] & b[69])^(a[208] & b[70])^(a[207] & b[71])^(a[206] & b[72])^(a[205] & b[73])^(a[204] & b[74])^(a[203] & b[75])^(a[202] & b[76])^(a[201] & b[77])^(a[200] & b[78])^(a[199] & b[79])^(a[198] & b[80])^(a[197] & b[81])^(a[196] & b[82])^(a[195] & b[83])^(a[194] & b[84])^(a[193] & b[85])^(a[192] & b[86])^(a[191] & b[87])^(a[190] & b[88])^(a[189] & b[89])^(a[188] & b[90])^(a[187] & b[91])^(a[186] & b[92])^(a[185] & b[93])^(a[184] & b[94])^(a[183] & b[95])^(a[182] & b[96])^(a[181] & b[97])^(a[180] & b[98])^(a[179] & b[99])^(a[178] & b[100])^(a[177] & b[101])^(a[176] & b[102])^(a[175] & b[103])^(a[174] & b[104])^(a[173] & b[105])^(a[172] & b[106])^(a[171] & b[107])^(a[170] & b[108])^(a[169] & b[109])^(a[168] & b[110])^(a[167] & b[111])^(a[166] & b[112])^(a[165] & b[113])^(a[164] & b[114])^(a[163] & b[115])^(a[162] & b[116])^(a[161] & b[117])^(a[160] & b[118])^(a[159] & b[119])^(a[158] & b[120])^(a[157] & b[121])^(a[156] & b[122])^(a[155] & b[123])^(a[154] & b[124])^(a[153] & b[125])^(a[152] & b[126])^(a[151] & b[127])^(a[150] & b[128])^(a[149] & b[129])^(a[148] & b[130])^(a[147] & b[131])^(a[146] & b[132])^(a[145] & b[133])^(a[144] & b[134])^(a[143] & b[135])^(a[142] & b[136])^(a[141] & b[137])^(a[140] & b[138])^(a[139] & b[139])^(a[138] & b[140])^(a[137] & b[141])^(a[136] & b[142])^(a[135] & b[143])^(a[134] & b[144])^(a[133] & b[145])^(a[132] & b[146])^(a[131] & b[147])^(a[130] & b[148])^(a[129] & b[149])^(a[128] & b[150])^(a[127] & b[151])^(a[126] & b[152])^(a[125] & b[153])^(a[124] & b[154])^(a[123] & b[155])^(a[122] & b[156])^(a[121] & b[157])^(a[120] & b[158])^(a[119] & b[159])^(a[118] & b[160])^(a[117] & b[161])^(a[116] & b[162])^(a[115] & b[163])^(a[114] & b[164])^(a[113] & b[165])^(a[112] & b[166])^(a[111] & b[167])^(a[110] & b[168])^(a[109] & b[169])^(a[108] & b[170])^(a[107] & b[171])^(a[106] & b[172])^(a[105] & b[173])^(a[104] & b[174])^(a[103] & b[175])^(a[102] & b[176])^(a[101] & b[177])^(a[100] & b[178])^(a[99] & b[179])^(a[98] & b[180])^(a[97] & b[181])^(a[96] & b[182])^(a[95] & b[183])^(a[94] & b[184])^(a[93] & b[185])^(a[92] & b[186])^(a[91] & b[187])^(a[90] & b[188])^(a[89] & b[189])^(a[88] & b[190])^(a[87] & b[191])^(a[86] & b[192])^(a[85] & b[193])^(a[84] & b[194])^(a[83] & b[195])^(a[82] & b[196])^(a[81] & b[197])^(a[80] & b[198])^(a[79] & b[199])^(a[78] & b[200])^(a[77] & b[201])^(a[76] & b[202])^(a[75] & b[203])^(a[74] & b[204])^(a[73] & b[205])^(a[72] & b[206])^(a[71] & b[207])^(a[70] & b[208])^(a[69] & b[209])^(a[68] & b[210])^(a[67] & b[211])^(a[66] & b[212])^(a[65] & b[213])^(a[64] & b[214])^(a[63] & b[215])^(a[62] & b[216])^(a[61] & b[217])^(a[60] & b[218])^(a[59] & b[219])^(a[58] & b[220])^(a[57] & b[221])^(a[56] & b[222])^(a[55] & b[223])^(a[54] & b[224])^(a[53] & b[225])^(a[52] & b[226])^(a[51] & b[227])^(a[50] & b[228])^(a[49] & b[229])^(a[48] & b[230])^(a[47] & b[231])^(a[46] & b[232]);
assign y[279] = (a[232] & b[47])^(a[231] & b[48])^(a[230] & b[49])^(a[229] & b[50])^(a[228] & b[51])^(a[227] & b[52])^(a[226] & b[53])^(a[225] & b[54])^(a[224] & b[55])^(a[223] & b[56])^(a[222] & b[57])^(a[221] & b[58])^(a[220] & b[59])^(a[219] & b[60])^(a[218] & b[61])^(a[217] & b[62])^(a[216] & b[63])^(a[215] & b[64])^(a[214] & b[65])^(a[213] & b[66])^(a[212] & b[67])^(a[211] & b[68])^(a[210] & b[69])^(a[209] & b[70])^(a[208] & b[71])^(a[207] & b[72])^(a[206] & b[73])^(a[205] & b[74])^(a[204] & b[75])^(a[203] & b[76])^(a[202] & b[77])^(a[201] & b[78])^(a[200] & b[79])^(a[199] & b[80])^(a[198] & b[81])^(a[197] & b[82])^(a[196] & b[83])^(a[195] & b[84])^(a[194] & b[85])^(a[193] & b[86])^(a[192] & b[87])^(a[191] & b[88])^(a[190] & b[89])^(a[189] & b[90])^(a[188] & b[91])^(a[187] & b[92])^(a[186] & b[93])^(a[185] & b[94])^(a[184] & b[95])^(a[183] & b[96])^(a[182] & b[97])^(a[181] & b[98])^(a[180] & b[99])^(a[179] & b[100])^(a[178] & b[101])^(a[177] & b[102])^(a[176] & b[103])^(a[175] & b[104])^(a[174] & b[105])^(a[173] & b[106])^(a[172] & b[107])^(a[171] & b[108])^(a[170] & b[109])^(a[169] & b[110])^(a[168] & b[111])^(a[167] & b[112])^(a[166] & b[113])^(a[165] & b[114])^(a[164] & b[115])^(a[163] & b[116])^(a[162] & b[117])^(a[161] & b[118])^(a[160] & b[119])^(a[159] & b[120])^(a[158] & b[121])^(a[157] & b[122])^(a[156] & b[123])^(a[155] & b[124])^(a[154] & b[125])^(a[153] & b[126])^(a[152] & b[127])^(a[151] & b[128])^(a[150] & b[129])^(a[149] & b[130])^(a[148] & b[131])^(a[147] & b[132])^(a[146] & b[133])^(a[145] & b[134])^(a[144] & b[135])^(a[143] & b[136])^(a[142] & b[137])^(a[141] & b[138])^(a[140] & b[139])^(a[139] & b[140])^(a[138] & b[141])^(a[137] & b[142])^(a[136] & b[143])^(a[135] & b[144])^(a[134] & b[145])^(a[133] & b[146])^(a[132] & b[147])^(a[131] & b[148])^(a[130] & b[149])^(a[129] & b[150])^(a[128] & b[151])^(a[127] & b[152])^(a[126] & b[153])^(a[125] & b[154])^(a[124] & b[155])^(a[123] & b[156])^(a[122] & b[157])^(a[121] & b[158])^(a[120] & b[159])^(a[119] & b[160])^(a[118] & b[161])^(a[117] & b[162])^(a[116] & b[163])^(a[115] & b[164])^(a[114] & b[165])^(a[113] & b[166])^(a[112] & b[167])^(a[111] & b[168])^(a[110] & b[169])^(a[109] & b[170])^(a[108] & b[171])^(a[107] & b[172])^(a[106] & b[173])^(a[105] & b[174])^(a[104] & b[175])^(a[103] & b[176])^(a[102] & b[177])^(a[101] & b[178])^(a[100] & b[179])^(a[99] & b[180])^(a[98] & b[181])^(a[97] & b[182])^(a[96] & b[183])^(a[95] & b[184])^(a[94] & b[185])^(a[93] & b[186])^(a[92] & b[187])^(a[91] & b[188])^(a[90] & b[189])^(a[89] & b[190])^(a[88] & b[191])^(a[87] & b[192])^(a[86] & b[193])^(a[85] & b[194])^(a[84] & b[195])^(a[83] & b[196])^(a[82] & b[197])^(a[81] & b[198])^(a[80] & b[199])^(a[79] & b[200])^(a[78] & b[201])^(a[77] & b[202])^(a[76] & b[203])^(a[75] & b[204])^(a[74] & b[205])^(a[73] & b[206])^(a[72] & b[207])^(a[71] & b[208])^(a[70] & b[209])^(a[69] & b[210])^(a[68] & b[211])^(a[67] & b[212])^(a[66] & b[213])^(a[65] & b[214])^(a[64] & b[215])^(a[63] & b[216])^(a[62] & b[217])^(a[61] & b[218])^(a[60] & b[219])^(a[59] & b[220])^(a[58] & b[221])^(a[57] & b[222])^(a[56] & b[223])^(a[55] & b[224])^(a[54] & b[225])^(a[53] & b[226])^(a[52] & b[227])^(a[51] & b[228])^(a[50] & b[229])^(a[49] & b[230])^(a[48] & b[231])^(a[47] & b[232]);
assign y[280] = (a[232] & b[48])^(a[231] & b[49])^(a[230] & b[50])^(a[229] & b[51])^(a[228] & b[52])^(a[227] & b[53])^(a[226] & b[54])^(a[225] & b[55])^(a[224] & b[56])^(a[223] & b[57])^(a[222] & b[58])^(a[221] & b[59])^(a[220] & b[60])^(a[219] & b[61])^(a[218] & b[62])^(a[217] & b[63])^(a[216] & b[64])^(a[215] & b[65])^(a[214] & b[66])^(a[213] & b[67])^(a[212] & b[68])^(a[211] & b[69])^(a[210] & b[70])^(a[209] & b[71])^(a[208] & b[72])^(a[207] & b[73])^(a[206] & b[74])^(a[205] & b[75])^(a[204] & b[76])^(a[203] & b[77])^(a[202] & b[78])^(a[201] & b[79])^(a[200] & b[80])^(a[199] & b[81])^(a[198] & b[82])^(a[197] & b[83])^(a[196] & b[84])^(a[195] & b[85])^(a[194] & b[86])^(a[193] & b[87])^(a[192] & b[88])^(a[191] & b[89])^(a[190] & b[90])^(a[189] & b[91])^(a[188] & b[92])^(a[187] & b[93])^(a[186] & b[94])^(a[185] & b[95])^(a[184] & b[96])^(a[183] & b[97])^(a[182] & b[98])^(a[181] & b[99])^(a[180] & b[100])^(a[179] & b[101])^(a[178] & b[102])^(a[177] & b[103])^(a[176] & b[104])^(a[175] & b[105])^(a[174] & b[106])^(a[173] & b[107])^(a[172] & b[108])^(a[171] & b[109])^(a[170] & b[110])^(a[169] & b[111])^(a[168] & b[112])^(a[167] & b[113])^(a[166] & b[114])^(a[165] & b[115])^(a[164] & b[116])^(a[163] & b[117])^(a[162] & b[118])^(a[161] & b[119])^(a[160] & b[120])^(a[159] & b[121])^(a[158] & b[122])^(a[157] & b[123])^(a[156] & b[124])^(a[155] & b[125])^(a[154] & b[126])^(a[153] & b[127])^(a[152] & b[128])^(a[151] & b[129])^(a[150] & b[130])^(a[149] & b[131])^(a[148] & b[132])^(a[147] & b[133])^(a[146] & b[134])^(a[145] & b[135])^(a[144] & b[136])^(a[143] & b[137])^(a[142] & b[138])^(a[141] & b[139])^(a[140] & b[140])^(a[139] & b[141])^(a[138] & b[142])^(a[137] & b[143])^(a[136] & b[144])^(a[135] & b[145])^(a[134] & b[146])^(a[133] & b[147])^(a[132] & b[148])^(a[131] & b[149])^(a[130] & b[150])^(a[129] & b[151])^(a[128] & b[152])^(a[127] & b[153])^(a[126] & b[154])^(a[125] & b[155])^(a[124] & b[156])^(a[123] & b[157])^(a[122] & b[158])^(a[121] & b[159])^(a[120] & b[160])^(a[119] & b[161])^(a[118] & b[162])^(a[117] & b[163])^(a[116] & b[164])^(a[115] & b[165])^(a[114] & b[166])^(a[113] & b[167])^(a[112] & b[168])^(a[111] & b[169])^(a[110] & b[170])^(a[109] & b[171])^(a[108] & b[172])^(a[107] & b[173])^(a[106] & b[174])^(a[105] & b[175])^(a[104] & b[176])^(a[103] & b[177])^(a[102] & b[178])^(a[101] & b[179])^(a[100] & b[180])^(a[99] & b[181])^(a[98] & b[182])^(a[97] & b[183])^(a[96] & b[184])^(a[95] & b[185])^(a[94] & b[186])^(a[93] & b[187])^(a[92] & b[188])^(a[91] & b[189])^(a[90] & b[190])^(a[89] & b[191])^(a[88] & b[192])^(a[87] & b[193])^(a[86] & b[194])^(a[85] & b[195])^(a[84] & b[196])^(a[83] & b[197])^(a[82] & b[198])^(a[81] & b[199])^(a[80] & b[200])^(a[79] & b[201])^(a[78] & b[202])^(a[77] & b[203])^(a[76] & b[204])^(a[75] & b[205])^(a[74] & b[206])^(a[73] & b[207])^(a[72] & b[208])^(a[71] & b[209])^(a[70] & b[210])^(a[69] & b[211])^(a[68] & b[212])^(a[67] & b[213])^(a[66] & b[214])^(a[65] & b[215])^(a[64] & b[216])^(a[63] & b[217])^(a[62] & b[218])^(a[61] & b[219])^(a[60] & b[220])^(a[59] & b[221])^(a[58] & b[222])^(a[57] & b[223])^(a[56] & b[224])^(a[55] & b[225])^(a[54] & b[226])^(a[53] & b[227])^(a[52] & b[228])^(a[51] & b[229])^(a[50] & b[230])^(a[49] & b[231])^(a[48] & b[232]);
assign y[281] = (a[232] & b[49])^(a[231] & b[50])^(a[230] & b[51])^(a[229] & b[52])^(a[228] & b[53])^(a[227] & b[54])^(a[226] & b[55])^(a[225] & b[56])^(a[224] & b[57])^(a[223] & b[58])^(a[222] & b[59])^(a[221] & b[60])^(a[220] & b[61])^(a[219] & b[62])^(a[218] & b[63])^(a[217] & b[64])^(a[216] & b[65])^(a[215] & b[66])^(a[214] & b[67])^(a[213] & b[68])^(a[212] & b[69])^(a[211] & b[70])^(a[210] & b[71])^(a[209] & b[72])^(a[208] & b[73])^(a[207] & b[74])^(a[206] & b[75])^(a[205] & b[76])^(a[204] & b[77])^(a[203] & b[78])^(a[202] & b[79])^(a[201] & b[80])^(a[200] & b[81])^(a[199] & b[82])^(a[198] & b[83])^(a[197] & b[84])^(a[196] & b[85])^(a[195] & b[86])^(a[194] & b[87])^(a[193] & b[88])^(a[192] & b[89])^(a[191] & b[90])^(a[190] & b[91])^(a[189] & b[92])^(a[188] & b[93])^(a[187] & b[94])^(a[186] & b[95])^(a[185] & b[96])^(a[184] & b[97])^(a[183] & b[98])^(a[182] & b[99])^(a[181] & b[100])^(a[180] & b[101])^(a[179] & b[102])^(a[178] & b[103])^(a[177] & b[104])^(a[176] & b[105])^(a[175] & b[106])^(a[174] & b[107])^(a[173] & b[108])^(a[172] & b[109])^(a[171] & b[110])^(a[170] & b[111])^(a[169] & b[112])^(a[168] & b[113])^(a[167] & b[114])^(a[166] & b[115])^(a[165] & b[116])^(a[164] & b[117])^(a[163] & b[118])^(a[162] & b[119])^(a[161] & b[120])^(a[160] & b[121])^(a[159] & b[122])^(a[158] & b[123])^(a[157] & b[124])^(a[156] & b[125])^(a[155] & b[126])^(a[154] & b[127])^(a[153] & b[128])^(a[152] & b[129])^(a[151] & b[130])^(a[150] & b[131])^(a[149] & b[132])^(a[148] & b[133])^(a[147] & b[134])^(a[146] & b[135])^(a[145] & b[136])^(a[144] & b[137])^(a[143] & b[138])^(a[142] & b[139])^(a[141] & b[140])^(a[140] & b[141])^(a[139] & b[142])^(a[138] & b[143])^(a[137] & b[144])^(a[136] & b[145])^(a[135] & b[146])^(a[134] & b[147])^(a[133] & b[148])^(a[132] & b[149])^(a[131] & b[150])^(a[130] & b[151])^(a[129] & b[152])^(a[128] & b[153])^(a[127] & b[154])^(a[126] & b[155])^(a[125] & b[156])^(a[124] & b[157])^(a[123] & b[158])^(a[122] & b[159])^(a[121] & b[160])^(a[120] & b[161])^(a[119] & b[162])^(a[118] & b[163])^(a[117] & b[164])^(a[116] & b[165])^(a[115] & b[166])^(a[114] & b[167])^(a[113] & b[168])^(a[112] & b[169])^(a[111] & b[170])^(a[110] & b[171])^(a[109] & b[172])^(a[108] & b[173])^(a[107] & b[174])^(a[106] & b[175])^(a[105] & b[176])^(a[104] & b[177])^(a[103] & b[178])^(a[102] & b[179])^(a[101] & b[180])^(a[100] & b[181])^(a[99] & b[182])^(a[98] & b[183])^(a[97] & b[184])^(a[96] & b[185])^(a[95] & b[186])^(a[94] & b[187])^(a[93] & b[188])^(a[92] & b[189])^(a[91] & b[190])^(a[90] & b[191])^(a[89] & b[192])^(a[88] & b[193])^(a[87] & b[194])^(a[86] & b[195])^(a[85] & b[196])^(a[84] & b[197])^(a[83] & b[198])^(a[82] & b[199])^(a[81] & b[200])^(a[80] & b[201])^(a[79] & b[202])^(a[78] & b[203])^(a[77] & b[204])^(a[76] & b[205])^(a[75] & b[206])^(a[74] & b[207])^(a[73] & b[208])^(a[72] & b[209])^(a[71] & b[210])^(a[70] & b[211])^(a[69] & b[212])^(a[68] & b[213])^(a[67] & b[214])^(a[66] & b[215])^(a[65] & b[216])^(a[64] & b[217])^(a[63] & b[218])^(a[62] & b[219])^(a[61] & b[220])^(a[60] & b[221])^(a[59] & b[222])^(a[58] & b[223])^(a[57] & b[224])^(a[56] & b[225])^(a[55] & b[226])^(a[54] & b[227])^(a[53] & b[228])^(a[52] & b[229])^(a[51] & b[230])^(a[50] & b[231])^(a[49] & b[232]);
assign y[282] = (a[232] & b[50])^(a[231] & b[51])^(a[230] & b[52])^(a[229] & b[53])^(a[228] & b[54])^(a[227] & b[55])^(a[226] & b[56])^(a[225] & b[57])^(a[224] & b[58])^(a[223] & b[59])^(a[222] & b[60])^(a[221] & b[61])^(a[220] & b[62])^(a[219] & b[63])^(a[218] & b[64])^(a[217] & b[65])^(a[216] & b[66])^(a[215] & b[67])^(a[214] & b[68])^(a[213] & b[69])^(a[212] & b[70])^(a[211] & b[71])^(a[210] & b[72])^(a[209] & b[73])^(a[208] & b[74])^(a[207] & b[75])^(a[206] & b[76])^(a[205] & b[77])^(a[204] & b[78])^(a[203] & b[79])^(a[202] & b[80])^(a[201] & b[81])^(a[200] & b[82])^(a[199] & b[83])^(a[198] & b[84])^(a[197] & b[85])^(a[196] & b[86])^(a[195] & b[87])^(a[194] & b[88])^(a[193] & b[89])^(a[192] & b[90])^(a[191] & b[91])^(a[190] & b[92])^(a[189] & b[93])^(a[188] & b[94])^(a[187] & b[95])^(a[186] & b[96])^(a[185] & b[97])^(a[184] & b[98])^(a[183] & b[99])^(a[182] & b[100])^(a[181] & b[101])^(a[180] & b[102])^(a[179] & b[103])^(a[178] & b[104])^(a[177] & b[105])^(a[176] & b[106])^(a[175] & b[107])^(a[174] & b[108])^(a[173] & b[109])^(a[172] & b[110])^(a[171] & b[111])^(a[170] & b[112])^(a[169] & b[113])^(a[168] & b[114])^(a[167] & b[115])^(a[166] & b[116])^(a[165] & b[117])^(a[164] & b[118])^(a[163] & b[119])^(a[162] & b[120])^(a[161] & b[121])^(a[160] & b[122])^(a[159] & b[123])^(a[158] & b[124])^(a[157] & b[125])^(a[156] & b[126])^(a[155] & b[127])^(a[154] & b[128])^(a[153] & b[129])^(a[152] & b[130])^(a[151] & b[131])^(a[150] & b[132])^(a[149] & b[133])^(a[148] & b[134])^(a[147] & b[135])^(a[146] & b[136])^(a[145] & b[137])^(a[144] & b[138])^(a[143] & b[139])^(a[142] & b[140])^(a[141] & b[141])^(a[140] & b[142])^(a[139] & b[143])^(a[138] & b[144])^(a[137] & b[145])^(a[136] & b[146])^(a[135] & b[147])^(a[134] & b[148])^(a[133] & b[149])^(a[132] & b[150])^(a[131] & b[151])^(a[130] & b[152])^(a[129] & b[153])^(a[128] & b[154])^(a[127] & b[155])^(a[126] & b[156])^(a[125] & b[157])^(a[124] & b[158])^(a[123] & b[159])^(a[122] & b[160])^(a[121] & b[161])^(a[120] & b[162])^(a[119] & b[163])^(a[118] & b[164])^(a[117] & b[165])^(a[116] & b[166])^(a[115] & b[167])^(a[114] & b[168])^(a[113] & b[169])^(a[112] & b[170])^(a[111] & b[171])^(a[110] & b[172])^(a[109] & b[173])^(a[108] & b[174])^(a[107] & b[175])^(a[106] & b[176])^(a[105] & b[177])^(a[104] & b[178])^(a[103] & b[179])^(a[102] & b[180])^(a[101] & b[181])^(a[100] & b[182])^(a[99] & b[183])^(a[98] & b[184])^(a[97] & b[185])^(a[96] & b[186])^(a[95] & b[187])^(a[94] & b[188])^(a[93] & b[189])^(a[92] & b[190])^(a[91] & b[191])^(a[90] & b[192])^(a[89] & b[193])^(a[88] & b[194])^(a[87] & b[195])^(a[86] & b[196])^(a[85] & b[197])^(a[84] & b[198])^(a[83] & b[199])^(a[82] & b[200])^(a[81] & b[201])^(a[80] & b[202])^(a[79] & b[203])^(a[78] & b[204])^(a[77] & b[205])^(a[76] & b[206])^(a[75] & b[207])^(a[74] & b[208])^(a[73] & b[209])^(a[72] & b[210])^(a[71] & b[211])^(a[70] & b[212])^(a[69] & b[213])^(a[68] & b[214])^(a[67] & b[215])^(a[66] & b[216])^(a[65] & b[217])^(a[64] & b[218])^(a[63] & b[219])^(a[62] & b[220])^(a[61] & b[221])^(a[60] & b[222])^(a[59] & b[223])^(a[58] & b[224])^(a[57] & b[225])^(a[56] & b[226])^(a[55] & b[227])^(a[54] & b[228])^(a[53] & b[229])^(a[52] & b[230])^(a[51] & b[231])^(a[50] & b[232]);
assign y[283] = (a[232] & b[51])^(a[231] & b[52])^(a[230] & b[53])^(a[229] & b[54])^(a[228] & b[55])^(a[227] & b[56])^(a[226] & b[57])^(a[225] & b[58])^(a[224] & b[59])^(a[223] & b[60])^(a[222] & b[61])^(a[221] & b[62])^(a[220] & b[63])^(a[219] & b[64])^(a[218] & b[65])^(a[217] & b[66])^(a[216] & b[67])^(a[215] & b[68])^(a[214] & b[69])^(a[213] & b[70])^(a[212] & b[71])^(a[211] & b[72])^(a[210] & b[73])^(a[209] & b[74])^(a[208] & b[75])^(a[207] & b[76])^(a[206] & b[77])^(a[205] & b[78])^(a[204] & b[79])^(a[203] & b[80])^(a[202] & b[81])^(a[201] & b[82])^(a[200] & b[83])^(a[199] & b[84])^(a[198] & b[85])^(a[197] & b[86])^(a[196] & b[87])^(a[195] & b[88])^(a[194] & b[89])^(a[193] & b[90])^(a[192] & b[91])^(a[191] & b[92])^(a[190] & b[93])^(a[189] & b[94])^(a[188] & b[95])^(a[187] & b[96])^(a[186] & b[97])^(a[185] & b[98])^(a[184] & b[99])^(a[183] & b[100])^(a[182] & b[101])^(a[181] & b[102])^(a[180] & b[103])^(a[179] & b[104])^(a[178] & b[105])^(a[177] & b[106])^(a[176] & b[107])^(a[175] & b[108])^(a[174] & b[109])^(a[173] & b[110])^(a[172] & b[111])^(a[171] & b[112])^(a[170] & b[113])^(a[169] & b[114])^(a[168] & b[115])^(a[167] & b[116])^(a[166] & b[117])^(a[165] & b[118])^(a[164] & b[119])^(a[163] & b[120])^(a[162] & b[121])^(a[161] & b[122])^(a[160] & b[123])^(a[159] & b[124])^(a[158] & b[125])^(a[157] & b[126])^(a[156] & b[127])^(a[155] & b[128])^(a[154] & b[129])^(a[153] & b[130])^(a[152] & b[131])^(a[151] & b[132])^(a[150] & b[133])^(a[149] & b[134])^(a[148] & b[135])^(a[147] & b[136])^(a[146] & b[137])^(a[145] & b[138])^(a[144] & b[139])^(a[143] & b[140])^(a[142] & b[141])^(a[141] & b[142])^(a[140] & b[143])^(a[139] & b[144])^(a[138] & b[145])^(a[137] & b[146])^(a[136] & b[147])^(a[135] & b[148])^(a[134] & b[149])^(a[133] & b[150])^(a[132] & b[151])^(a[131] & b[152])^(a[130] & b[153])^(a[129] & b[154])^(a[128] & b[155])^(a[127] & b[156])^(a[126] & b[157])^(a[125] & b[158])^(a[124] & b[159])^(a[123] & b[160])^(a[122] & b[161])^(a[121] & b[162])^(a[120] & b[163])^(a[119] & b[164])^(a[118] & b[165])^(a[117] & b[166])^(a[116] & b[167])^(a[115] & b[168])^(a[114] & b[169])^(a[113] & b[170])^(a[112] & b[171])^(a[111] & b[172])^(a[110] & b[173])^(a[109] & b[174])^(a[108] & b[175])^(a[107] & b[176])^(a[106] & b[177])^(a[105] & b[178])^(a[104] & b[179])^(a[103] & b[180])^(a[102] & b[181])^(a[101] & b[182])^(a[100] & b[183])^(a[99] & b[184])^(a[98] & b[185])^(a[97] & b[186])^(a[96] & b[187])^(a[95] & b[188])^(a[94] & b[189])^(a[93] & b[190])^(a[92] & b[191])^(a[91] & b[192])^(a[90] & b[193])^(a[89] & b[194])^(a[88] & b[195])^(a[87] & b[196])^(a[86] & b[197])^(a[85] & b[198])^(a[84] & b[199])^(a[83] & b[200])^(a[82] & b[201])^(a[81] & b[202])^(a[80] & b[203])^(a[79] & b[204])^(a[78] & b[205])^(a[77] & b[206])^(a[76] & b[207])^(a[75] & b[208])^(a[74] & b[209])^(a[73] & b[210])^(a[72] & b[211])^(a[71] & b[212])^(a[70] & b[213])^(a[69] & b[214])^(a[68] & b[215])^(a[67] & b[216])^(a[66] & b[217])^(a[65] & b[218])^(a[64] & b[219])^(a[63] & b[220])^(a[62] & b[221])^(a[61] & b[222])^(a[60] & b[223])^(a[59] & b[224])^(a[58] & b[225])^(a[57] & b[226])^(a[56] & b[227])^(a[55] & b[228])^(a[54] & b[229])^(a[53] & b[230])^(a[52] & b[231])^(a[51] & b[232]);
assign y[284] = (a[232] & b[52])^(a[231] & b[53])^(a[230] & b[54])^(a[229] & b[55])^(a[228] & b[56])^(a[227] & b[57])^(a[226] & b[58])^(a[225] & b[59])^(a[224] & b[60])^(a[223] & b[61])^(a[222] & b[62])^(a[221] & b[63])^(a[220] & b[64])^(a[219] & b[65])^(a[218] & b[66])^(a[217] & b[67])^(a[216] & b[68])^(a[215] & b[69])^(a[214] & b[70])^(a[213] & b[71])^(a[212] & b[72])^(a[211] & b[73])^(a[210] & b[74])^(a[209] & b[75])^(a[208] & b[76])^(a[207] & b[77])^(a[206] & b[78])^(a[205] & b[79])^(a[204] & b[80])^(a[203] & b[81])^(a[202] & b[82])^(a[201] & b[83])^(a[200] & b[84])^(a[199] & b[85])^(a[198] & b[86])^(a[197] & b[87])^(a[196] & b[88])^(a[195] & b[89])^(a[194] & b[90])^(a[193] & b[91])^(a[192] & b[92])^(a[191] & b[93])^(a[190] & b[94])^(a[189] & b[95])^(a[188] & b[96])^(a[187] & b[97])^(a[186] & b[98])^(a[185] & b[99])^(a[184] & b[100])^(a[183] & b[101])^(a[182] & b[102])^(a[181] & b[103])^(a[180] & b[104])^(a[179] & b[105])^(a[178] & b[106])^(a[177] & b[107])^(a[176] & b[108])^(a[175] & b[109])^(a[174] & b[110])^(a[173] & b[111])^(a[172] & b[112])^(a[171] & b[113])^(a[170] & b[114])^(a[169] & b[115])^(a[168] & b[116])^(a[167] & b[117])^(a[166] & b[118])^(a[165] & b[119])^(a[164] & b[120])^(a[163] & b[121])^(a[162] & b[122])^(a[161] & b[123])^(a[160] & b[124])^(a[159] & b[125])^(a[158] & b[126])^(a[157] & b[127])^(a[156] & b[128])^(a[155] & b[129])^(a[154] & b[130])^(a[153] & b[131])^(a[152] & b[132])^(a[151] & b[133])^(a[150] & b[134])^(a[149] & b[135])^(a[148] & b[136])^(a[147] & b[137])^(a[146] & b[138])^(a[145] & b[139])^(a[144] & b[140])^(a[143] & b[141])^(a[142] & b[142])^(a[141] & b[143])^(a[140] & b[144])^(a[139] & b[145])^(a[138] & b[146])^(a[137] & b[147])^(a[136] & b[148])^(a[135] & b[149])^(a[134] & b[150])^(a[133] & b[151])^(a[132] & b[152])^(a[131] & b[153])^(a[130] & b[154])^(a[129] & b[155])^(a[128] & b[156])^(a[127] & b[157])^(a[126] & b[158])^(a[125] & b[159])^(a[124] & b[160])^(a[123] & b[161])^(a[122] & b[162])^(a[121] & b[163])^(a[120] & b[164])^(a[119] & b[165])^(a[118] & b[166])^(a[117] & b[167])^(a[116] & b[168])^(a[115] & b[169])^(a[114] & b[170])^(a[113] & b[171])^(a[112] & b[172])^(a[111] & b[173])^(a[110] & b[174])^(a[109] & b[175])^(a[108] & b[176])^(a[107] & b[177])^(a[106] & b[178])^(a[105] & b[179])^(a[104] & b[180])^(a[103] & b[181])^(a[102] & b[182])^(a[101] & b[183])^(a[100] & b[184])^(a[99] & b[185])^(a[98] & b[186])^(a[97] & b[187])^(a[96] & b[188])^(a[95] & b[189])^(a[94] & b[190])^(a[93] & b[191])^(a[92] & b[192])^(a[91] & b[193])^(a[90] & b[194])^(a[89] & b[195])^(a[88] & b[196])^(a[87] & b[197])^(a[86] & b[198])^(a[85] & b[199])^(a[84] & b[200])^(a[83] & b[201])^(a[82] & b[202])^(a[81] & b[203])^(a[80] & b[204])^(a[79] & b[205])^(a[78] & b[206])^(a[77] & b[207])^(a[76] & b[208])^(a[75] & b[209])^(a[74] & b[210])^(a[73] & b[211])^(a[72] & b[212])^(a[71] & b[213])^(a[70] & b[214])^(a[69] & b[215])^(a[68] & b[216])^(a[67] & b[217])^(a[66] & b[218])^(a[65] & b[219])^(a[64] & b[220])^(a[63] & b[221])^(a[62] & b[222])^(a[61] & b[223])^(a[60] & b[224])^(a[59] & b[225])^(a[58] & b[226])^(a[57] & b[227])^(a[56] & b[228])^(a[55] & b[229])^(a[54] & b[230])^(a[53] & b[231])^(a[52] & b[232]);
assign y[285] = (a[232] & b[53])^(a[231] & b[54])^(a[230] & b[55])^(a[229] & b[56])^(a[228] & b[57])^(a[227] & b[58])^(a[226] & b[59])^(a[225] & b[60])^(a[224] & b[61])^(a[223] & b[62])^(a[222] & b[63])^(a[221] & b[64])^(a[220] & b[65])^(a[219] & b[66])^(a[218] & b[67])^(a[217] & b[68])^(a[216] & b[69])^(a[215] & b[70])^(a[214] & b[71])^(a[213] & b[72])^(a[212] & b[73])^(a[211] & b[74])^(a[210] & b[75])^(a[209] & b[76])^(a[208] & b[77])^(a[207] & b[78])^(a[206] & b[79])^(a[205] & b[80])^(a[204] & b[81])^(a[203] & b[82])^(a[202] & b[83])^(a[201] & b[84])^(a[200] & b[85])^(a[199] & b[86])^(a[198] & b[87])^(a[197] & b[88])^(a[196] & b[89])^(a[195] & b[90])^(a[194] & b[91])^(a[193] & b[92])^(a[192] & b[93])^(a[191] & b[94])^(a[190] & b[95])^(a[189] & b[96])^(a[188] & b[97])^(a[187] & b[98])^(a[186] & b[99])^(a[185] & b[100])^(a[184] & b[101])^(a[183] & b[102])^(a[182] & b[103])^(a[181] & b[104])^(a[180] & b[105])^(a[179] & b[106])^(a[178] & b[107])^(a[177] & b[108])^(a[176] & b[109])^(a[175] & b[110])^(a[174] & b[111])^(a[173] & b[112])^(a[172] & b[113])^(a[171] & b[114])^(a[170] & b[115])^(a[169] & b[116])^(a[168] & b[117])^(a[167] & b[118])^(a[166] & b[119])^(a[165] & b[120])^(a[164] & b[121])^(a[163] & b[122])^(a[162] & b[123])^(a[161] & b[124])^(a[160] & b[125])^(a[159] & b[126])^(a[158] & b[127])^(a[157] & b[128])^(a[156] & b[129])^(a[155] & b[130])^(a[154] & b[131])^(a[153] & b[132])^(a[152] & b[133])^(a[151] & b[134])^(a[150] & b[135])^(a[149] & b[136])^(a[148] & b[137])^(a[147] & b[138])^(a[146] & b[139])^(a[145] & b[140])^(a[144] & b[141])^(a[143] & b[142])^(a[142] & b[143])^(a[141] & b[144])^(a[140] & b[145])^(a[139] & b[146])^(a[138] & b[147])^(a[137] & b[148])^(a[136] & b[149])^(a[135] & b[150])^(a[134] & b[151])^(a[133] & b[152])^(a[132] & b[153])^(a[131] & b[154])^(a[130] & b[155])^(a[129] & b[156])^(a[128] & b[157])^(a[127] & b[158])^(a[126] & b[159])^(a[125] & b[160])^(a[124] & b[161])^(a[123] & b[162])^(a[122] & b[163])^(a[121] & b[164])^(a[120] & b[165])^(a[119] & b[166])^(a[118] & b[167])^(a[117] & b[168])^(a[116] & b[169])^(a[115] & b[170])^(a[114] & b[171])^(a[113] & b[172])^(a[112] & b[173])^(a[111] & b[174])^(a[110] & b[175])^(a[109] & b[176])^(a[108] & b[177])^(a[107] & b[178])^(a[106] & b[179])^(a[105] & b[180])^(a[104] & b[181])^(a[103] & b[182])^(a[102] & b[183])^(a[101] & b[184])^(a[100] & b[185])^(a[99] & b[186])^(a[98] & b[187])^(a[97] & b[188])^(a[96] & b[189])^(a[95] & b[190])^(a[94] & b[191])^(a[93] & b[192])^(a[92] & b[193])^(a[91] & b[194])^(a[90] & b[195])^(a[89] & b[196])^(a[88] & b[197])^(a[87] & b[198])^(a[86] & b[199])^(a[85] & b[200])^(a[84] & b[201])^(a[83] & b[202])^(a[82] & b[203])^(a[81] & b[204])^(a[80] & b[205])^(a[79] & b[206])^(a[78] & b[207])^(a[77] & b[208])^(a[76] & b[209])^(a[75] & b[210])^(a[74] & b[211])^(a[73] & b[212])^(a[72] & b[213])^(a[71] & b[214])^(a[70] & b[215])^(a[69] & b[216])^(a[68] & b[217])^(a[67] & b[218])^(a[66] & b[219])^(a[65] & b[220])^(a[64] & b[221])^(a[63] & b[222])^(a[62] & b[223])^(a[61] & b[224])^(a[60] & b[225])^(a[59] & b[226])^(a[58] & b[227])^(a[57] & b[228])^(a[56] & b[229])^(a[55] & b[230])^(a[54] & b[231])^(a[53] & b[232]);
assign y[286] = (a[232] & b[54])^(a[231] & b[55])^(a[230] & b[56])^(a[229] & b[57])^(a[228] & b[58])^(a[227] & b[59])^(a[226] & b[60])^(a[225] & b[61])^(a[224] & b[62])^(a[223] & b[63])^(a[222] & b[64])^(a[221] & b[65])^(a[220] & b[66])^(a[219] & b[67])^(a[218] & b[68])^(a[217] & b[69])^(a[216] & b[70])^(a[215] & b[71])^(a[214] & b[72])^(a[213] & b[73])^(a[212] & b[74])^(a[211] & b[75])^(a[210] & b[76])^(a[209] & b[77])^(a[208] & b[78])^(a[207] & b[79])^(a[206] & b[80])^(a[205] & b[81])^(a[204] & b[82])^(a[203] & b[83])^(a[202] & b[84])^(a[201] & b[85])^(a[200] & b[86])^(a[199] & b[87])^(a[198] & b[88])^(a[197] & b[89])^(a[196] & b[90])^(a[195] & b[91])^(a[194] & b[92])^(a[193] & b[93])^(a[192] & b[94])^(a[191] & b[95])^(a[190] & b[96])^(a[189] & b[97])^(a[188] & b[98])^(a[187] & b[99])^(a[186] & b[100])^(a[185] & b[101])^(a[184] & b[102])^(a[183] & b[103])^(a[182] & b[104])^(a[181] & b[105])^(a[180] & b[106])^(a[179] & b[107])^(a[178] & b[108])^(a[177] & b[109])^(a[176] & b[110])^(a[175] & b[111])^(a[174] & b[112])^(a[173] & b[113])^(a[172] & b[114])^(a[171] & b[115])^(a[170] & b[116])^(a[169] & b[117])^(a[168] & b[118])^(a[167] & b[119])^(a[166] & b[120])^(a[165] & b[121])^(a[164] & b[122])^(a[163] & b[123])^(a[162] & b[124])^(a[161] & b[125])^(a[160] & b[126])^(a[159] & b[127])^(a[158] & b[128])^(a[157] & b[129])^(a[156] & b[130])^(a[155] & b[131])^(a[154] & b[132])^(a[153] & b[133])^(a[152] & b[134])^(a[151] & b[135])^(a[150] & b[136])^(a[149] & b[137])^(a[148] & b[138])^(a[147] & b[139])^(a[146] & b[140])^(a[145] & b[141])^(a[144] & b[142])^(a[143] & b[143])^(a[142] & b[144])^(a[141] & b[145])^(a[140] & b[146])^(a[139] & b[147])^(a[138] & b[148])^(a[137] & b[149])^(a[136] & b[150])^(a[135] & b[151])^(a[134] & b[152])^(a[133] & b[153])^(a[132] & b[154])^(a[131] & b[155])^(a[130] & b[156])^(a[129] & b[157])^(a[128] & b[158])^(a[127] & b[159])^(a[126] & b[160])^(a[125] & b[161])^(a[124] & b[162])^(a[123] & b[163])^(a[122] & b[164])^(a[121] & b[165])^(a[120] & b[166])^(a[119] & b[167])^(a[118] & b[168])^(a[117] & b[169])^(a[116] & b[170])^(a[115] & b[171])^(a[114] & b[172])^(a[113] & b[173])^(a[112] & b[174])^(a[111] & b[175])^(a[110] & b[176])^(a[109] & b[177])^(a[108] & b[178])^(a[107] & b[179])^(a[106] & b[180])^(a[105] & b[181])^(a[104] & b[182])^(a[103] & b[183])^(a[102] & b[184])^(a[101] & b[185])^(a[100] & b[186])^(a[99] & b[187])^(a[98] & b[188])^(a[97] & b[189])^(a[96] & b[190])^(a[95] & b[191])^(a[94] & b[192])^(a[93] & b[193])^(a[92] & b[194])^(a[91] & b[195])^(a[90] & b[196])^(a[89] & b[197])^(a[88] & b[198])^(a[87] & b[199])^(a[86] & b[200])^(a[85] & b[201])^(a[84] & b[202])^(a[83] & b[203])^(a[82] & b[204])^(a[81] & b[205])^(a[80] & b[206])^(a[79] & b[207])^(a[78] & b[208])^(a[77] & b[209])^(a[76] & b[210])^(a[75] & b[211])^(a[74] & b[212])^(a[73] & b[213])^(a[72] & b[214])^(a[71] & b[215])^(a[70] & b[216])^(a[69] & b[217])^(a[68] & b[218])^(a[67] & b[219])^(a[66] & b[220])^(a[65] & b[221])^(a[64] & b[222])^(a[63] & b[223])^(a[62] & b[224])^(a[61] & b[225])^(a[60] & b[226])^(a[59] & b[227])^(a[58] & b[228])^(a[57] & b[229])^(a[56] & b[230])^(a[55] & b[231])^(a[54] & b[232]);
assign y[287] = (a[232] & b[55])^(a[231] & b[56])^(a[230] & b[57])^(a[229] & b[58])^(a[228] & b[59])^(a[227] & b[60])^(a[226] & b[61])^(a[225] & b[62])^(a[224] & b[63])^(a[223] & b[64])^(a[222] & b[65])^(a[221] & b[66])^(a[220] & b[67])^(a[219] & b[68])^(a[218] & b[69])^(a[217] & b[70])^(a[216] & b[71])^(a[215] & b[72])^(a[214] & b[73])^(a[213] & b[74])^(a[212] & b[75])^(a[211] & b[76])^(a[210] & b[77])^(a[209] & b[78])^(a[208] & b[79])^(a[207] & b[80])^(a[206] & b[81])^(a[205] & b[82])^(a[204] & b[83])^(a[203] & b[84])^(a[202] & b[85])^(a[201] & b[86])^(a[200] & b[87])^(a[199] & b[88])^(a[198] & b[89])^(a[197] & b[90])^(a[196] & b[91])^(a[195] & b[92])^(a[194] & b[93])^(a[193] & b[94])^(a[192] & b[95])^(a[191] & b[96])^(a[190] & b[97])^(a[189] & b[98])^(a[188] & b[99])^(a[187] & b[100])^(a[186] & b[101])^(a[185] & b[102])^(a[184] & b[103])^(a[183] & b[104])^(a[182] & b[105])^(a[181] & b[106])^(a[180] & b[107])^(a[179] & b[108])^(a[178] & b[109])^(a[177] & b[110])^(a[176] & b[111])^(a[175] & b[112])^(a[174] & b[113])^(a[173] & b[114])^(a[172] & b[115])^(a[171] & b[116])^(a[170] & b[117])^(a[169] & b[118])^(a[168] & b[119])^(a[167] & b[120])^(a[166] & b[121])^(a[165] & b[122])^(a[164] & b[123])^(a[163] & b[124])^(a[162] & b[125])^(a[161] & b[126])^(a[160] & b[127])^(a[159] & b[128])^(a[158] & b[129])^(a[157] & b[130])^(a[156] & b[131])^(a[155] & b[132])^(a[154] & b[133])^(a[153] & b[134])^(a[152] & b[135])^(a[151] & b[136])^(a[150] & b[137])^(a[149] & b[138])^(a[148] & b[139])^(a[147] & b[140])^(a[146] & b[141])^(a[145] & b[142])^(a[144] & b[143])^(a[143] & b[144])^(a[142] & b[145])^(a[141] & b[146])^(a[140] & b[147])^(a[139] & b[148])^(a[138] & b[149])^(a[137] & b[150])^(a[136] & b[151])^(a[135] & b[152])^(a[134] & b[153])^(a[133] & b[154])^(a[132] & b[155])^(a[131] & b[156])^(a[130] & b[157])^(a[129] & b[158])^(a[128] & b[159])^(a[127] & b[160])^(a[126] & b[161])^(a[125] & b[162])^(a[124] & b[163])^(a[123] & b[164])^(a[122] & b[165])^(a[121] & b[166])^(a[120] & b[167])^(a[119] & b[168])^(a[118] & b[169])^(a[117] & b[170])^(a[116] & b[171])^(a[115] & b[172])^(a[114] & b[173])^(a[113] & b[174])^(a[112] & b[175])^(a[111] & b[176])^(a[110] & b[177])^(a[109] & b[178])^(a[108] & b[179])^(a[107] & b[180])^(a[106] & b[181])^(a[105] & b[182])^(a[104] & b[183])^(a[103] & b[184])^(a[102] & b[185])^(a[101] & b[186])^(a[100] & b[187])^(a[99] & b[188])^(a[98] & b[189])^(a[97] & b[190])^(a[96] & b[191])^(a[95] & b[192])^(a[94] & b[193])^(a[93] & b[194])^(a[92] & b[195])^(a[91] & b[196])^(a[90] & b[197])^(a[89] & b[198])^(a[88] & b[199])^(a[87] & b[200])^(a[86] & b[201])^(a[85] & b[202])^(a[84] & b[203])^(a[83] & b[204])^(a[82] & b[205])^(a[81] & b[206])^(a[80] & b[207])^(a[79] & b[208])^(a[78] & b[209])^(a[77] & b[210])^(a[76] & b[211])^(a[75] & b[212])^(a[74] & b[213])^(a[73] & b[214])^(a[72] & b[215])^(a[71] & b[216])^(a[70] & b[217])^(a[69] & b[218])^(a[68] & b[219])^(a[67] & b[220])^(a[66] & b[221])^(a[65] & b[222])^(a[64] & b[223])^(a[63] & b[224])^(a[62] & b[225])^(a[61] & b[226])^(a[60] & b[227])^(a[59] & b[228])^(a[58] & b[229])^(a[57] & b[230])^(a[56] & b[231])^(a[55] & b[232]);
assign y[288] = (a[232] & b[56])^(a[231] & b[57])^(a[230] & b[58])^(a[229] & b[59])^(a[228] & b[60])^(a[227] & b[61])^(a[226] & b[62])^(a[225] & b[63])^(a[224] & b[64])^(a[223] & b[65])^(a[222] & b[66])^(a[221] & b[67])^(a[220] & b[68])^(a[219] & b[69])^(a[218] & b[70])^(a[217] & b[71])^(a[216] & b[72])^(a[215] & b[73])^(a[214] & b[74])^(a[213] & b[75])^(a[212] & b[76])^(a[211] & b[77])^(a[210] & b[78])^(a[209] & b[79])^(a[208] & b[80])^(a[207] & b[81])^(a[206] & b[82])^(a[205] & b[83])^(a[204] & b[84])^(a[203] & b[85])^(a[202] & b[86])^(a[201] & b[87])^(a[200] & b[88])^(a[199] & b[89])^(a[198] & b[90])^(a[197] & b[91])^(a[196] & b[92])^(a[195] & b[93])^(a[194] & b[94])^(a[193] & b[95])^(a[192] & b[96])^(a[191] & b[97])^(a[190] & b[98])^(a[189] & b[99])^(a[188] & b[100])^(a[187] & b[101])^(a[186] & b[102])^(a[185] & b[103])^(a[184] & b[104])^(a[183] & b[105])^(a[182] & b[106])^(a[181] & b[107])^(a[180] & b[108])^(a[179] & b[109])^(a[178] & b[110])^(a[177] & b[111])^(a[176] & b[112])^(a[175] & b[113])^(a[174] & b[114])^(a[173] & b[115])^(a[172] & b[116])^(a[171] & b[117])^(a[170] & b[118])^(a[169] & b[119])^(a[168] & b[120])^(a[167] & b[121])^(a[166] & b[122])^(a[165] & b[123])^(a[164] & b[124])^(a[163] & b[125])^(a[162] & b[126])^(a[161] & b[127])^(a[160] & b[128])^(a[159] & b[129])^(a[158] & b[130])^(a[157] & b[131])^(a[156] & b[132])^(a[155] & b[133])^(a[154] & b[134])^(a[153] & b[135])^(a[152] & b[136])^(a[151] & b[137])^(a[150] & b[138])^(a[149] & b[139])^(a[148] & b[140])^(a[147] & b[141])^(a[146] & b[142])^(a[145] & b[143])^(a[144] & b[144])^(a[143] & b[145])^(a[142] & b[146])^(a[141] & b[147])^(a[140] & b[148])^(a[139] & b[149])^(a[138] & b[150])^(a[137] & b[151])^(a[136] & b[152])^(a[135] & b[153])^(a[134] & b[154])^(a[133] & b[155])^(a[132] & b[156])^(a[131] & b[157])^(a[130] & b[158])^(a[129] & b[159])^(a[128] & b[160])^(a[127] & b[161])^(a[126] & b[162])^(a[125] & b[163])^(a[124] & b[164])^(a[123] & b[165])^(a[122] & b[166])^(a[121] & b[167])^(a[120] & b[168])^(a[119] & b[169])^(a[118] & b[170])^(a[117] & b[171])^(a[116] & b[172])^(a[115] & b[173])^(a[114] & b[174])^(a[113] & b[175])^(a[112] & b[176])^(a[111] & b[177])^(a[110] & b[178])^(a[109] & b[179])^(a[108] & b[180])^(a[107] & b[181])^(a[106] & b[182])^(a[105] & b[183])^(a[104] & b[184])^(a[103] & b[185])^(a[102] & b[186])^(a[101] & b[187])^(a[100] & b[188])^(a[99] & b[189])^(a[98] & b[190])^(a[97] & b[191])^(a[96] & b[192])^(a[95] & b[193])^(a[94] & b[194])^(a[93] & b[195])^(a[92] & b[196])^(a[91] & b[197])^(a[90] & b[198])^(a[89] & b[199])^(a[88] & b[200])^(a[87] & b[201])^(a[86] & b[202])^(a[85] & b[203])^(a[84] & b[204])^(a[83] & b[205])^(a[82] & b[206])^(a[81] & b[207])^(a[80] & b[208])^(a[79] & b[209])^(a[78] & b[210])^(a[77] & b[211])^(a[76] & b[212])^(a[75] & b[213])^(a[74] & b[214])^(a[73] & b[215])^(a[72] & b[216])^(a[71] & b[217])^(a[70] & b[218])^(a[69] & b[219])^(a[68] & b[220])^(a[67] & b[221])^(a[66] & b[222])^(a[65] & b[223])^(a[64] & b[224])^(a[63] & b[225])^(a[62] & b[226])^(a[61] & b[227])^(a[60] & b[228])^(a[59] & b[229])^(a[58] & b[230])^(a[57] & b[231])^(a[56] & b[232]);
assign y[289] = (a[232] & b[57])^(a[231] & b[58])^(a[230] & b[59])^(a[229] & b[60])^(a[228] & b[61])^(a[227] & b[62])^(a[226] & b[63])^(a[225] & b[64])^(a[224] & b[65])^(a[223] & b[66])^(a[222] & b[67])^(a[221] & b[68])^(a[220] & b[69])^(a[219] & b[70])^(a[218] & b[71])^(a[217] & b[72])^(a[216] & b[73])^(a[215] & b[74])^(a[214] & b[75])^(a[213] & b[76])^(a[212] & b[77])^(a[211] & b[78])^(a[210] & b[79])^(a[209] & b[80])^(a[208] & b[81])^(a[207] & b[82])^(a[206] & b[83])^(a[205] & b[84])^(a[204] & b[85])^(a[203] & b[86])^(a[202] & b[87])^(a[201] & b[88])^(a[200] & b[89])^(a[199] & b[90])^(a[198] & b[91])^(a[197] & b[92])^(a[196] & b[93])^(a[195] & b[94])^(a[194] & b[95])^(a[193] & b[96])^(a[192] & b[97])^(a[191] & b[98])^(a[190] & b[99])^(a[189] & b[100])^(a[188] & b[101])^(a[187] & b[102])^(a[186] & b[103])^(a[185] & b[104])^(a[184] & b[105])^(a[183] & b[106])^(a[182] & b[107])^(a[181] & b[108])^(a[180] & b[109])^(a[179] & b[110])^(a[178] & b[111])^(a[177] & b[112])^(a[176] & b[113])^(a[175] & b[114])^(a[174] & b[115])^(a[173] & b[116])^(a[172] & b[117])^(a[171] & b[118])^(a[170] & b[119])^(a[169] & b[120])^(a[168] & b[121])^(a[167] & b[122])^(a[166] & b[123])^(a[165] & b[124])^(a[164] & b[125])^(a[163] & b[126])^(a[162] & b[127])^(a[161] & b[128])^(a[160] & b[129])^(a[159] & b[130])^(a[158] & b[131])^(a[157] & b[132])^(a[156] & b[133])^(a[155] & b[134])^(a[154] & b[135])^(a[153] & b[136])^(a[152] & b[137])^(a[151] & b[138])^(a[150] & b[139])^(a[149] & b[140])^(a[148] & b[141])^(a[147] & b[142])^(a[146] & b[143])^(a[145] & b[144])^(a[144] & b[145])^(a[143] & b[146])^(a[142] & b[147])^(a[141] & b[148])^(a[140] & b[149])^(a[139] & b[150])^(a[138] & b[151])^(a[137] & b[152])^(a[136] & b[153])^(a[135] & b[154])^(a[134] & b[155])^(a[133] & b[156])^(a[132] & b[157])^(a[131] & b[158])^(a[130] & b[159])^(a[129] & b[160])^(a[128] & b[161])^(a[127] & b[162])^(a[126] & b[163])^(a[125] & b[164])^(a[124] & b[165])^(a[123] & b[166])^(a[122] & b[167])^(a[121] & b[168])^(a[120] & b[169])^(a[119] & b[170])^(a[118] & b[171])^(a[117] & b[172])^(a[116] & b[173])^(a[115] & b[174])^(a[114] & b[175])^(a[113] & b[176])^(a[112] & b[177])^(a[111] & b[178])^(a[110] & b[179])^(a[109] & b[180])^(a[108] & b[181])^(a[107] & b[182])^(a[106] & b[183])^(a[105] & b[184])^(a[104] & b[185])^(a[103] & b[186])^(a[102] & b[187])^(a[101] & b[188])^(a[100] & b[189])^(a[99] & b[190])^(a[98] & b[191])^(a[97] & b[192])^(a[96] & b[193])^(a[95] & b[194])^(a[94] & b[195])^(a[93] & b[196])^(a[92] & b[197])^(a[91] & b[198])^(a[90] & b[199])^(a[89] & b[200])^(a[88] & b[201])^(a[87] & b[202])^(a[86] & b[203])^(a[85] & b[204])^(a[84] & b[205])^(a[83] & b[206])^(a[82] & b[207])^(a[81] & b[208])^(a[80] & b[209])^(a[79] & b[210])^(a[78] & b[211])^(a[77] & b[212])^(a[76] & b[213])^(a[75] & b[214])^(a[74] & b[215])^(a[73] & b[216])^(a[72] & b[217])^(a[71] & b[218])^(a[70] & b[219])^(a[69] & b[220])^(a[68] & b[221])^(a[67] & b[222])^(a[66] & b[223])^(a[65] & b[224])^(a[64] & b[225])^(a[63] & b[226])^(a[62] & b[227])^(a[61] & b[228])^(a[60] & b[229])^(a[59] & b[230])^(a[58] & b[231])^(a[57] & b[232]);
assign y[290] = (a[232] & b[58])^(a[231] & b[59])^(a[230] & b[60])^(a[229] & b[61])^(a[228] & b[62])^(a[227] & b[63])^(a[226] & b[64])^(a[225] & b[65])^(a[224] & b[66])^(a[223] & b[67])^(a[222] & b[68])^(a[221] & b[69])^(a[220] & b[70])^(a[219] & b[71])^(a[218] & b[72])^(a[217] & b[73])^(a[216] & b[74])^(a[215] & b[75])^(a[214] & b[76])^(a[213] & b[77])^(a[212] & b[78])^(a[211] & b[79])^(a[210] & b[80])^(a[209] & b[81])^(a[208] & b[82])^(a[207] & b[83])^(a[206] & b[84])^(a[205] & b[85])^(a[204] & b[86])^(a[203] & b[87])^(a[202] & b[88])^(a[201] & b[89])^(a[200] & b[90])^(a[199] & b[91])^(a[198] & b[92])^(a[197] & b[93])^(a[196] & b[94])^(a[195] & b[95])^(a[194] & b[96])^(a[193] & b[97])^(a[192] & b[98])^(a[191] & b[99])^(a[190] & b[100])^(a[189] & b[101])^(a[188] & b[102])^(a[187] & b[103])^(a[186] & b[104])^(a[185] & b[105])^(a[184] & b[106])^(a[183] & b[107])^(a[182] & b[108])^(a[181] & b[109])^(a[180] & b[110])^(a[179] & b[111])^(a[178] & b[112])^(a[177] & b[113])^(a[176] & b[114])^(a[175] & b[115])^(a[174] & b[116])^(a[173] & b[117])^(a[172] & b[118])^(a[171] & b[119])^(a[170] & b[120])^(a[169] & b[121])^(a[168] & b[122])^(a[167] & b[123])^(a[166] & b[124])^(a[165] & b[125])^(a[164] & b[126])^(a[163] & b[127])^(a[162] & b[128])^(a[161] & b[129])^(a[160] & b[130])^(a[159] & b[131])^(a[158] & b[132])^(a[157] & b[133])^(a[156] & b[134])^(a[155] & b[135])^(a[154] & b[136])^(a[153] & b[137])^(a[152] & b[138])^(a[151] & b[139])^(a[150] & b[140])^(a[149] & b[141])^(a[148] & b[142])^(a[147] & b[143])^(a[146] & b[144])^(a[145] & b[145])^(a[144] & b[146])^(a[143] & b[147])^(a[142] & b[148])^(a[141] & b[149])^(a[140] & b[150])^(a[139] & b[151])^(a[138] & b[152])^(a[137] & b[153])^(a[136] & b[154])^(a[135] & b[155])^(a[134] & b[156])^(a[133] & b[157])^(a[132] & b[158])^(a[131] & b[159])^(a[130] & b[160])^(a[129] & b[161])^(a[128] & b[162])^(a[127] & b[163])^(a[126] & b[164])^(a[125] & b[165])^(a[124] & b[166])^(a[123] & b[167])^(a[122] & b[168])^(a[121] & b[169])^(a[120] & b[170])^(a[119] & b[171])^(a[118] & b[172])^(a[117] & b[173])^(a[116] & b[174])^(a[115] & b[175])^(a[114] & b[176])^(a[113] & b[177])^(a[112] & b[178])^(a[111] & b[179])^(a[110] & b[180])^(a[109] & b[181])^(a[108] & b[182])^(a[107] & b[183])^(a[106] & b[184])^(a[105] & b[185])^(a[104] & b[186])^(a[103] & b[187])^(a[102] & b[188])^(a[101] & b[189])^(a[100] & b[190])^(a[99] & b[191])^(a[98] & b[192])^(a[97] & b[193])^(a[96] & b[194])^(a[95] & b[195])^(a[94] & b[196])^(a[93] & b[197])^(a[92] & b[198])^(a[91] & b[199])^(a[90] & b[200])^(a[89] & b[201])^(a[88] & b[202])^(a[87] & b[203])^(a[86] & b[204])^(a[85] & b[205])^(a[84] & b[206])^(a[83] & b[207])^(a[82] & b[208])^(a[81] & b[209])^(a[80] & b[210])^(a[79] & b[211])^(a[78] & b[212])^(a[77] & b[213])^(a[76] & b[214])^(a[75] & b[215])^(a[74] & b[216])^(a[73] & b[217])^(a[72] & b[218])^(a[71] & b[219])^(a[70] & b[220])^(a[69] & b[221])^(a[68] & b[222])^(a[67] & b[223])^(a[66] & b[224])^(a[65] & b[225])^(a[64] & b[226])^(a[63] & b[227])^(a[62] & b[228])^(a[61] & b[229])^(a[60] & b[230])^(a[59] & b[231])^(a[58] & b[232]);
assign y[291] = (a[232] & b[59])^(a[231] & b[60])^(a[230] & b[61])^(a[229] & b[62])^(a[228] & b[63])^(a[227] & b[64])^(a[226] & b[65])^(a[225] & b[66])^(a[224] & b[67])^(a[223] & b[68])^(a[222] & b[69])^(a[221] & b[70])^(a[220] & b[71])^(a[219] & b[72])^(a[218] & b[73])^(a[217] & b[74])^(a[216] & b[75])^(a[215] & b[76])^(a[214] & b[77])^(a[213] & b[78])^(a[212] & b[79])^(a[211] & b[80])^(a[210] & b[81])^(a[209] & b[82])^(a[208] & b[83])^(a[207] & b[84])^(a[206] & b[85])^(a[205] & b[86])^(a[204] & b[87])^(a[203] & b[88])^(a[202] & b[89])^(a[201] & b[90])^(a[200] & b[91])^(a[199] & b[92])^(a[198] & b[93])^(a[197] & b[94])^(a[196] & b[95])^(a[195] & b[96])^(a[194] & b[97])^(a[193] & b[98])^(a[192] & b[99])^(a[191] & b[100])^(a[190] & b[101])^(a[189] & b[102])^(a[188] & b[103])^(a[187] & b[104])^(a[186] & b[105])^(a[185] & b[106])^(a[184] & b[107])^(a[183] & b[108])^(a[182] & b[109])^(a[181] & b[110])^(a[180] & b[111])^(a[179] & b[112])^(a[178] & b[113])^(a[177] & b[114])^(a[176] & b[115])^(a[175] & b[116])^(a[174] & b[117])^(a[173] & b[118])^(a[172] & b[119])^(a[171] & b[120])^(a[170] & b[121])^(a[169] & b[122])^(a[168] & b[123])^(a[167] & b[124])^(a[166] & b[125])^(a[165] & b[126])^(a[164] & b[127])^(a[163] & b[128])^(a[162] & b[129])^(a[161] & b[130])^(a[160] & b[131])^(a[159] & b[132])^(a[158] & b[133])^(a[157] & b[134])^(a[156] & b[135])^(a[155] & b[136])^(a[154] & b[137])^(a[153] & b[138])^(a[152] & b[139])^(a[151] & b[140])^(a[150] & b[141])^(a[149] & b[142])^(a[148] & b[143])^(a[147] & b[144])^(a[146] & b[145])^(a[145] & b[146])^(a[144] & b[147])^(a[143] & b[148])^(a[142] & b[149])^(a[141] & b[150])^(a[140] & b[151])^(a[139] & b[152])^(a[138] & b[153])^(a[137] & b[154])^(a[136] & b[155])^(a[135] & b[156])^(a[134] & b[157])^(a[133] & b[158])^(a[132] & b[159])^(a[131] & b[160])^(a[130] & b[161])^(a[129] & b[162])^(a[128] & b[163])^(a[127] & b[164])^(a[126] & b[165])^(a[125] & b[166])^(a[124] & b[167])^(a[123] & b[168])^(a[122] & b[169])^(a[121] & b[170])^(a[120] & b[171])^(a[119] & b[172])^(a[118] & b[173])^(a[117] & b[174])^(a[116] & b[175])^(a[115] & b[176])^(a[114] & b[177])^(a[113] & b[178])^(a[112] & b[179])^(a[111] & b[180])^(a[110] & b[181])^(a[109] & b[182])^(a[108] & b[183])^(a[107] & b[184])^(a[106] & b[185])^(a[105] & b[186])^(a[104] & b[187])^(a[103] & b[188])^(a[102] & b[189])^(a[101] & b[190])^(a[100] & b[191])^(a[99] & b[192])^(a[98] & b[193])^(a[97] & b[194])^(a[96] & b[195])^(a[95] & b[196])^(a[94] & b[197])^(a[93] & b[198])^(a[92] & b[199])^(a[91] & b[200])^(a[90] & b[201])^(a[89] & b[202])^(a[88] & b[203])^(a[87] & b[204])^(a[86] & b[205])^(a[85] & b[206])^(a[84] & b[207])^(a[83] & b[208])^(a[82] & b[209])^(a[81] & b[210])^(a[80] & b[211])^(a[79] & b[212])^(a[78] & b[213])^(a[77] & b[214])^(a[76] & b[215])^(a[75] & b[216])^(a[74] & b[217])^(a[73] & b[218])^(a[72] & b[219])^(a[71] & b[220])^(a[70] & b[221])^(a[69] & b[222])^(a[68] & b[223])^(a[67] & b[224])^(a[66] & b[225])^(a[65] & b[226])^(a[64] & b[227])^(a[63] & b[228])^(a[62] & b[229])^(a[61] & b[230])^(a[60] & b[231])^(a[59] & b[232]);
assign y[292] = (a[232] & b[60])^(a[231] & b[61])^(a[230] & b[62])^(a[229] & b[63])^(a[228] & b[64])^(a[227] & b[65])^(a[226] & b[66])^(a[225] & b[67])^(a[224] & b[68])^(a[223] & b[69])^(a[222] & b[70])^(a[221] & b[71])^(a[220] & b[72])^(a[219] & b[73])^(a[218] & b[74])^(a[217] & b[75])^(a[216] & b[76])^(a[215] & b[77])^(a[214] & b[78])^(a[213] & b[79])^(a[212] & b[80])^(a[211] & b[81])^(a[210] & b[82])^(a[209] & b[83])^(a[208] & b[84])^(a[207] & b[85])^(a[206] & b[86])^(a[205] & b[87])^(a[204] & b[88])^(a[203] & b[89])^(a[202] & b[90])^(a[201] & b[91])^(a[200] & b[92])^(a[199] & b[93])^(a[198] & b[94])^(a[197] & b[95])^(a[196] & b[96])^(a[195] & b[97])^(a[194] & b[98])^(a[193] & b[99])^(a[192] & b[100])^(a[191] & b[101])^(a[190] & b[102])^(a[189] & b[103])^(a[188] & b[104])^(a[187] & b[105])^(a[186] & b[106])^(a[185] & b[107])^(a[184] & b[108])^(a[183] & b[109])^(a[182] & b[110])^(a[181] & b[111])^(a[180] & b[112])^(a[179] & b[113])^(a[178] & b[114])^(a[177] & b[115])^(a[176] & b[116])^(a[175] & b[117])^(a[174] & b[118])^(a[173] & b[119])^(a[172] & b[120])^(a[171] & b[121])^(a[170] & b[122])^(a[169] & b[123])^(a[168] & b[124])^(a[167] & b[125])^(a[166] & b[126])^(a[165] & b[127])^(a[164] & b[128])^(a[163] & b[129])^(a[162] & b[130])^(a[161] & b[131])^(a[160] & b[132])^(a[159] & b[133])^(a[158] & b[134])^(a[157] & b[135])^(a[156] & b[136])^(a[155] & b[137])^(a[154] & b[138])^(a[153] & b[139])^(a[152] & b[140])^(a[151] & b[141])^(a[150] & b[142])^(a[149] & b[143])^(a[148] & b[144])^(a[147] & b[145])^(a[146] & b[146])^(a[145] & b[147])^(a[144] & b[148])^(a[143] & b[149])^(a[142] & b[150])^(a[141] & b[151])^(a[140] & b[152])^(a[139] & b[153])^(a[138] & b[154])^(a[137] & b[155])^(a[136] & b[156])^(a[135] & b[157])^(a[134] & b[158])^(a[133] & b[159])^(a[132] & b[160])^(a[131] & b[161])^(a[130] & b[162])^(a[129] & b[163])^(a[128] & b[164])^(a[127] & b[165])^(a[126] & b[166])^(a[125] & b[167])^(a[124] & b[168])^(a[123] & b[169])^(a[122] & b[170])^(a[121] & b[171])^(a[120] & b[172])^(a[119] & b[173])^(a[118] & b[174])^(a[117] & b[175])^(a[116] & b[176])^(a[115] & b[177])^(a[114] & b[178])^(a[113] & b[179])^(a[112] & b[180])^(a[111] & b[181])^(a[110] & b[182])^(a[109] & b[183])^(a[108] & b[184])^(a[107] & b[185])^(a[106] & b[186])^(a[105] & b[187])^(a[104] & b[188])^(a[103] & b[189])^(a[102] & b[190])^(a[101] & b[191])^(a[100] & b[192])^(a[99] & b[193])^(a[98] & b[194])^(a[97] & b[195])^(a[96] & b[196])^(a[95] & b[197])^(a[94] & b[198])^(a[93] & b[199])^(a[92] & b[200])^(a[91] & b[201])^(a[90] & b[202])^(a[89] & b[203])^(a[88] & b[204])^(a[87] & b[205])^(a[86] & b[206])^(a[85] & b[207])^(a[84] & b[208])^(a[83] & b[209])^(a[82] & b[210])^(a[81] & b[211])^(a[80] & b[212])^(a[79] & b[213])^(a[78] & b[214])^(a[77] & b[215])^(a[76] & b[216])^(a[75] & b[217])^(a[74] & b[218])^(a[73] & b[219])^(a[72] & b[220])^(a[71] & b[221])^(a[70] & b[222])^(a[69] & b[223])^(a[68] & b[224])^(a[67] & b[225])^(a[66] & b[226])^(a[65] & b[227])^(a[64] & b[228])^(a[63] & b[229])^(a[62] & b[230])^(a[61] & b[231])^(a[60] & b[232]);
assign y[293] = (a[232] & b[61])^(a[231] & b[62])^(a[230] & b[63])^(a[229] & b[64])^(a[228] & b[65])^(a[227] & b[66])^(a[226] & b[67])^(a[225] & b[68])^(a[224] & b[69])^(a[223] & b[70])^(a[222] & b[71])^(a[221] & b[72])^(a[220] & b[73])^(a[219] & b[74])^(a[218] & b[75])^(a[217] & b[76])^(a[216] & b[77])^(a[215] & b[78])^(a[214] & b[79])^(a[213] & b[80])^(a[212] & b[81])^(a[211] & b[82])^(a[210] & b[83])^(a[209] & b[84])^(a[208] & b[85])^(a[207] & b[86])^(a[206] & b[87])^(a[205] & b[88])^(a[204] & b[89])^(a[203] & b[90])^(a[202] & b[91])^(a[201] & b[92])^(a[200] & b[93])^(a[199] & b[94])^(a[198] & b[95])^(a[197] & b[96])^(a[196] & b[97])^(a[195] & b[98])^(a[194] & b[99])^(a[193] & b[100])^(a[192] & b[101])^(a[191] & b[102])^(a[190] & b[103])^(a[189] & b[104])^(a[188] & b[105])^(a[187] & b[106])^(a[186] & b[107])^(a[185] & b[108])^(a[184] & b[109])^(a[183] & b[110])^(a[182] & b[111])^(a[181] & b[112])^(a[180] & b[113])^(a[179] & b[114])^(a[178] & b[115])^(a[177] & b[116])^(a[176] & b[117])^(a[175] & b[118])^(a[174] & b[119])^(a[173] & b[120])^(a[172] & b[121])^(a[171] & b[122])^(a[170] & b[123])^(a[169] & b[124])^(a[168] & b[125])^(a[167] & b[126])^(a[166] & b[127])^(a[165] & b[128])^(a[164] & b[129])^(a[163] & b[130])^(a[162] & b[131])^(a[161] & b[132])^(a[160] & b[133])^(a[159] & b[134])^(a[158] & b[135])^(a[157] & b[136])^(a[156] & b[137])^(a[155] & b[138])^(a[154] & b[139])^(a[153] & b[140])^(a[152] & b[141])^(a[151] & b[142])^(a[150] & b[143])^(a[149] & b[144])^(a[148] & b[145])^(a[147] & b[146])^(a[146] & b[147])^(a[145] & b[148])^(a[144] & b[149])^(a[143] & b[150])^(a[142] & b[151])^(a[141] & b[152])^(a[140] & b[153])^(a[139] & b[154])^(a[138] & b[155])^(a[137] & b[156])^(a[136] & b[157])^(a[135] & b[158])^(a[134] & b[159])^(a[133] & b[160])^(a[132] & b[161])^(a[131] & b[162])^(a[130] & b[163])^(a[129] & b[164])^(a[128] & b[165])^(a[127] & b[166])^(a[126] & b[167])^(a[125] & b[168])^(a[124] & b[169])^(a[123] & b[170])^(a[122] & b[171])^(a[121] & b[172])^(a[120] & b[173])^(a[119] & b[174])^(a[118] & b[175])^(a[117] & b[176])^(a[116] & b[177])^(a[115] & b[178])^(a[114] & b[179])^(a[113] & b[180])^(a[112] & b[181])^(a[111] & b[182])^(a[110] & b[183])^(a[109] & b[184])^(a[108] & b[185])^(a[107] & b[186])^(a[106] & b[187])^(a[105] & b[188])^(a[104] & b[189])^(a[103] & b[190])^(a[102] & b[191])^(a[101] & b[192])^(a[100] & b[193])^(a[99] & b[194])^(a[98] & b[195])^(a[97] & b[196])^(a[96] & b[197])^(a[95] & b[198])^(a[94] & b[199])^(a[93] & b[200])^(a[92] & b[201])^(a[91] & b[202])^(a[90] & b[203])^(a[89] & b[204])^(a[88] & b[205])^(a[87] & b[206])^(a[86] & b[207])^(a[85] & b[208])^(a[84] & b[209])^(a[83] & b[210])^(a[82] & b[211])^(a[81] & b[212])^(a[80] & b[213])^(a[79] & b[214])^(a[78] & b[215])^(a[77] & b[216])^(a[76] & b[217])^(a[75] & b[218])^(a[74] & b[219])^(a[73] & b[220])^(a[72] & b[221])^(a[71] & b[222])^(a[70] & b[223])^(a[69] & b[224])^(a[68] & b[225])^(a[67] & b[226])^(a[66] & b[227])^(a[65] & b[228])^(a[64] & b[229])^(a[63] & b[230])^(a[62] & b[231])^(a[61] & b[232]);
assign y[294] = (a[232] & b[62])^(a[231] & b[63])^(a[230] & b[64])^(a[229] & b[65])^(a[228] & b[66])^(a[227] & b[67])^(a[226] & b[68])^(a[225] & b[69])^(a[224] & b[70])^(a[223] & b[71])^(a[222] & b[72])^(a[221] & b[73])^(a[220] & b[74])^(a[219] & b[75])^(a[218] & b[76])^(a[217] & b[77])^(a[216] & b[78])^(a[215] & b[79])^(a[214] & b[80])^(a[213] & b[81])^(a[212] & b[82])^(a[211] & b[83])^(a[210] & b[84])^(a[209] & b[85])^(a[208] & b[86])^(a[207] & b[87])^(a[206] & b[88])^(a[205] & b[89])^(a[204] & b[90])^(a[203] & b[91])^(a[202] & b[92])^(a[201] & b[93])^(a[200] & b[94])^(a[199] & b[95])^(a[198] & b[96])^(a[197] & b[97])^(a[196] & b[98])^(a[195] & b[99])^(a[194] & b[100])^(a[193] & b[101])^(a[192] & b[102])^(a[191] & b[103])^(a[190] & b[104])^(a[189] & b[105])^(a[188] & b[106])^(a[187] & b[107])^(a[186] & b[108])^(a[185] & b[109])^(a[184] & b[110])^(a[183] & b[111])^(a[182] & b[112])^(a[181] & b[113])^(a[180] & b[114])^(a[179] & b[115])^(a[178] & b[116])^(a[177] & b[117])^(a[176] & b[118])^(a[175] & b[119])^(a[174] & b[120])^(a[173] & b[121])^(a[172] & b[122])^(a[171] & b[123])^(a[170] & b[124])^(a[169] & b[125])^(a[168] & b[126])^(a[167] & b[127])^(a[166] & b[128])^(a[165] & b[129])^(a[164] & b[130])^(a[163] & b[131])^(a[162] & b[132])^(a[161] & b[133])^(a[160] & b[134])^(a[159] & b[135])^(a[158] & b[136])^(a[157] & b[137])^(a[156] & b[138])^(a[155] & b[139])^(a[154] & b[140])^(a[153] & b[141])^(a[152] & b[142])^(a[151] & b[143])^(a[150] & b[144])^(a[149] & b[145])^(a[148] & b[146])^(a[147] & b[147])^(a[146] & b[148])^(a[145] & b[149])^(a[144] & b[150])^(a[143] & b[151])^(a[142] & b[152])^(a[141] & b[153])^(a[140] & b[154])^(a[139] & b[155])^(a[138] & b[156])^(a[137] & b[157])^(a[136] & b[158])^(a[135] & b[159])^(a[134] & b[160])^(a[133] & b[161])^(a[132] & b[162])^(a[131] & b[163])^(a[130] & b[164])^(a[129] & b[165])^(a[128] & b[166])^(a[127] & b[167])^(a[126] & b[168])^(a[125] & b[169])^(a[124] & b[170])^(a[123] & b[171])^(a[122] & b[172])^(a[121] & b[173])^(a[120] & b[174])^(a[119] & b[175])^(a[118] & b[176])^(a[117] & b[177])^(a[116] & b[178])^(a[115] & b[179])^(a[114] & b[180])^(a[113] & b[181])^(a[112] & b[182])^(a[111] & b[183])^(a[110] & b[184])^(a[109] & b[185])^(a[108] & b[186])^(a[107] & b[187])^(a[106] & b[188])^(a[105] & b[189])^(a[104] & b[190])^(a[103] & b[191])^(a[102] & b[192])^(a[101] & b[193])^(a[100] & b[194])^(a[99] & b[195])^(a[98] & b[196])^(a[97] & b[197])^(a[96] & b[198])^(a[95] & b[199])^(a[94] & b[200])^(a[93] & b[201])^(a[92] & b[202])^(a[91] & b[203])^(a[90] & b[204])^(a[89] & b[205])^(a[88] & b[206])^(a[87] & b[207])^(a[86] & b[208])^(a[85] & b[209])^(a[84] & b[210])^(a[83] & b[211])^(a[82] & b[212])^(a[81] & b[213])^(a[80] & b[214])^(a[79] & b[215])^(a[78] & b[216])^(a[77] & b[217])^(a[76] & b[218])^(a[75] & b[219])^(a[74] & b[220])^(a[73] & b[221])^(a[72] & b[222])^(a[71] & b[223])^(a[70] & b[224])^(a[69] & b[225])^(a[68] & b[226])^(a[67] & b[227])^(a[66] & b[228])^(a[65] & b[229])^(a[64] & b[230])^(a[63] & b[231])^(a[62] & b[232]);
assign y[295] = (a[232] & b[63])^(a[231] & b[64])^(a[230] & b[65])^(a[229] & b[66])^(a[228] & b[67])^(a[227] & b[68])^(a[226] & b[69])^(a[225] & b[70])^(a[224] & b[71])^(a[223] & b[72])^(a[222] & b[73])^(a[221] & b[74])^(a[220] & b[75])^(a[219] & b[76])^(a[218] & b[77])^(a[217] & b[78])^(a[216] & b[79])^(a[215] & b[80])^(a[214] & b[81])^(a[213] & b[82])^(a[212] & b[83])^(a[211] & b[84])^(a[210] & b[85])^(a[209] & b[86])^(a[208] & b[87])^(a[207] & b[88])^(a[206] & b[89])^(a[205] & b[90])^(a[204] & b[91])^(a[203] & b[92])^(a[202] & b[93])^(a[201] & b[94])^(a[200] & b[95])^(a[199] & b[96])^(a[198] & b[97])^(a[197] & b[98])^(a[196] & b[99])^(a[195] & b[100])^(a[194] & b[101])^(a[193] & b[102])^(a[192] & b[103])^(a[191] & b[104])^(a[190] & b[105])^(a[189] & b[106])^(a[188] & b[107])^(a[187] & b[108])^(a[186] & b[109])^(a[185] & b[110])^(a[184] & b[111])^(a[183] & b[112])^(a[182] & b[113])^(a[181] & b[114])^(a[180] & b[115])^(a[179] & b[116])^(a[178] & b[117])^(a[177] & b[118])^(a[176] & b[119])^(a[175] & b[120])^(a[174] & b[121])^(a[173] & b[122])^(a[172] & b[123])^(a[171] & b[124])^(a[170] & b[125])^(a[169] & b[126])^(a[168] & b[127])^(a[167] & b[128])^(a[166] & b[129])^(a[165] & b[130])^(a[164] & b[131])^(a[163] & b[132])^(a[162] & b[133])^(a[161] & b[134])^(a[160] & b[135])^(a[159] & b[136])^(a[158] & b[137])^(a[157] & b[138])^(a[156] & b[139])^(a[155] & b[140])^(a[154] & b[141])^(a[153] & b[142])^(a[152] & b[143])^(a[151] & b[144])^(a[150] & b[145])^(a[149] & b[146])^(a[148] & b[147])^(a[147] & b[148])^(a[146] & b[149])^(a[145] & b[150])^(a[144] & b[151])^(a[143] & b[152])^(a[142] & b[153])^(a[141] & b[154])^(a[140] & b[155])^(a[139] & b[156])^(a[138] & b[157])^(a[137] & b[158])^(a[136] & b[159])^(a[135] & b[160])^(a[134] & b[161])^(a[133] & b[162])^(a[132] & b[163])^(a[131] & b[164])^(a[130] & b[165])^(a[129] & b[166])^(a[128] & b[167])^(a[127] & b[168])^(a[126] & b[169])^(a[125] & b[170])^(a[124] & b[171])^(a[123] & b[172])^(a[122] & b[173])^(a[121] & b[174])^(a[120] & b[175])^(a[119] & b[176])^(a[118] & b[177])^(a[117] & b[178])^(a[116] & b[179])^(a[115] & b[180])^(a[114] & b[181])^(a[113] & b[182])^(a[112] & b[183])^(a[111] & b[184])^(a[110] & b[185])^(a[109] & b[186])^(a[108] & b[187])^(a[107] & b[188])^(a[106] & b[189])^(a[105] & b[190])^(a[104] & b[191])^(a[103] & b[192])^(a[102] & b[193])^(a[101] & b[194])^(a[100] & b[195])^(a[99] & b[196])^(a[98] & b[197])^(a[97] & b[198])^(a[96] & b[199])^(a[95] & b[200])^(a[94] & b[201])^(a[93] & b[202])^(a[92] & b[203])^(a[91] & b[204])^(a[90] & b[205])^(a[89] & b[206])^(a[88] & b[207])^(a[87] & b[208])^(a[86] & b[209])^(a[85] & b[210])^(a[84] & b[211])^(a[83] & b[212])^(a[82] & b[213])^(a[81] & b[214])^(a[80] & b[215])^(a[79] & b[216])^(a[78] & b[217])^(a[77] & b[218])^(a[76] & b[219])^(a[75] & b[220])^(a[74] & b[221])^(a[73] & b[222])^(a[72] & b[223])^(a[71] & b[224])^(a[70] & b[225])^(a[69] & b[226])^(a[68] & b[227])^(a[67] & b[228])^(a[66] & b[229])^(a[65] & b[230])^(a[64] & b[231])^(a[63] & b[232]);
assign y[296] = (a[232] & b[64])^(a[231] & b[65])^(a[230] & b[66])^(a[229] & b[67])^(a[228] & b[68])^(a[227] & b[69])^(a[226] & b[70])^(a[225] & b[71])^(a[224] & b[72])^(a[223] & b[73])^(a[222] & b[74])^(a[221] & b[75])^(a[220] & b[76])^(a[219] & b[77])^(a[218] & b[78])^(a[217] & b[79])^(a[216] & b[80])^(a[215] & b[81])^(a[214] & b[82])^(a[213] & b[83])^(a[212] & b[84])^(a[211] & b[85])^(a[210] & b[86])^(a[209] & b[87])^(a[208] & b[88])^(a[207] & b[89])^(a[206] & b[90])^(a[205] & b[91])^(a[204] & b[92])^(a[203] & b[93])^(a[202] & b[94])^(a[201] & b[95])^(a[200] & b[96])^(a[199] & b[97])^(a[198] & b[98])^(a[197] & b[99])^(a[196] & b[100])^(a[195] & b[101])^(a[194] & b[102])^(a[193] & b[103])^(a[192] & b[104])^(a[191] & b[105])^(a[190] & b[106])^(a[189] & b[107])^(a[188] & b[108])^(a[187] & b[109])^(a[186] & b[110])^(a[185] & b[111])^(a[184] & b[112])^(a[183] & b[113])^(a[182] & b[114])^(a[181] & b[115])^(a[180] & b[116])^(a[179] & b[117])^(a[178] & b[118])^(a[177] & b[119])^(a[176] & b[120])^(a[175] & b[121])^(a[174] & b[122])^(a[173] & b[123])^(a[172] & b[124])^(a[171] & b[125])^(a[170] & b[126])^(a[169] & b[127])^(a[168] & b[128])^(a[167] & b[129])^(a[166] & b[130])^(a[165] & b[131])^(a[164] & b[132])^(a[163] & b[133])^(a[162] & b[134])^(a[161] & b[135])^(a[160] & b[136])^(a[159] & b[137])^(a[158] & b[138])^(a[157] & b[139])^(a[156] & b[140])^(a[155] & b[141])^(a[154] & b[142])^(a[153] & b[143])^(a[152] & b[144])^(a[151] & b[145])^(a[150] & b[146])^(a[149] & b[147])^(a[148] & b[148])^(a[147] & b[149])^(a[146] & b[150])^(a[145] & b[151])^(a[144] & b[152])^(a[143] & b[153])^(a[142] & b[154])^(a[141] & b[155])^(a[140] & b[156])^(a[139] & b[157])^(a[138] & b[158])^(a[137] & b[159])^(a[136] & b[160])^(a[135] & b[161])^(a[134] & b[162])^(a[133] & b[163])^(a[132] & b[164])^(a[131] & b[165])^(a[130] & b[166])^(a[129] & b[167])^(a[128] & b[168])^(a[127] & b[169])^(a[126] & b[170])^(a[125] & b[171])^(a[124] & b[172])^(a[123] & b[173])^(a[122] & b[174])^(a[121] & b[175])^(a[120] & b[176])^(a[119] & b[177])^(a[118] & b[178])^(a[117] & b[179])^(a[116] & b[180])^(a[115] & b[181])^(a[114] & b[182])^(a[113] & b[183])^(a[112] & b[184])^(a[111] & b[185])^(a[110] & b[186])^(a[109] & b[187])^(a[108] & b[188])^(a[107] & b[189])^(a[106] & b[190])^(a[105] & b[191])^(a[104] & b[192])^(a[103] & b[193])^(a[102] & b[194])^(a[101] & b[195])^(a[100] & b[196])^(a[99] & b[197])^(a[98] & b[198])^(a[97] & b[199])^(a[96] & b[200])^(a[95] & b[201])^(a[94] & b[202])^(a[93] & b[203])^(a[92] & b[204])^(a[91] & b[205])^(a[90] & b[206])^(a[89] & b[207])^(a[88] & b[208])^(a[87] & b[209])^(a[86] & b[210])^(a[85] & b[211])^(a[84] & b[212])^(a[83] & b[213])^(a[82] & b[214])^(a[81] & b[215])^(a[80] & b[216])^(a[79] & b[217])^(a[78] & b[218])^(a[77] & b[219])^(a[76] & b[220])^(a[75] & b[221])^(a[74] & b[222])^(a[73] & b[223])^(a[72] & b[224])^(a[71] & b[225])^(a[70] & b[226])^(a[69] & b[227])^(a[68] & b[228])^(a[67] & b[229])^(a[66] & b[230])^(a[65] & b[231])^(a[64] & b[232]);
assign y[297] = (a[232] & b[65])^(a[231] & b[66])^(a[230] & b[67])^(a[229] & b[68])^(a[228] & b[69])^(a[227] & b[70])^(a[226] & b[71])^(a[225] & b[72])^(a[224] & b[73])^(a[223] & b[74])^(a[222] & b[75])^(a[221] & b[76])^(a[220] & b[77])^(a[219] & b[78])^(a[218] & b[79])^(a[217] & b[80])^(a[216] & b[81])^(a[215] & b[82])^(a[214] & b[83])^(a[213] & b[84])^(a[212] & b[85])^(a[211] & b[86])^(a[210] & b[87])^(a[209] & b[88])^(a[208] & b[89])^(a[207] & b[90])^(a[206] & b[91])^(a[205] & b[92])^(a[204] & b[93])^(a[203] & b[94])^(a[202] & b[95])^(a[201] & b[96])^(a[200] & b[97])^(a[199] & b[98])^(a[198] & b[99])^(a[197] & b[100])^(a[196] & b[101])^(a[195] & b[102])^(a[194] & b[103])^(a[193] & b[104])^(a[192] & b[105])^(a[191] & b[106])^(a[190] & b[107])^(a[189] & b[108])^(a[188] & b[109])^(a[187] & b[110])^(a[186] & b[111])^(a[185] & b[112])^(a[184] & b[113])^(a[183] & b[114])^(a[182] & b[115])^(a[181] & b[116])^(a[180] & b[117])^(a[179] & b[118])^(a[178] & b[119])^(a[177] & b[120])^(a[176] & b[121])^(a[175] & b[122])^(a[174] & b[123])^(a[173] & b[124])^(a[172] & b[125])^(a[171] & b[126])^(a[170] & b[127])^(a[169] & b[128])^(a[168] & b[129])^(a[167] & b[130])^(a[166] & b[131])^(a[165] & b[132])^(a[164] & b[133])^(a[163] & b[134])^(a[162] & b[135])^(a[161] & b[136])^(a[160] & b[137])^(a[159] & b[138])^(a[158] & b[139])^(a[157] & b[140])^(a[156] & b[141])^(a[155] & b[142])^(a[154] & b[143])^(a[153] & b[144])^(a[152] & b[145])^(a[151] & b[146])^(a[150] & b[147])^(a[149] & b[148])^(a[148] & b[149])^(a[147] & b[150])^(a[146] & b[151])^(a[145] & b[152])^(a[144] & b[153])^(a[143] & b[154])^(a[142] & b[155])^(a[141] & b[156])^(a[140] & b[157])^(a[139] & b[158])^(a[138] & b[159])^(a[137] & b[160])^(a[136] & b[161])^(a[135] & b[162])^(a[134] & b[163])^(a[133] & b[164])^(a[132] & b[165])^(a[131] & b[166])^(a[130] & b[167])^(a[129] & b[168])^(a[128] & b[169])^(a[127] & b[170])^(a[126] & b[171])^(a[125] & b[172])^(a[124] & b[173])^(a[123] & b[174])^(a[122] & b[175])^(a[121] & b[176])^(a[120] & b[177])^(a[119] & b[178])^(a[118] & b[179])^(a[117] & b[180])^(a[116] & b[181])^(a[115] & b[182])^(a[114] & b[183])^(a[113] & b[184])^(a[112] & b[185])^(a[111] & b[186])^(a[110] & b[187])^(a[109] & b[188])^(a[108] & b[189])^(a[107] & b[190])^(a[106] & b[191])^(a[105] & b[192])^(a[104] & b[193])^(a[103] & b[194])^(a[102] & b[195])^(a[101] & b[196])^(a[100] & b[197])^(a[99] & b[198])^(a[98] & b[199])^(a[97] & b[200])^(a[96] & b[201])^(a[95] & b[202])^(a[94] & b[203])^(a[93] & b[204])^(a[92] & b[205])^(a[91] & b[206])^(a[90] & b[207])^(a[89] & b[208])^(a[88] & b[209])^(a[87] & b[210])^(a[86] & b[211])^(a[85] & b[212])^(a[84] & b[213])^(a[83] & b[214])^(a[82] & b[215])^(a[81] & b[216])^(a[80] & b[217])^(a[79] & b[218])^(a[78] & b[219])^(a[77] & b[220])^(a[76] & b[221])^(a[75] & b[222])^(a[74] & b[223])^(a[73] & b[224])^(a[72] & b[225])^(a[71] & b[226])^(a[70] & b[227])^(a[69] & b[228])^(a[68] & b[229])^(a[67] & b[230])^(a[66] & b[231])^(a[65] & b[232]);
assign y[298] = (a[232] & b[66])^(a[231] & b[67])^(a[230] & b[68])^(a[229] & b[69])^(a[228] & b[70])^(a[227] & b[71])^(a[226] & b[72])^(a[225] & b[73])^(a[224] & b[74])^(a[223] & b[75])^(a[222] & b[76])^(a[221] & b[77])^(a[220] & b[78])^(a[219] & b[79])^(a[218] & b[80])^(a[217] & b[81])^(a[216] & b[82])^(a[215] & b[83])^(a[214] & b[84])^(a[213] & b[85])^(a[212] & b[86])^(a[211] & b[87])^(a[210] & b[88])^(a[209] & b[89])^(a[208] & b[90])^(a[207] & b[91])^(a[206] & b[92])^(a[205] & b[93])^(a[204] & b[94])^(a[203] & b[95])^(a[202] & b[96])^(a[201] & b[97])^(a[200] & b[98])^(a[199] & b[99])^(a[198] & b[100])^(a[197] & b[101])^(a[196] & b[102])^(a[195] & b[103])^(a[194] & b[104])^(a[193] & b[105])^(a[192] & b[106])^(a[191] & b[107])^(a[190] & b[108])^(a[189] & b[109])^(a[188] & b[110])^(a[187] & b[111])^(a[186] & b[112])^(a[185] & b[113])^(a[184] & b[114])^(a[183] & b[115])^(a[182] & b[116])^(a[181] & b[117])^(a[180] & b[118])^(a[179] & b[119])^(a[178] & b[120])^(a[177] & b[121])^(a[176] & b[122])^(a[175] & b[123])^(a[174] & b[124])^(a[173] & b[125])^(a[172] & b[126])^(a[171] & b[127])^(a[170] & b[128])^(a[169] & b[129])^(a[168] & b[130])^(a[167] & b[131])^(a[166] & b[132])^(a[165] & b[133])^(a[164] & b[134])^(a[163] & b[135])^(a[162] & b[136])^(a[161] & b[137])^(a[160] & b[138])^(a[159] & b[139])^(a[158] & b[140])^(a[157] & b[141])^(a[156] & b[142])^(a[155] & b[143])^(a[154] & b[144])^(a[153] & b[145])^(a[152] & b[146])^(a[151] & b[147])^(a[150] & b[148])^(a[149] & b[149])^(a[148] & b[150])^(a[147] & b[151])^(a[146] & b[152])^(a[145] & b[153])^(a[144] & b[154])^(a[143] & b[155])^(a[142] & b[156])^(a[141] & b[157])^(a[140] & b[158])^(a[139] & b[159])^(a[138] & b[160])^(a[137] & b[161])^(a[136] & b[162])^(a[135] & b[163])^(a[134] & b[164])^(a[133] & b[165])^(a[132] & b[166])^(a[131] & b[167])^(a[130] & b[168])^(a[129] & b[169])^(a[128] & b[170])^(a[127] & b[171])^(a[126] & b[172])^(a[125] & b[173])^(a[124] & b[174])^(a[123] & b[175])^(a[122] & b[176])^(a[121] & b[177])^(a[120] & b[178])^(a[119] & b[179])^(a[118] & b[180])^(a[117] & b[181])^(a[116] & b[182])^(a[115] & b[183])^(a[114] & b[184])^(a[113] & b[185])^(a[112] & b[186])^(a[111] & b[187])^(a[110] & b[188])^(a[109] & b[189])^(a[108] & b[190])^(a[107] & b[191])^(a[106] & b[192])^(a[105] & b[193])^(a[104] & b[194])^(a[103] & b[195])^(a[102] & b[196])^(a[101] & b[197])^(a[100] & b[198])^(a[99] & b[199])^(a[98] & b[200])^(a[97] & b[201])^(a[96] & b[202])^(a[95] & b[203])^(a[94] & b[204])^(a[93] & b[205])^(a[92] & b[206])^(a[91] & b[207])^(a[90] & b[208])^(a[89] & b[209])^(a[88] & b[210])^(a[87] & b[211])^(a[86] & b[212])^(a[85] & b[213])^(a[84] & b[214])^(a[83] & b[215])^(a[82] & b[216])^(a[81] & b[217])^(a[80] & b[218])^(a[79] & b[219])^(a[78] & b[220])^(a[77] & b[221])^(a[76] & b[222])^(a[75] & b[223])^(a[74] & b[224])^(a[73] & b[225])^(a[72] & b[226])^(a[71] & b[227])^(a[70] & b[228])^(a[69] & b[229])^(a[68] & b[230])^(a[67] & b[231])^(a[66] & b[232]);
assign y[299] = (a[232] & b[67])^(a[231] & b[68])^(a[230] & b[69])^(a[229] & b[70])^(a[228] & b[71])^(a[227] & b[72])^(a[226] & b[73])^(a[225] & b[74])^(a[224] & b[75])^(a[223] & b[76])^(a[222] & b[77])^(a[221] & b[78])^(a[220] & b[79])^(a[219] & b[80])^(a[218] & b[81])^(a[217] & b[82])^(a[216] & b[83])^(a[215] & b[84])^(a[214] & b[85])^(a[213] & b[86])^(a[212] & b[87])^(a[211] & b[88])^(a[210] & b[89])^(a[209] & b[90])^(a[208] & b[91])^(a[207] & b[92])^(a[206] & b[93])^(a[205] & b[94])^(a[204] & b[95])^(a[203] & b[96])^(a[202] & b[97])^(a[201] & b[98])^(a[200] & b[99])^(a[199] & b[100])^(a[198] & b[101])^(a[197] & b[102])^(a[196] & b[103])^(a[195] & b[104])^(a[194] & b[105])^(a[193] & b[106])^(a[192] & b[107])^(a[191] & b[108])^(a[190] & b[109])^(a[189] & b[110])^(a[188] & b[111])^(a[187] & b[112])^(a[186] & b[113])^(a[185] & b[114])^(a[184] & b[115])^(a[183] & b[116])^(a[182] & b[117])^(a[181] & b[118])^(a[180] & b[119])^(a[179] & b[120])^(a[178] & b[121])^(a[177] & b[122])^(a[176] & b[123])^(a[175] & b[124])^(a[174] & b[125])^(a[173] & b[126])^(a[172] & b[127])^(a[171] & b[128])^(a[170] & b[129])^(a[169] & b[130])^(a[168] & b[131])^(a[167] & b[132])^(a[166] & b[133])^(a[165] & b[134])^(a[164] & b[135])^(a[163] & b[136])^(a[162] & b[137])^(a[161] & b[138])^(a[160] & b[139])^(a[159] & b[140])^(a[158] & b[141])^(a[157] & b[142])^(a[156] & b[143])^(a[155] & b[144])^(a[154] & b[145])^(a[153] & b[146])^(a[152] & b[147])^(a[151] & b[148])^(a[150] & b[149])^(a[149] & b[150])^(a[148] & b[151])^(a[147] & b[152])^(a[146] & b[153])^(a[145] & b[154])^(a[144] & b[155])^(a[143] & b[156])^(a[142] & b[157])^(a[141] & b[158])^(a[140] & b[159])^(a[139] & b[160])^(a[138] & b[161])^(a[137] & b[162])^(a[136] & b[163])^(a[135] & b[164])^(a[134] & b[165])^(a[133] & b[166])^(a[132] & b[167])^(a[131] & b[168])^(a[130] & b[169])^(a[129] & b[170])^(a[128] & b[171])^(a[127] & b[172])^(a[126] & b[173])^(a[125] & b[174])^(a[124] & b[175])^(a[123] & b[176])^(a[122] & b[177])^(a[121] & b[178])^(a[120] & b[179])^(a[119] & b[180])^(a[118] & b[181])^(a[117] & b[182])^(a[116] & b[183])^(a[115] & b[184])^(a[114] & b[185])^(a[113] & b[186])^(a[112] & b[187])^(a[111] & b[188])^(a[110] & b[189])^(a[109] & b[190])^(a[108] & b[191])^(a[107] & b[192])^(a[106] & b[193])^(a[105] & b[194])^(a[104] & b[195])^(a[103] & b[196])^(a[102] & b[197])^(a[101] & b[198])^(a[100] & b[199])^(a[99] & b[200])^(a[98] & b[201])^(a[97] & b[202])^(a[96] & b[203])^(a[95] & b[204])^(a[94] & b[205])^(a[93] & b[206])^(a[92] & b[207])^(a[91] & b[208])^(a[90] & b[209])^(a[89] & b[210])^(a[88] & b[211])^(a[87] & b[212])^(a[86] & b[213])^(a[85] & b[214])^(a[84] & b[215])^(a[83] & b[216])^(a[82] & b[217])^(a[81] & b[218])^(a[80] & b[219])^(a[79] & b[220])^(a[78] & b[221])^(a[77] & b[222])^(a[76] & b[223])^(a[75] & b[224])^(a[74] & b[225])^(a[73] & b[226])^(a[72] & b[227])^(a[71] & b[228])^(a[70] & b[229])^(a[69] & b[230])^(a[68] & b[231])^(a[67] & b[232]);
assign y[300] = (a[232] & b[68])^(a[231] & b[69])^(a[230] & b[70])^(a[229] & b[71])^(a[228] & b[72])^(a[227] & b[73])^(a[226] & b[74])^(a[225] & b[75])^(a[224] & b[76])^(a[223] & b[77])^(a[222] & b[78])^(a[221] & b[79])^(a[220] & b[80])^(a[219] & b[81])^(a[218] & b[82])^(a[217] & b[83])^(a[216] & b[84])^(a[215] & b[85])^(a[214] & b[86])^(a[213] & b[87])^(a[212] & b[88])^(a[211] & b[89])^(a[210] & b[90])^(a[209] & b[91])^(a[208] & b[92])^(a[207] & b[93])^(a[206] & b[94])^(a[205] & b[95])^(a[204] & b[96])^(a[203] & b[97])^(a[202] & b[98])^(a[201] & b[99])^(a[200] & b[100])^(a[199] & b[101])^(a[198] & b[102])^(a[197] & b[103])^(a[196] & b[104])^(a[195] & b[105])^(a[194] & b[106])^(a[193] & b[107])^(a[192] & b[108])^(a[191] & b[109])^(a[190] & b[110])^(a[189] & b[111])^(a[188] & b[112])^(a[187] & b[113])^(a[186] & b[114])^(a[185] & b[115])^(a[184] & b[116])^(a[183] & b[117])^(a[182] & b[118])^(a[181] & b[119])^(a[180] & b[120])^(a[179] & b[121])^(a[178] & b[122])^(a[177] & b[123])^(a[176] & b[124])^(a[175] & b[125])^(a[174] & b[126])^(a[173] & b[127])^(a[172] & b[128])^(a[171] & b[129])^(a[170] & b[130])^(a[169] & b[131])^(a[168] & b[132])^(a[167] & b[133])^(a[166] & b[134])^(a[165] & b[135])^(a[164] & b[136])^(a[163] & b[137])^(a[162] & b[138])^(a[161] & b[139])^(a[160] & b[140])^(a[159] & b[141])^(a[158] & b[142])^(a[157] & b[143])^(a[156] & b[144])^(a[155] & b[145])^(a[154] & b[146])^(a[153] & b[147])^(a[152] & b[148])^(a[151] & b[149])^(a[150] & b[150])^(a[149] & b[151])^(a[148] & b[152])^(a[147] & b[153])^(a[146] & b[154])^(a[145] & b[155])^(a[144] & b[156])^(a[143] & b[157])^(a[142] & b[158])^(a[141] & b[159])^(a[140] & b[160])^(a[139] & b[161])^(a[138] & b[162])^(a[137] & b[163])^(a[136] & b[164])^(a[135] & b[165])^(a[134] & b[166])^(a[133] & b[167])^(a[132] & b[168])^(a[131] & b[169])^(a[130] & b[170])^(a[129] & b[171])^(a[128] & b[172])^(a[127] & b[173])^(a[126] & b[174])^(a[125] & b[175])^(a[124] & b[176])^(a[123] & b[177])^(a[122] & b[178])^(a[121] & b[179])^(a[120] & b[180])^(a[119] & b[181])^(a[118] & b[182])^(a[117] & b[183])^(a[116] & b[184])^(a[115] & b[185])^(a[114] & b[186])^(a[113] & b[187])^(a[112] & b[188])^(a[111] & b[189])^(a[110] & b[190])^(a[109] & b[191])^(a[108] & b[192])^(a[107] & b[193])^(a[106] & b[194])^(a[105] & b[195])^(a[104] & b[196])^(a[103] & b[197])^(a[102] & b[198])^(a[101] & b[199])^(a[100] & b[200])^(a[99] & b[201])^(a[98] & b[202])^(a[97] & b[203])^(a[96] & b[204])^(a[95] & b[205])^(a[94] & b[206])^(a[93] & b[207])^(a[92] & b[208])^(a[91] & b[209])^(a[90] & b[210])^(a[89] & b[211])^(a[88] & b[212])^(a[87] & b[213])^(a[86] & b[214])^(a[85] & b[215])^(a[84] & b[216])^(a[83] & b[217])^(a[82] & b[218])^(a[81] & b[219])^(a[80] & b[220])^(a[79] & b[221])^(a[78] & b[222])^(a[77] & b[223])^(a[76] & b[224])^(a[75] & b[225])^(a[74] & b[226])^(a[73] & b[227])^(a[72] & b[228])^(a[71] & b[229])^(a[70] & b[230])^(a[69] & b[231])^(a[68] & b[232]);
assign y[301] = (a[232] & b[69])^(a[231] & b[70])^(a[230] & b[71])^(a[229] & b[72])^(a[228] & b[73])^(a[227] & b[74])^(a[226] & b[75])^(a[225] & b[76])^(a[224] & b[77])^(a[223] & b[78])^(a[222] & b[79])^(a[221] & b[80])^(a[220] & b[81])^(a[219] & b[82])^(a[218] & b[83])^(a[217] & b[84])^(a[216] & b[85])^(a[215] & b[86])^(a[214] & b[87])^(a[213] & b[88])^(a[212] & b[89])^(a[211] & b[90])^(a[210] & b[91])^(a[209] & b[92])^(a[208] & b[93])^(a[207] & b[94])^(a[206] & b[95])^(a[205] & b[96])^(a[204] & b[97])^(a[203] & b[98])^(a[202] & b[99])^(a[201] & b[100])^(a[200] & b[101])^(a[199] & b[102])^(a[198] & b[103])^(a[197] & b[104])^(a[196] & b[105])^(a[195] & b[106])^(a[194] & b[107])^(a[193] & b[108])^(a[192] & b[109])^(a[191] & b[110])^(a[190] & b[111])^(a[189] & b[112])^(a[188] & b[113])^(a[187] & b[114])^(a[186] & b[115])^(a[185] & b[116])^(a[184] & b[117])^(a[183] & b[118])^(a[182] & b[119])^(a[181] & b[120])^(a[180] & b[121])^(a[179] & b[122])^(a[178] & b[123])^(a[177] & b[124])^(a[176] & b[125])^(a[175] & b[126])^(a[174] & b[127])^(a[173] & b[128])^(a[172] & b[129])^(a[171] & b[130])^(a[170] & b[131])^(a[169] & b[132])^(a[168] & b[133])^(a[167] & b[134])^(a[166] & b[135])^(a[165] & b[136])^(a[164] & b[137])^(a[163] & b[138])^(a[162] & b[139])^(a[161] & b[140])^(a[160] & b[141])^(a[159] & b[142])^(a[158] & b[143])^(a[157] & b[144])^(a[156] & b[145])^(a[155] & b[146])^(a[154] & b[147])^(a[153] & b[148])^(a[152] & b[149])^(a[151] & b[150])^(a[150] & b[151])^(a[149] & b[152])^(a[148] & b[153])^(a[147] & b[154])^(a[146] & b[155])^(a[145] & b[156])^(a[144] & b[157])^(a[143] & b[158])^(a[142] & b[159])^(a[141] & b[160])^(a[140] & b[161])^(a[139] & b[162])^(a[138] & b[163])^(a[137] & b[164])^(a[136] & b[165])^(a[135] & b[166])^(a[134] & b[167])^(a[133] & b[168])^(a[132] & b[169])^(a[131] & b[170])^(a[130] & b[171])^(a[129] & b[172])^(a[128] & b[173])^(a[127] & b[174])^(a[126] & b[175])^(a[125] & b[176])^(a[124] & b[177])^(a[123] & b[178])^(a[122] & b[179])^(a[121] & b[180])^(a[120] & b[181])^(a[119] & b[182])^(a[118] & b[183])^(a[117] & b[184])^(a[116] & b[185])^(a[115] & b[186])^(a[114] & b[187])^(a[113] & b[188])^(a[112] & b[189])^(a[111] & b[190])^(a[110] & b[191])^(a[109] & b[192])^(a[108] & b[193])^(a[107] & b[194])^(a[106] & b[195])^(a[105] & b[196])^(a[104] & b[197])^(a[103] & b[198])^(a[102] & b[199])^(a[101] & b[200])^(a[100] & b[201])^(a[99] & b[202])^(a[98] & b[203])^(a[97] & b[204])^(a[96] & b[205])^(a[95] & b[206])^(a[94] & b[207])^(a[93] & b[208])^(a[92] & b[209])^(a[91] & b[210])^(a[90] & b[211])^(a[89] & b[212])^(a[88] & b[213])^(a[87] & b[214])^(a[86] & b[215])^(a[85] & b[216])^(a[84] & b[217])^(a[83] & b[218])^(a[82] & b[219])^(a[81] & b[220])^(a[80] & b[221])^(a[79] & b[222])^(a[78] & b[223])^(a[77] & b[224])^(a[76] & b[225])^(a[75] & b[226])^(a[74] & b[227])^(a[73] & b[228])^(a[72] & b[229])^(a[71] & b[230])^(a[70] & b[231])^(a[69] & b[232]);
assign y[302] = (a[232] & b[70])^(a[231] & b[71])^(a[230] & b[72])^(a[229] & b[73])^(a[228] & b[74])^(a[227] & b[75])^(a[226] & b[76])^(a[225] & b[77])^(a[224] & b[78])^(a[223] & b[79])^(a[222] & b[80])^(a[221] & b[81])^(a[220] & b[82])^(a[219] & b[83])^(a[218] & b[84])^(a[217] & b[85])^(a[216] & b[86])^(a[215] & b[87])^(a[214] & b[88])^(a[213] & b[89])^(a[212] & b[90])^(a[211] & b[91])^(a[210] & b[92])^(a[209] & b[93])^(a[208] & b[94])^(a[207] & b[95])^(a[206] & b[96])^(a[205] & b[97])^(a[204] & b[98])^(a[203] & b[99])^(a[202] & b[100])^(a[201] & b[101])^(a[200] & b[102])^(a[199] & b[103])^(a[198] & b[104])^(a[197] & b[105])^(a[196] & b[106])^(a[195] & b[107])^(a[194] & b[108])^(a[193] & b[109])^(a[192] & b[110])^(a[191] & b[111])^(a[190] & b[112])^(a[189] & b[113])^(a[188] & b[114])^(a[187] & b[115])^(a[186] & b[116])^(a[185] & b[117])^(a[184] & b[118])^(a[183] & b[119])^(a[182] & b[120])^(a[181] & b[121])^(a[180] & b[122])^(a[179] & b[123])^(a[178] & b[124])^(a[177] & b[125])^(a[176] & b[126])^(a[175] & b[127])^(a[174] & b[128])^(a[173] & b[129])^(a[172] & b[130])^(a[171] & b[131])^(a[170] & b[132])^(a[169] & b[133])^(a[168] & b[134])^(a[167] & b[135])^(a[166] & b[136])^(a[165] & b[137])^(a[164] & b[138])^(a[163] & b[139])^(a[162] & b[140])^(a[161] & b[141])^(a[160] & b[142])^(a[159] & b[143])^(a[158] & b[144])^(a[157] & b[145])^(a[156] & b[146])^(a[155] & b[147])^(a[154] & b[148])^(a[153] & b[149])^(a[152] & b[150])^(a[151] & b[151])^(a[150] & b[152])^(a[149] & b[153])^(a[148] & b[154])^(a[147] & b[155])^(a[146] & b[156])^(a[145] & b[157])^(a[144] & b[158])^(a[143] & b[159])^(a[142] & b[160])^(a[141] & b[161])^(a[140] & b[162])^(a[139] & b[163])^(a[138] & b[164])^(a[137] & b[165])^(a[136] & b[166])^(a[135] & b[167])^(a[134] & b[168])^(a[133] & b[169])^(a[132] & b[170])^(a[131] & b[171])^(a[130] & b[172])^(a[129] & b[173])^(a[128] & b[174])^(a[127] & b[175])^(a[126] & b[176])^(a[125] & b[177])^(a[124] & b[178])^(a[123] & b[179])^(a[122] & b[180])^(a[121] & b[181])^(a[120] & b[182])^(a[119] & b[183])^(a[118] & b[184])^(a[117] & b[185])^(a[116] & b[186])^(a[115] & b[187])^(a[114] & b[188])^(a[113] & b[189])^(a[112] & b[190])^(a[111] & b[191])^(a[110] & b[192])^(a[109] & b[193])^(a[108] & b[194])^(a[107] & b[195])^(a[106] & b[196])^(a[105] & b[197])^(a[104] & b[198])^(a[103] & b[199])^(a[102] & b[200])^(a[101] & b[201])^(a[100] & b[202])^(a[99] & b[203])^(a[98] & b[204])^(a[97] & b[205])^(a[96] & b[206])^(a[95] & b[207])^(a[94] & b[208])^(a[93] & b[209])^(a[92] & b[210])^(a[91] & b[211])^(a[90] & b[212])^(a[89] & b[213])^(a[88] & b[214])^(a[87] & b[215])^(a[86] & b[216])^(a[85] & b[217])^(a[84] & b[218])^(a[83] & b[219])^(a[82] & b[220])^(a[81] & b[221])^(a[80] & b[222])^(a[79] & b[223])^(a[78] & b[224])^(a[77] & b[225])^(a[76] & b[226])^(a[75] & b[227])^(a[74] & b[228])^(a[73] & b[229])^(a[72] & b[230])^(a[71] & b[231])^(a[70] & b[232]);
assign y[303] = (a[232] & b[71])^(a[231] & b[72])^(a[230] & b[73])^(a[229] & b[74])^(a[228] & b[75])^(a[227] & b[76])^(a[226] & b[77])^(a[225] & b[78])^(a[224] & b[79])^(a[223] & b[80])^(a[222] & b[81])^(a[221] & b[82])^(a[220] & b[83])^(a[219] & b[84])^(a[218] & b[85])^(a[217] & b[86])^(a[216] & b[87])^(a[215] & b[88])^(a[214] & b[89])^(a[213] & b[90])^(a[212] & b[91])^(a[211] & b[92])^(a[210] & b[93])^(a[209] & b[94])^(a[208] & b[95])^(a[207] & b[96])^(a[206] & b[97])^(a[205] & b[98])^(a[204] & b[99])^(a[203] & b[100])^(a[202] & b[101])^(a[201] & b[102])^(a[200] & b[103])^(a[199] & b[104])^(a[198] & b[105])^(a[197] & b[106])^(a[196] & b[107])^(a[195] & b[108])^(a[194] & b[109])^(a[193] & b[110])^(a[192] & b[111])^(a[191] & b[112])^(a[190] & b[113])^(a[189] & b[114])^(a[188] & b[115])^(a[187] & b[116])^(a[186] & b[117])^(a[185] & b[118])^(a[184] & b[119])^(a[183] & b[120])^(a[182] & b[121])^(a[181] & b[122])^(a[180] & b[123])^(a[179] & b[124])^(a[178] & b[125])^(a[177] & b[126])^(a[176] & b[127])^(a[175] & b[128])^(a[174] & b[129])^(a[173] & b[130])^(a[172] & b[131])^(a[171] & b[132])^(a[170] & b[133])^(a[169] & b[134])^(a[168] & b[135])^(a[167] & b[136])^(a[166] & b[137])^(a[165] & b[138])^(a[164] & b[139])^(a[163] & b[140])^(a[162] & b[141])^(a[161] & b[142])^(a[160] & b[143])^(a[159] & b[144])^(a[158] & b[145])^(a[157] & b[146])^(a[156] & b[147])^(a[155] & b[148])^(a[154] & b[149])^(a[153] & b[150])^(a[152] & b[151])^(a[151] & b[152])^(a[150] & b[153])^(a[149] & b[154])^(a[148] & b[155])^(a[147] & b[156])^(a[146] & b[157])^(a[145] & b[158])^(a[144] & b[159])^(a[143] & b[160])^(a[142] & b[161])^(a[141] & b[162])^(a[140] & b[163])^(a[139] & b[164])^(a[138] & b[165])^(a[137] & b[166])^(a[136] & b[167])^(a[135] & b[168])^(a[134] & b[169])^(a[133] & b[170])^(a[132] & b[171])^(a[131] & b[172])^(a[130] & b[173])^(a[129] & b[174])^(a[128] & b[175])^(a[127] & b[176])^(a[126] & b[177])^(a[125] & b[178])^(a[124] & b[179])^(a[123] & b[180])^(a[122] & b[181])^(a[121] & b[182])^(a[120] & b[183])^(a[119] & b[184])^(a[118] & b[185])^(a[117] & b[186])^(a[116] & b[187])^(a[115] & b[188])^(a[114] & b[189])^(a[113] & b[190])^(a[112] & b[191])^(a[111] & b[192])^(a[110] & b[193])^(a[109] & b[194])^(a[108] & b[195])^(a[107] & b[196])^(a[106] & b[197])^(a[105] & b[198])^(a[104] & b[199])^(a[103] & b[200])^(a[102] & b[201])^(a[101] & b[202])^(a[100] & b[203])^(a[99] & b[204])^(a[98] & b[205])^(a[97] & b[206])^(a[96] & b[207])^(a[95] & b[208])^(a[94] & b[209])^(a[93] & b[210])^(a[92] & b[211])^(a[91] & b[212])^(a[90] & b[213])^(a[89] & b[214])^(a[88] & b[215])^(a[87] & b[216])^(a[86] & b[217])^(a[85] & b[218])^(a[84] & b[219])^(a[83] & b[220])^(a[82] & b[221])^(a[81] & b[222])^(a[80] & b[223])^(a[79] & b[224])^(a[78] & b[225])^(a[77] & b[226])^(a[76] & b[227])^(a[75] & b[228])^(a[74] & b[229])^(a[73] & b[230])^(a[72] & b[231])^(a[71] & b[232]);
assign y[304] = (a[232] & b[72])^(a[231] & b[73])^(a[230] & b[74])^(a[229] & b[75])^(a[228] & b[76])^(a[227] & b[77])^(a[226] & b[78])^(a[225] & b[79])^(a[224] & b[80])^(a[223] & b[81])^(a[222] & b[82])^(a[221] & b[83])^(a[220] & b[84])^(a[219] & b[85])^(a[218] & b[86])^(a[217] & b[87])^(a[216] & b[88])^(a[215] & b[89])^(a[214] & b[90])^(a[213] & b[91])^(a[212] & b[92])^(a[211] & b[93])^(a[210] & b[94])^(a[209] & b[95])^(a[208] & b[96])^(a[207] & b[97])^(a[206] & b[98])^(a[205] & b[99])^(a[204] & b[100])^(a[203] & b[101])^(a[202] & b[102])^(a[201] & b[103])^(a[200] & b[104])^(a[199] & b[105])^(a[198] & b[106])^(a[197] & b[107])^(a[196] & b[108])^(a[195] & b[109])^(a[194] & b[110])^(a[193] & b[111])^(a[192] & b[112])^(a[191] & b[113])^(a[190] & b[114])^(a[189] & b[115])^(a[188] & b[116])^(a[187] & b[117])^(a[186] & b[118])^(a[185] & b[119])^(a[184] & b[120])^(a[183] & b[121])^(a[182] & b[122])^(a[181] & b[123])^(a[180] & b[124])^(a[179] & b[125])^(a[178] & b[126])^(a[177] & b[127])^(a[176] & b[128])^(a[175] & b[129])^(a[174] & b[130])^(a[173] & b[131])^(a[172] & b[132])^(a[171] & b[133])^(a[170] & b[134])^(a[169] & b[135])^(a[168] & b[136])^(a[167] & b[137])^(a[166] & b[138])^(a[165] & b[139])^(a[164] & b[140])^(a[163] & b[141])^(a[162] & b[142])^(a[161] & b[143])^(a[160] & b[144])^(a[159] & b[145])^(a[158] & b[146])^(a[157] & b[147])^(a[156] & b[148])^(a[155] & b[149])^(a[154] & b[150])^(a[153] & b[151])^(a[152] & b[152])^(a[151] & b[153])^(a[150] & b[154])^(a[149] & b[155])^(a[148] & b[156])^(a[147] & b[157])^(a[146] & b[158])^(a[145] & b[159])^(a[144] & b[160])^(a[143] & b[161])^(a[142] & b[162])^(a[141] & b[163])^(a[140] & b[164])^(a[139] & b[165])^(a[138] & b[166])^(a[137] & b[167])^(a[136] & b[168])^(a[135] & b[169])^(a[134] & b[170])^(a[133] & b[171])^(a[132] & b[172])^(a[131] & b[173])^(a[130] & b[174])^(a[129] & b[175])^(a[128] & b[176])^(a[127] & b[177])^(a[126] & b[178])^(a[125] & b[179])^(a[124] & b[180])^(a[123] & b[181])^(a[122] & b[182])^(a[121] & b[183])^(a[120] & b[184])^(a[119] & b[185])^(a[118] & b[186])^(a[117] & b[187])^(a[116] & b[188])^(a[115] & b[189])^(a[114] & b[190])^(a[113] & b[191])^(a[112] & b[192])^(a[111] & b[193])^(a[110] & b[194])^(a[109] & b[195])^(a[108] & b[196])^(a[107] & b[197])^(a[106] & b[198])^(a[105] & b[199])^(a[104] & b[200])^(a[103] & b[201])^(a[102] & b[202])^(a[101] & b[203])^(a[100] & b[204])^(a[99] & b[205])^(a[98] & b[206])^(a[97] & b[207])^(a[96] & b[208])^(a[95] & b[209])^(a[94] & b[210])^(a[93] & b[211])^(a[92] & b[212])^(a[91] & b[213])^(a[90] & b[214])^(a[89] & b[215])^(a[88] & b[216])^(a[87] & b[217])^(a[86] & b[218])^(a[85] & b[219])^(a[84] & b[220])^(a[83] & b[221])^(a[82] & b[222])^(a[81] & b[223])^(a[80] & b[224])^(a[79] & b[225])^(a[78] & b[226])^(a[77] & b[227])^(a[76] & b[228])^(a[75] & b[229])^(a[74] & b[230])^(a[73] & b[231])^(a[72] & b[232]);
assign y[305] = (a[232] & b[73])^(a[231] & b[74])^(a[230] & b[75])^(a[229] & b[76])^(a[228] & b[77])^(a[227] & b[78])^(a[226] & b[79])^(a[225] & b[80])^(a[224] & b[81])^(a[223] & b[82])^(a[222] & b[83])^(a[221] & b[84])^(a[220] & b[85])^(a[219] & b[86])^(a[218] & b[87])^(a[217] & b[88])^(a[216] & b[89])^(a[215] & b[90])^(a[214] & b[91])^(a[213] & b[92])^(a[212] & b[93])^(a[211] & b[94])^(a[210] & b[95])^(a[209] & b[96])^(a[208] & b[97])^(a[207] & b[98])^(a[206] & b[99])^(a[205] & b[100])^(a[204] & b[101])^(a[203] & b[102])^(a[202] & b[103])^(a[201] & b[104])^(a[200] & b[105])^(a[199] & b[106])^(a[198] & b[107])^(a[197] & b[108])^(a[196] & b[109])^(a[195] & b[110])^(a[194] & b[111])^(a[193] & b[112])^(a[192] & b[113])^(a[191] & b[114])^(a[190] & b[115])^(a[189] & b[116])^(a[188] & b[117])^(a[187] & b[118])^(a[186] & b[119])^(a[185] & b[120])^(a[184] & b[121])^(a[183] & b[122])^(a[182] & b[123])^(a[181] & b[124])^(a[180] & b[125])^(a[179] & b[126])^(a[178] & b[127])^(a[177] & b[128])^(a[176] & b[129])^(a[175] & b[130])^(a[174] & b[131])^(a[173] & b[132])^(a[172] & b[133])^(a[171] & b[134])^(a[170] & b[135])^(a[169] & b[136])^(a[168] & b[137])^(a[167] & b[138])^(a[166] & b[139])^(a[165] & b[140])^(a[164] & b[141])^(a[163] & b[142])^(a[162] & b[143])^(a[161] & b[144])^(a[160] & b[145])^(a[159] & b[146])^(a[158] & b[147])^(a[157] & b[148])^(a[156] & b[149])^(a[155] & b[150])^(a[154] & b[151])^(a[153] & b[152])^(a[152] & b[153])^(a[151] & b[154])^(a[150] & b[155])^(a[149] & b[156])^(a[148] & b[157])^(a[147] & b[158])^(a[146] & b[159])^(a[145] & b[160])^(a[144] & b[161])^(a[143] & b[162])^(a[142] & b[163])^(a[141] & b[164])^(a[140] & b[165])^(a[139] & b[166])^(a[138] & b[167])^(a[137] & b[168])^(a[136] & b[169])^(a[135] & b[170])^(a[134] & b[171])^(a[133] & b[172])^(a[132] & b[173])^(a[131] & b[174])^(a[130] & b[175])^(a[129] & b[176])^(a[128] & b[177])^(a[127] & b[178])^(a[126] & b[179])^(a[125] & b[180])^(a[124] & b[181])^(a[123] & b[182])^(a[122] & b[183])^(a[121] & b[184])^(a[120] & b[185])^(a[119] & b[186])^(a[118] & b[187])^(a[117] & b[188])^(a[116] & b[189])^(a[115] & b[190])^(a[114] & b[191])^(a[113] & b[192])^(a[112] & b[193])^(a[111] & b[194])^(a[110] & b[195])^(a[109] & b[196])^(a[108] & b[197])^(a[107] & b[198])^(a[106] & b[199])^(a[105] & b[200])^(a[104] & b[201])^(a[103] & b[202])^(a[102] & b[203])^(a[101] & b[204])^(a[100] & b[205])^(a[99] & b[206])^(a[98] & b[207])^(a[97] & b[208])^(a[96] & b[209])^(a[95] & b[210])^(a[94] & b[211])^(a[93] & b[212])^(a[92] & b[213])^(a[91] & b[214])^(a[90] & b[215])^(a[89] & b[216])^(a[88] & b[217])^(a[87] & b[218])^(a[86] & b[219])^(a[85] & b[220])^(a[84] & b[221])^(a[83] & b[222])^(a[82] & b[223])^(a[81] & b[224])^(a[80] & b[225])^(a[79] & b[226])^(a[78] & b[227])^(a[77] & b[228])^(a[76] & b[229])^(a[75] & b[230])^(a[74] & b[231])^(a[73] & b[232]);
assign y[306] = (a[232] & b[74])^(a[231] & b[75])^(a[230] & b[76])^(a[229] & b[77])^(a[228] & b[78])^(a[227] & b[79])^(a[226] & b[80])^(a[225] & b[81])^(a[224] & b[82])^(a[223] & b[83])^(a[222] & b[84])^(a[221] & b[85])^(a[220] & b[86])^(a[219] & b[87])^(a[218] & b[88])^(a[217] & b[89])^(a[216] & b[90])^(a[215] & b[91])^(a[214] & b[92])^(a[213] & b[93])^(a[212] & b[94])^(a[211] & b[95])^(a[210] & b[96])^(a[209] & b[97])^(a[208] & b[98])^(a[207] & b[99])^(a[206] & b[100])^(a[205] & b[101])^(a[204] & b[102])^(a[203] & b[103])^(a[202] & b[104])^(a[201] & b[105])^(a[200] & b[106])^(a[199] & b[107])^(a[198] & b[108])^(a[197] & b[109])^(a[196] & b[110])^(a[195] & b[111])^(a[194] & b[112])^(a[193] & b[113])^(a[192] & b[114])^(a[191] & b[115])^(a[190] & b[116])^(a[189] & b[117])^(a[188] & b[118])^(a[187] & b[119])^(a[186] & b[120])^(a[185] & b[121])^(a[184] & b[122])^(a[183] & b[123])^(a[182] & b[124])^(a[181] & b[125])^(a[180] & b[126])^(a[179] & b[127])^(a[178] & b[128])^(a[177] & b[129])^(a[176] & b[130])^(a[175] & b[131])^(a[174] & b[132])^(a[173] & b[133])^(a[172] & b[134])^(a[171] & b[135])^(a[170] & b[136])^(a[169] & b[137])^(a[168] & b[138])^(a[167] & b[139])^(a[166] & b[140])^(a[165] & b[141])^(a[164] & b[142])^(a[163] & b[143])^(a[162] & b[144])^(a[161] & b[145])^(a[160] & b[146])^(a[159] & b[147])^(a[158] & b[148])^(a[157] & b[149])^(a[156] & b[150])^(a[155] & b[151])^(a[154] & b[152])^(a[153] & b[153])^(a[152] & b[154])^(a[151] & b[155])^(a[150] & b[156])^(a[149] & b[157])^(a[148] & b[158])^(a[147] & b[159])^(a[146] & b[160])^(a[145] & b[161])^(a[144] & b[162])^(a[143] & b[163])^(a[142] & b[164])^(a[141] & b[165])^(a[140] & b[166])^(a[139] & b[167])^(a[138] & b[168])^(a[137] & b[169])^(a[136] & b[170])^(a[135] & b[171])^(a[134] & b[172])^(a[133] & b[173])^(a[132] & b[174])^(a[131] & b[175])^(a[130] & b[176])^(a[129] & b[177])^(a[128] & b[178])^(a[127] & b[179])^(a[126] & b[180])^(a[125] & b[181])^(a[124] & b[182])^(a[123] & b[183])^(a[122] & b[184])^(a[121] & b[185])^(a[120] & b[186])^(a[119] & b[187])^(a[118] & b[188])^(a[117] & b[189])^(a[116] & b[190])^(a[115] & b[191])^(a[114] & b[192])^(a[113] & b[193])^(a[112] & b[194])^(a[111] & b[195])^(a[110] & b[196])^(a[109] & b[197])^(a[108] & b[198])^(a[107] & b[199])^(a[106] & b[200])^(a[105] & b[201])^(a[104] & b[202])^(a[103] & b[203])^(a[102] & b[204])^(a[101] & b[205])^(a[100] & b[206])^(a[99] & b[207])^(a[98] & b[208])^(a[97] & b[209])^(a[96] & b[210])^(a[95] & b[211])^(a[94] & b[212])^(a[93] & b[213])^(a[92] & b[214])^(a[91] & b[215])^(a[90] & b[216])^(a[89] & b[217])^(a[88] & b[218])^(a[87] & b[219])^(a[86] & b[220])^(a[85] & b[221])^(a[84] & b[222])^(a[83] & b[223])^(a[82] & b[224])^(a[81] & b[225])^(a[80] & b[226])^(a[79] & b[227])^(a[78] & b[228])^(a[77] & b[229])^(a[76] & b[230])^(a[75] & b[231])^(a[74] & b[232]);
assign y[307] = (a[232] & b[75])^(a[231] & b[76])^(a[230] & b[77])^(a[229] & b[78])^(a[228] & b[79])^(a[227] & b[80])^(a[226] & b[81])^(a[225] & b[82])^(a[224] & b[83])^(a[223] & b[84])^(a[222] & b[85])^(a[221] & b[86])^(a[220] & b[87])^(a[219] & b[88])^(a[218] & b[89])^(a[217] & b[90])^(a[216] & b[91])^(a[215] & b[92])^(a[214] & b[93])^(a[213] & b[94])^(a[212] & b[95])^(a[211] & b[96])^(a[210] & b[97])^(a[209] & b[98])^(a[208] & b[99])^(a[207] & b[100])^(a[206] & b[101])^(a[205] & b[102])^(a[204] & b[103])^(a[203] & b[104])^(a[202] & b[105])^(a[201] & b[106])^(a[200] & b[107])^(a[199] & b[108])^(a[198] & b[109])^(a[197] & b[110])^(a[196] & b[111])^(a[195] & b[112])^(a[194] & b[113])^(a[193] & b[114])^(a[192] & b[115])^(a[191] & b[116])^(a[190] & b[117])^(a[189] & b[118])^(a[188] & b[119])^(a[187] & b[120])^(a[186] & b[121])^(a[185] & b[122])^(a[184] & b[123])^(a[183] & b[124])^(a[182] & b[125])^(a[181] & b[126])^(a[180] & b[127])^(a[179] & b[128])^(a[178] & b[129])^(a[177] & b[130])^(a[176] & b[131])^(a[175] & b[132])^(a[174] & b[133])^(a[173] & b[134])^(a[172] & b[135])^(a[171] & b[136])^(a[170] & b[137])^(a[169] & b[138])^(a[168] & b[139])^(a[167] & b[140])^(a[166] & b[141])^(a[165] & b[142])^(a[164] & b[143])^(a[163] & b[144])^(a[162] & b[145])^(a[161] & b[146])^(a[160] & b[147])^(a[159] & b[148])^(a[158] & b[149])^(a[157] & b[150])^(a[156] & b[151])^(a[155] & b[152])^(a[154] & b[153])^(a[153] & b[154])^(a[152] & b[155])^(a[151] & b[156])^(a[150] & b[157])^(a[149] & b[158])^(a[148] & b[159])^(a[147] & b[160])^(a[146] & b[161])^(a[145] & b[162])^(a[144] & b[163])^(a[143] & b[164])^(a[142] & b[165])^(a[141] & b[166])^(a[140] & b[167])^(a[139] & b[168])^(a[138] & b[169])^(a[137] & b[170])^(a[136] & b[171])^(a[135] & b[172])^(a[134] & b[173])^(a[133] & b[174])^(a[132] & b[175])^(a[131] & b[176])^(a[130] & b[177])^(a[129] & b[178])^(a[128] & b[179])^(a[127] & b[180])^(a[126] & b[181])^(a[125] & b[182])^(a[124] & b[183])^(a[123] & b[184])^(a[122] & b[185])^(a[121] & b[186])^(a[120] & b[187])^(a[119] & b[188])^(a[118] & b[189])^(a[117] & b[190])^(a[116] & b[191])^(a[115] & b[192])^(a[114] & b[193])^(a[113] & b[194])^(a[112] & b[195])^(a[111] & b[196])^(a[110] & b[197])^(a[109] & b[198])^(a[108] & b[199])^(a[107] & b[200])^(a[106] & b[201])^(a[105] & b[202])^(a[104] & b[203])^(a[103] & b[204])^(a[102] & b[205])^(a[101] & b[206])^(a[100] & b[207])^(a[99] & b[208])^(a[98] & b[209])^(a[97] & b[210])^(a[96] & b[211])^(a[95] & b[212])^(a[94] & b[213])^(a[93] & b[214])^(a[92] & b[215])^(a[91] & b[216])^(a[90] & b[217])^(a[89] & b[218])^(a[88] & b[219])^(a[87] & b[220])^(a[86] & b[221])^(a[85] & b[222])^(a[84] & b[223])^(a[83] & b[224])^(a[82] & b[225])^(a[81] & b[226])^(a[80] & b[227])^(a[79] & b[228])^(a[78] & b[229])^(a[77] & b[230])^(a[76] & b[231])^(a[75] & b[232]);
assign y[308] = (a[232] & b[76])^(a[231] & b[77])^(a[230] & b[78])^(a[229] & b[79])^(a[228] & b[80])^(a[227] & b[81])^(a[226] & b[82])^(a[225] & b[83])^(a[224] & b[84])^(a[223] & b[85])^(a[222] & b[86])^(a[221] & b[87])^(a[220] & b[88])^(a[219] & b[89])^(a[218] & b[90])^(a[217] & b[91])^(a[216] & b[92])^(a[215] & b[93])^(a[214] & b[94])^(a[213] & b[95])^(a[212] & b[96])^(a[211] & b[97])^(a[210] & b[98])^(a[209] & b[99])^(a[208] & b[100])^(a[207] & b[101])^(a[206] & b[102])^(a[205] & b[103])^(a[204] & b[104])^(a[203] & b[105])^(a[202] & b[106])^(a[201] & b[107])^(a[200] & b[108])^(a[199] & b[109])^(a[198] & b[110])^(a[197] & b[111])^(a[196] & b[112])^(a[195] & b[113])^(a[194] & b[114])^(a[193] & b[115])^(a[192] & b[116])^(a[191] & b[117])^(a[190] & b[118])^(a[189] & b[119])^(a[188] & b[120])^(a[187] & b[121])^(a[186] & b[122])^(a[185] & b[123])^(a[184] & b[124])^(a[183] & b[125])^(a[182] & b[126])^(a[181] & b[127])^(a[180] & b[128])^(a[179] & b[129])^(a[178] & b[130])^(a[177] & b[131])^(a[176] & b[132])^(a[175] & b[133])^(a[174] & b[134])^(a[173] & b[135])^(a[172] & b[136])^(a[171] & b[137])^(a[170] & b[138])^(a[169] & b[139])^(a[168] & b[140])^(a[167] & b[141])^(a[166] & b[142])^(a[165] & b[143])^(a[164] & b[144])^(a[163] & b[145])^(a[162] & b[146])^(a[161] & b[147])^(a[160] & b[148])^(a[159] & b[149])^(a[158] & b[150])^(a[157] & b[151])^(a[156] & b[152])^(a[155] & b[153])^(a[154] & b[154])^(a[153] & b[155])^(a[152] & b[156])^(a[151] & b[157])^(a[150] & b[158])^(a[149] & b[159])^(a[148] & b[160])^(a[147] & b[161])^(a[146] & b[162])^(a[145] & b[163])^(a[144] & b[164])^(a[143] & b[165])^(a[142] & b[166])^(a[141] & b[167])^(a[140] & b[168])^(a[139] & b[169])^(a[138] & b[170])^(a[137] & b[171])^(a[136] & b[172])^(a[135] & b[173])^(a[134] & b[174])^(a[133] & b[175])^(a[132] & b[176])^(a[131] & b[177])^(a[130] & b[178])^(a[129] & b[179])^(a[128] & b[180])^(a[127] & b[181])^(a[126] & b[182])^(a[125] & b[183])^(a[124] & b[184])^(a[123] & b[185])^(a[122] & b[186])^(a[121] & b[187])^(a[120] & b[188])^(a[119] & b[189])^(a[118] & b[190])^(a[117] & b[191])^(a[116] & b[192])^(a[115] & b[193])^(a[114] & b[194])^(a[113] & b[195])^(a[112] & b[196])^(a[111] & b[197])^(a[110] & b[198])^(a[109] & b[199])^(a[108] & b[200])^(a[107] & b[201])^(a[106] & b[202])^(a[105] & b[203])^(a[104] & b[204])^(a[103] & b[205])^(a[102] & b[206])^(a[101] & b[207])^(a[100] & b[208])^(a[99] & b[209])^(a[98] & b[210])^(a[97] & b[211])^(a[96] & b[212])^(a[95] & b[213])^(a[94] & b[214])^(a[93] & b[215])^(a[92] & b[216])^(a[91] & b[217])^(a[90] & b[218])^(a[89] & b[219])^(a[88] & b[220])^(a[87] & b[221])^(a[86] & b[222])^(a[85] & b[223])^(a[84] & b[224])^(a[83] & b[225])^(a[82] & b[226])^(a[81] & b[227])^(a[80] & b[228])^(a[79] & b[229])^(a[78] & b[230])^(a[77] & b[231])^(a[76] & b[232]);
assign y[309] = (a[232] & b[77])^(a[231] & b[78])^(a[230] & b[79])^(a[229] & b[80])^(a[228] & b[81])^(a[227] & b[82])^(a[226] & b[83])^(a[225] & b[84])^(a[224] & b[85])^(a[223] & b[86])^(a[222] & b[87])^(a[221] & b[88])^(a[220] & b[89])^(a[219] & b[90])^(a[218] & b[91])^(a[217] & b[92])^(a[216] & b[93])^(a[215] & b[94])^(a[214] & b[95])^(a[213] & b[96])^(a[212] & b[97])^(a[211] & b[98])^(a[210] & b[99])^(a[209] & b[100])^(a[208] & b[101])^(a[207] & b[102])^(a[206] & b[103])^(a[205] & b[104])^(a[204] & b[105])^(a[203] & b[106])^(a[202] & b[107])^(a[201] & b[108])^(a[200] & b[109])^(a[199] & b[110])^(a[198] & b[111])^(a[197] & b[112])^(a[196] & b[113])^(a[195] & b[114])^(a[194] & b[115])^(a[193] & b[116])^(a[192] & b[117])^(a[191] & b[118])^(a[190] & b[119])^(a[189] & b[120])^(a[188] & b[121])^(a[187] & b[122])^(a[186] & b[123])^(a[185] & b[124])^(a[184] & b[125])^(a[183] & b[126])^(a[182] & b[127])^(a[181] & b[128])^(a[180] & b[129])^(a[179] & b[130])^(a[178] & b[131])^(a[177] & b[132])^(a[176] & b[133])^(a[175] & b[134])^(a[174] & b[135])^(a[173] & b[136])^(a[172] & b[137])^(a[171] & b[138])^(a[170] & b[139])^(a[169] & b[140])^(a[168] & b[141])^(a[167] & b[142])^(a[166] & b[143])^(a[165] & b[144])^(a[164] & b[145])^(a[163] & b[146])^(a[162] & b[147])^(a[161] & b[148])^(a[160] & b[149])^(a[159] & b[150])^(a[158] & b[151])^(a[157] & b[152])^(a[156] & b[153])^(a[155] & b[154])^(a[154] & b[155])^(a[153] & b[156])^(a[152] & b[157])^(a[151] & b[158])^(a[150] & b[159])^(a[149] & b[160])^(a[148] & b[161])^(a[147] & b[162])^(a[146] & b[163])^(a[145] & b[164])^(a[144] & b[165])^(a[143] & b[166])^(a[142] & b[167])^(a[141] & b[168])^(a[140] & b[169])^(a[139] & b[170])^(a[138] & b[171])^(a[137] & b[172])^(a[136] & b[173])^(a[135] & b[174])^(a[134] & b[175])^(a[133] & b[176])^(a[132] & b[177])^(a[131] & b[178])^(a[130] & b[179])^(a[129] & b[180])^(a[128] & b[181])^(a[127] & b[182])^(a[126] & b[183])^(a[125] & b[184])^(a[124] & b[185])^(a[123] & b[186])^(a[122] & b[187])^(a[121] & b[188])^(a[120] & b[189])^(a[119] & b[190])^(a[118] & b[191])^(a[117] & b[192])^(a[116] & b[193])^(a[115] & b[194])^(a[114] & b[195])^(a[113] & b[196])^(a[112] & b[197])^(a[111] & b[198])^(a[110] & b[199])^(a[109] & b[200])^(a[108] & b[201])^(a[107] & b[202])^(a[106] & b[203])^(a[105] & b[204])^(a[104] & b[205])^(a[103] & b[206])^(a[102] & b[207])^(a[101] & b[208])^(a[100] & b[209])^(a[99] & b[210])^(a[98] & b[211])^(a[97] & b[212])^(a[96] & b[213])^(a[95] & b[214])^(a[94] & b[215])^(a[93] & b[216])^(a[92] & b[217])^(a[91] & b[218])^(a[90] & b[219])^(a[89] & b[220])^(a[88] & b[221])^(a[87] & b[222])^(a[86] & b[223])^(a[85] & b[224])^(a[84] & b[225])^(a[83] & b[226])^(a[82] & b[227])^(a[81] & b[228])^(a[80] & b[229])^(a[79] & b[230])^(a[78] & b[231])^(a[77] & b[232]);
assign y[310] = (a[232] & b[78])^(a[231] & b[79])^(a[230] & b[80])^(a[229] & b[81])^(a[228] & b[82])^(a[227] & b[83])^(a[226] & b[84])^(a[225] & b[85])^(a[224] & b[86])^(a[223] & b[87])^(a[222] & b[88])^(a[221] & b[89])^(a[220] & b[90])^(a[219] & b[91])^(a[218] & b[92])^(a[217] & b[93])^(a[216] & b[94])^(a[215] & b[95])^(a[214] & b[96])^(a[213] & b[97])^(a[212] & b[98])^(a[211] & b[99])^(a[210] & b[100])^(a[209] & b[101])^(a[208] & b[102])^(a[207] & b[103])^(a[206] & b[104])^(a[205] & b[105])^(a[204] & b[106])^(a[203] & b[107])^(a[202] & b[108])^(a[201] & b[109])^(a[200] & b[110])^(a[199] & b[111])^(a[198] & b[112])^(a[197] & b[113])^(a[196] & b[114])^(a[195] & b[115])^(a[194] & b[116])^(a[193] & b[117])^(a[192] & b[118])^(a[191] & b[119])^(a[190] & b[120])^(a[189] & b[121])^(a[188] & b[122])^(a[187] & b[123])^(a[186] & b[124])^(a[185] & b[125])^(a[184] & b[126])^(a[183] & b[127])^(a[182] & b[128])^(a[181] & b[129])^(a[180] & b[130])^(a[179] & b[131])^(a[178] & b[132])^(a[177] & b[133])^(a[176] & b[134])^(a[175] & b[135])^(a[174] & b[136])^(a[173] & b[137])^(a[172] & b[138])^(a[171] & b[139])^(a[170] & b[140])^(a[169] & b[141])^(a[168] & b[142])^(a[167] & b[143])^(a[166] & b[144])^(a[165] & b[145])^(a[164] & b[146])^(a[163] & b[147])^(a[162] & b[148])^(a[161] & b[149])^(a[160] & b[150])^(a[159] & b[151])^(a[158] & b[152])^(a[157] & b[153])^(a[156] & b[154])^(a[155] & b[155])^(a[154] & b[156])^(a[153] & b[157])^(a[152] & b[158])^(a[151] & b[159])^(a[150] & b[160])^(a[149] & b[161])^(a[148] & b[162])^(a[147] & b[163])^(a[146] & b[164])^(a[145] & b[165])^(a[144] & b[166])^(a[143] & b[167])^(a[142] & b[168])^(a[141] & b[169])^(a[140] & b[170])^(a[139] & b[171])^(a[138] & b[172])^(a[137] & b[173])^(a[136] & b[174])^(a[135] & b[175])^(a[134] & b[176])^(a[133] & b[177])^(a[132] & b[178])^(a[131] & b[179])^(a[130] & b[180])^(a[129] & b[181])^(a[128] & b[182])^(a[127] & b[183])^(a[126] & b[184])^(a[125] & b[185])^(a[124] & b[186])^(a[123] & b[187])^(a[122] & b[188])^(a[121] & b[189])^(a[120] & b[190])^(a[119] & b[191])^(a[118] & b[192])^(a[117] & b[193])^(a[116] & b[194])^(a[115] & b[195])^(a[114] & b[196])^(a[113] & b[197])^(a[112] & b[198])^(a[111] & b[199])^(a[110] & b[200])^(a[109] & b[201])^(a[108] & b[202])^(a[107] & b[203])^(a[106] & b[204])^(a[105] & b[205])^(a[104] & b[206])^(a[103] & b[207])^(a[102] & b[208])^(a[101] & b[209])^(a[100] & b[210])^(a[99] & b[211])^(a[98] & b[212])^(a[97] & b[213])^(a[96] & b[214])^(a[95] & b[215])^(a[94] & b[216])^(a[93] & b[217])^(a[92] & b[218])^(a[91] & b[219])^(a[90] & b[220])^(a[89] & b[221])^(a[88] & b[222])^(a[87] & b[223])^(a[86] & b[224])^(a[85] & b[225])^(a[84] & b[226])^(a[83] & b[227])^(a[82] & b[228])^(a[81] & b[229])^(a[80] & b[230])^(a[79] & b[231])^(a[78] & b[232]);
assign y[311] = (a[232] & b[79])^(a[231] & b[80])^(a[230] & b[81])^(a[229] & b[82])^(a[228] & b[83])^(a[227] & b[84])^(a[226] & b[85])^(a[225] & b[86])^(a[224] & b[87])^(a[223] & b[88])^(a[222] & b[89])^(a[221] & b[90])^(a[220] & b[91])^(a[219] & b[92])^(a[218] & b[93])^(a[217] & b[94])^(a[216] & b[95])^(a[215] & b[96])^(a[214] & b[97])^(a[213] & b[98])^(a[212] & b[99])^(a[211] & b[100])^(a[210] & b[101])^(a[209] & b[102])^(a[208] & b[103])^(a[207] & b[104])^(a[206] & b[105])^(a[205] & b[106])^(a[204] & b[107])^(a[203] & b[108])^(a[202] & b[109])^(a[201] & b[110])^(a[200] & b[111])^(a[199] & b[112])^(a[198] & b[113])^(a[197] & b[114])^(a[196] & b[115])^(a[195] & b[116])^(a[194] & b[117])^(a[193] & b[118])^(a[192] & b[119])^(a[191] & b[120])^(a[190] & b[121])^(a[189] & b[122])^(a[188] & b[123])^(a[187] & b[124])^(a[186] & b[125])^(a[185] & b[126])^(a[184] & b[127])^(a[183] & b[128])^(a[182] & b[129])^(a[181] & b[130])^(a[180] & b[131])^(a[179] & b[132])^(a[178] & b[133])^(a[177] & b[134])^(a[176] & b[135])^(a[175] & b[136])^(a[174] & b[137])^(a[173] & b[138])^(a[172] & b[139])^(a[171] & b[140])^(a[170] & b[141])^(a[169] & b[142])^(a[168] & b[143])^(a[167] & b[144])^(a[166] & b[145])^(a[165] & b[146])^(a[164] & b[147])^(a[163] & b[148])^(a[162] & b[149])^(a[161] & b[150])^(a[160] & b[151])^(a[159] & b[152])^(a[158] & b[153])^(a[157] & b[154])^(a[156] & b[155])^(a[155] & b[156])^(a[154] & b[157])^(a[153] & b[158])^(a[152] & b[159])^(a[151] & b[160])^(a[150] & b[161])^(a[149] & b[162])^(a[148] & b[163])^(a[147] & b[164])^(a[146] & b[165])^(a[145] & b[166])^(a[144] & b[167])^(a[143] & b[168])^(a[142] & b[169])^(a[141] & b[170])^(a[140] & b[171])^(a[139] & b[172])^(a[138] & b[173])^(a[137] & b[174])^(a[136] & b[175])^(a[135] & b[176])^(a[134] & b[177])^(a[133] & b[178])^(a[132] & b[179])^(a[131] & b[180])^(a[130] & b[181])^(a[129] & b[182])^(a[128] & b[183])^(a[127] & b[184])^(a[126] & b[185])^(a[125] & b[186])^(a[124] & b[187])^(a[123] & b[188])^(a[122] & b[189])^(a[121] & b[190])^(a[120] & b[191])^(a[119] & b[192])^(a[118] & b[193])^(a[117] & b[194])^(a[116] & b[195])^(a[115] & b[196])^(a[114] & b[197])^(a[113] & b[198])^(a[112] & b[199])^(a[111] & b[200])^(a[110] & b[201])^(a[109] & b[202])^(a[108] & b[203])^(a[107] & b[204])^(a[106] & b[205])^(a[105] & b[206])^(a[104] & b[207])^(a[103] & b[208])^(a[102] & b[209])^(a[101] & b[210])^(a[100] & b[211])^(a[99] & b[212])^(a[98] & b[213])^(a[97] & b[214])^(a[96] & b[215])^(a[95] & b[216])^(a[94] & b[217])^(a[93] & b[218])^(a[92] & b[219])^(a[91] & b[220])^(a[90] & b[221])^(a[89] & b[222])^(a[88] & b[223])^(a[87] & b[224])^(a[86] & b[225])^(a[85] & b[226])^(a[84] & b[227])^(a[83] & b[228])^(a[82] & b[229])^(a[81] & b[230])^(a[80] & b[231])^(a[79] & b[232]);
assign y[312] = (a[232] & b[80])^(a[231] & b[81])^(a[230] & b[82])^(a[229] & b[83])^(a[228] & b[84])^(a[227] & b[85])^(a[226] & b[86])^(a[225] & b[87])^(a[224] & b[88])^(a[223] & b[89])^(a[222] & b[90])^(a[221] & b[91])^(a[220] & b[92])^(a[219] & b[93])^(a[218] & b[94])^(a[217] & b[95])^(a[216] & b[96])^(a[215] & b[97])^(a[214] & b[98])^(a[213] & b[99])^(a[212] & b[100])^(a[211] & b[101])^(a[210] & b[102])^(a[209] & b[103])^(a[208] & b[104])^(a[207] & b[105])^(a[206] & b[106])^(a[205] & b[107])^(a[204] & b[108])^(a[203] & b[109])^(a[202] & b[110])^(a[201] & b[111])^(a[200] & b[112])^(a[199] & b[113])^(a[198] & b[114])^(a[197] & b[115])^(a[196] & b[116])^(a[195] & b[117])^(a[194] & b[118])^(a[193] & b[119])^(a[192] & b[120])^(a[191] & b[121])^(a[190] & b[122])^(a[189] & b[123])^(a[188] & b[124])^(a[187] & b[125])^(a[186] & b[126])^(a[185] & b[127])^(a[184] & b[128])^(a[183] & b[129])^(a[182] & b[130])^(a[181] & b[131])^(a[180] & b[132])^(a[179] & b[133])^(a[178] & b[134])^(a[177] & b[135])^(a[176] & b[136])^(a[175] & b[137])^(a[174] & b[138])^(a[173] & b[139])^(a[172] & b[140])^(a[171] & b[141])^(a[170] & b[142])^(a[169] & b[143])^(a[168] & b[144])^(a[167] & b[145])^(a[166] & b[146])^(a[165] & b[147])^(a[164] & b[148])^(a[163] & b[149])^(a[162] & b[150])^(a[161] & b[151])^(a[160] & b[152])^(a[159] & b[153])^(a[158] & b[154])^(a[157] & b[155])^(a[156] & b[156])^(a[155] & b[157])^(a[154] & b[158])^(a[153] & b[159])^(a[152] & b[160])^(a[151] & b[161])^(a[150] & b[162])^(a[149] & b[163])^(a[148] & b[164])^(a[147] & b[165])^(a[146] & b[166])^(a[145] & b[167])^(a[144] & b[168])^(a[143] & b[169])^(a[142] & b[170])^(a[141] & b[171])^(a[140] & b[172])^(a[139] & b[173])^(a[138] & b[174])^(a[137] & b[175])^(a[136] & b[176])^(a[135] & b[177])^(a[134] & b[178])^(a[133] & b[179])^(a[132] & b[180])^(a[131] & b[181])^(a[130] & b[182])^(a[129] & b[183])^(a[128] & b[184])^(a[127] & b[185])^(a[126] & b[186])^(a[125] & b[187])^(a[124] & b[188])^(a[123] & b[189])^(a[122] & b[190])^(a[121] & b[191])^(a[120] & b[192])^(a[119] & b[193])^(a[118] & b[194])^(a[117] & b[195])^(a[116] & b[196])^(a[115] & b[197])^(a[114] & b[198])^(a[113] & b[199])^(a[112] & b[200])^(a[111] & b[201])^(a[110] & b[202])^(a[109] & b[203])^(a[108] & b[204])^(a[107] & b[205])^(a[106] & b[206])^(a[105] & b[207])^(a[104] & b[208])^(a[103] & b[209])^(a[102] & b[210])^(a[101] & b[211])^(a[100] & b[212])^(a[99] & b[213])^(a[98] & b[214])^(a[97] & b[215])^(a[96] & b[216])^(a[95] & b[217])^(a[94] & b[218])^(a[93] & b[219])^(a[92] & b[220])^(a[91] & b[221])^(a[90] & b[222])^(a[89] & b[223])^(a[88] & b[224])^(a[87] & b[225])^(a[86] & b[226])^(a[85] & b[227])^(a[84] & b[228])^(a[83] & b[229])^(a[82] & b[230])^(a[81] & b[231])^(a[80] & b[232]);
assign y[313] = (a[232] & b[81])^(a[231] & b[82])^(a[230] & b[83])^(a[229] & b[84])^(a[228] & b[85])^(a[227] & b[86])^(a[226] & b[87])^(a[225] & b[88])^(a[224] & b[89])^(a[223] & b[90])^(a[222] & b[91])^(a[221] & b[92])^(a[220] & b[93])^(a[219] & b[94])^(a[218] & b[95])^(a[217] & b[96])^(a[216] & b[97])^(a[215] & b[98])^(a[214] & b[99])^(a[213] & b[100])^(a[212] & b[101])^(a[211] & b[102])^(a[210] & b[103])^(a[209] & b[104])^(a[208] & b[105])^(a[207] & b[106])^(a[206] & b[107])^(a[205] & b[108])^(a[204] & b[109])^(a[203] & b[110])^(a[202] & b[111])^(a[201] & b[112])^(a[200] & b[113])^(a[199] & b[114])^(a[198] & b[115])^(a[197] & b[116])^(a[196] & b[117])^(a[195] & b[118])^(a[194] & b[119])^(a[193] & b[120])^(a[192] & b[121])^(a[191] & b[122])^(a[190] & b[123])^(a[189] & b[124])^(a[188] & b[125])^(a[187] & b[126])^(a[186] & b[127])^(a[185] & b[128])^(a[184] & b[129])^(a[183] & b[130])^(a[182] & b[131])^(a[181] & b[132])^(a[180] & b[133])^(a[179] & b[134])^(a[178] & b[135])^(a[177] & b[136])^(a[176] & b[137])^(a[175] & b[138])^(a[174] & b[139])^(a[173] & b[140])^(a[172] & b[141])^(a[171] & b[142])^(a[170] & b[143])^(a[169] & b[144])^(a[168] & b[145])^(a[167] & b[146])^(a[166] & b[147])^(a[165] & b[148])^(a[164] & b[149])^(a[163] & b[150])^(a[162] & b[151])^(a[161] & b[152])^(a[160] & b[153])^(a[159] & b[154])^(a[158] & b[155])^(a[157] & b[156])^(a[156] & b[157])^(a[155] & b[158])^(a[154] & b[159])^(a[153] & b[160])^(a[152] & b[161])^(a[151] & b[162])^(a[150] & b[163])^(a[149] & b[164])^(a[148] & b[165])^(a[147] & b[166])^(a[146] & b[167])^(a[145] & b[168])^(a[144] & b[169])^(a[143] & b[170])^(a[142] & b[171])^(a[141] & b[172])^(a[140] & b[173])^(a[139] & b[174])^(a[138] & b[175])^(a[137] & b[176])^(a[136] & b[177])^(a[135] & b[178])^(a[134] & b[179])^(a[133] & b[180])^(a[132] & b[181])^(a[131] & b[182])^(a[130] & b[183])^(a[129] & b[184])^(a[128] & b[185])^(a[127] & b[186])^(a[126] & b[187])^(a[125] & b[188])^(a[124] & b[189])^(a[123] & b[190])^(a[122] & b[191])^(a[121] & b[192])^(a[120] & b[193])^(a[119] & b[194])^(a[118] & b[195])^(a[117] & b[196])^(a[116] & b[197])^(a[115] & b[198])^(a[114] & b[199])^(a[113] & b[200])^(a[112] & b[201])^(a[111] & b[202])^(a[110] & b[203])^(a[109] & b[204])^(a[108] & b[205])^(a[107] & b[206])^(a[106] & b[207])^(a[105] & b[208])^(a[104] & b[209])^(a[103] & b[210])^(a[102] & b[211])^(a[101] & b[212])^(a[100] & b[213])^(a[99] & b[214])^(a[98] & b[215])^(a[97] & b[216])^(a[96] & b[217])^(a[95] & b[218])^(a[94] & b[219])^(a[93] & b[220])^(a[92] & b[221])^(a[91] & b[222])^(a[90] & b[223])^(a[89] & b[224])^(a[88] & b[225])^(a[87] & b[226])^(a[86] & b[227])^(a[85] & b[228])^(a[84] & b[229])^(a[83] & b[230])^(a[82] & b[231])^(a[81] & b[232]);
assign y[314] = (a[232] & b[82])^(a[231] & b[83])^(a[230] & b[84])^(a[229] & b[85])^(a[228] & b[86])^(a[227] & b[87])^(a[226] & b[88])^(a[225] & b[89])^(a[224] & b[90])^(a[223] & b[91])^(a[222] & b[92])^(a[221] & b[93])^(a[220] & b[94])^(a[219] & b[95])^(a[218] & b[96])^(a[217] & b[97])^(a[216] & b[98])^(a[215] & b[99])^(a[214] & b[100])^(a[213] & b[101])^(a[212] & b[102])^(a[211] & b[103])^(a[210] & b[104])^(a[209] & b[105])^(a[208] & b[106])^(a[207] & b[107])^(a[206] & b[108])^(a[205] & b[109])^(a[204] & b[110])^(a[203] & b[111])^(a[202] & b[112])^(a[201] & b[113])^(a[200] & b[114])^(a[199] & b[115])^(a[198] & b[116])^(a[197] & b[117])^(a[196] & b[118])^(a[195] & b[119])^(a[194] & b[120])^(a[193] & b[121])^(a[192] & b[122])^(a[191] & b[123])^(a[190] & b[124])^(a[189] & b[125])^(a[188] & b[126])^(a[187] & b[127])^(a[186] & b[128])^(a[185] & b[129])^(a[184] & b[130])^(a[183] & b[131])^(a[182] & b[132])^(a[181] & b[133])^(a[180] & b[134])^(a[179] & b[135])^(a[178] & b[136])^(a[177] & b[137])^(a[176] & b[138])^(a[175] & b[139])^(a[174] & b[140])^(a[173] & b[141])^(a[172] & b[142])^(a[171] & b[143])^(a[170] & b[144])^(a[169] & b[145])^(a[168] & b[146])^(a[167] & b[147])^(a[166] & b[148])^(a[165] & b[149])^(a[164] & b[150])^(a[163] & b[151])^(a[162] & b[152])^(a[161] & b[153])^(a[160] & b[154])^(a[159] & b[155])^(a[158] & b[156])^(a[157] & b[157])^(a[156] & b[158])^(a[155] & b[159])^(a[154] & b[160])^(a[153] & b[161])^(a[152] & b[162])^(a[151] & b[163])^(a[150] & b[164])^(a[149] & b[165])^(a[148] & b[166])^(a[147] & b[167])^(a[146] & b[168])^(a[145] & b[169])^(a[144] & b[170])^(a[143] & b[171])^(a[142] & b[172])^(a[141] & b[173])^(a[140] & b[174])^(a[139] & b[175])^(a[138] & b[176])^(a[137] & b[177])^(a[136] & b[178])^(a[135] & b[179])^(a[134] & b[180])^(a[133] & b[181])^(a[132] & b[182])^(a[131] & b[183])^(a[130] & b[184])^(a[129] & b[185])^(a[128] & b[186])^(a[127] & b[187])^(a[126] & b[188])^(a[125] & b[189])^(a[124] & b[190])^(a[123] & b[191])^(a[122] & b[192])^(a[121] & b[193])^(a[120] & b[194])^(a[119] & b[195])^(a[118] & b[196])^(a[117] & b[197])^(a[116] & b[198])^(a[115] & b[199])^(a[114] & b[200])^(a[113] & b[201])^(a[112] & b[202])^(a[111] & b[203])^(a[110] & b[204])^(a[109] & b[205])^(a[108] & b[206])^(a[107] & b[207])^(a[106] & b[208])^(a[105] & b[209])^(a[104] & b[210])^(a[103] & b[211])^(a[102] & b[212])^(a[101] & b[213])^(a[100] & b[214])^(a[99] & b[215])^(a[98] & b[216])^(a[97] & b[217])^(a[96] & b[218])^(a[95] & b[219])^(a[94] & b[220])^(a[93] & b[221])^(a[92] & b[222])^(a[91] & b[223])^(a[90] & b[224])^(a[89] & b[225])^(a[88] & b[226])^(a[87] & b[227])^(a[86] & b[228])^(a[85] & b[229])^(a[84] & b[230])^(a[83] & b[231])^(a[82] & b[232]);
assign y[315] = (a[232] & b[83])^(a[231] & b[84])^(a[230] & b[85])^(a[229] & b[86])^(a[228] & b[87])^(a[227] & b[88])^(a[226] & b[89])^(a[225] & b[90])^(a[224] & b[91])^(a[223] & b[92])^(a[222] & b[93])^(a[221] & b[94])^(a[220] & b[95])^(a[219] & b[96])^(a[218] & b[97])^(a[217] & b[98])^(a[216] & b[99])^(a[215] & b[100])^(a[214] & b[101])^(a[213] & b[102])^(a[212] & b[103])^(a[211] & b[104])^(a[210] & b[105])^(a[209] & b[106])^(a[208] & b[107])^(a[207] & b[108])^(a[206] & b[109])^(a[205] & b[110])^(a[204] & b[111])^(a[203] & b[112])^(a[202] & b[113])^(a[201] & b[114])^(a[200] & b[115])^(a[199] & b[116])^(a[198] & b[117])^(a[197] & b[118])^(a[196] & b[119])^(a[195] & b[120])^(a[194] & b[121])^(a[193] & b[122])^(a[192] & b[123])^(a[191] & b[124])^(a[190] & b[125])^(a[189] & b[126])^(a[188] & b[127])^(a[187] & b[128])^(a[186] & b[129])^(a[185] & b[130])^(a[184] & b[131])^(a[183] & b[132])^(a[182] & b[133])^(a[181] & b[134])^(a[180] & b[135])^(a[179] & b[136])^(a[178] & b[137])^(a[177] & b[138])^(a[176] & b[139])^(a[175] & b[140])^(a[174] & b[141])^(a[173] & b[142])^(a[172] & b[143])^(a[171] & b[144])^(a[170] & b[145])^(a[169] & b[146])^(a[168] & b[147])^(a[167] & b[148])^(a[166] & b[149])^(a[165] & b[150])^(a[164] & b[151])^(a[163] & b[152])^(a[162] & b[153])^(a[161] & b[154])^(a[160] & b[155])^(a[159] & b[156])^(a[158] & b[157])^(a[157] & b[158])^(a[156] & b[159])^(a[155] & b[160])^(a[154] & b[161])^(a[153] & b[162])^(a[152] & b[163])^(a[151] & b[164])^(a[150] & b[165])^(a[149] & b[166])^(a[148] & b[167])^(a[147] & b[168])^(a[146] & b[169])^(a[145] & b[170])^(a[144] & b[171])^(a[143] & b[172])^(a[142] & b[173])^(a[141] & b[174])^(a[140] & b[175])^(a[139] & b[176])^(a[138] & b[177])^(a[137] & b[178])^(a[136] & b[179])^(a[135] & b[180])^(a[134] & b[181])^(a[133] & b[182])^(a[132] & b[183])^(a[131] & b[184])^(a[130] & b[185])^(a[129] & b[186])^(a[128] & b[187])^(a[127] & b[188])^(a[126] & b[189])^(a[125] & b[190])^(a[124] & b[191])^(a[123] & b[192])^(a[122] & b[193])^(a[121] & b[194])^(a[120] & b[195])^(a[119] & b[196])^(a[118] & b[197])^(a[117] & b[198])^(a[116] & b[199])^(a[115] & b[200])^(a[114] & b[201])^(a[113] & b[202])^(a[112] & b[203])^(a[111] & b[204])^(a[110] & b[205])^(a[109] & b[206])^(a[108] & b[207])^(a[107] & b[208])^(a[106] & b[209])^(a[105] & b[210])^(a[104] & b[211])^(a[103] & b[212])^(a[102] & b[213])^(a[101] & b[214])^(a[100] & b[215])^(a[99] & b[216])^(a[98] & b[217])^(a[97] & b[218])^(a[96] & b[219])^(a[95] & b[220])^(a[94] & b[221])^(a[93] & b[222])^(a[92] & b[223])^(a[91] & b[224])^(a[90] & b[225])^(a[89] & b[226])^(a[88] & b[227])^(a[87] & b[228])^(a[86] & b[229])^(a[85] & b[230])^(a[84] & b[231])^(a[83] & b[232]);
assign y[316] = (a[232] & b[84])^(a[231] & b[85])^(a[230] & b[86])^(a[229] & b[87])^(a[228] & b[88])^(a[227] & b[89])^(a[226] & b[90])^(a[225] & b[91])^(a[224] & b[92])^(a[223] & b[93])^(a[222] & b[94])^(a[221] & b[95])^(a[220] & b[96])^(a[219] & b[97])^(a[218] & b[98])^(a[217] & b[99])^(a[216] & b[100])^(a[215] & b[101])^(a[214] & b[102])^(a[213] & b[103])^(a[212] & b[104])^(a[211] & b[105])^(a[210] & b[106])^(a[209] & b[107])^(a[208] & b[108])^(a[207] & b[109])^(a[206] & b[110])^(a[205] & b[111])^(a[204] & b[112])^(a[203] & b[113])^(a[202] & b[114])^(a[201] & b[115])^(a[200] & b[116])^(a[199] & b[117])^(a[198] & b[118])^(a[197] & b[119])^(a[196] & b[120])^(a[195] & b[121])^(a[194] & b[122])^(a[193] & b[123])^(a[192] & b[124])^(a[191] & b[125])^(a[190] & b[126])^(a[189] & b[127])^(a[188] & b[128])^(a[187] & b[129])^(a[186] & b[130])^(a[185] & b[131])^(a[184] & b[132])^(a[183] & b[133])^(a[182] & b[134])^(a[181] & b[135])^(a[180] & b[136])^(a[179] & b[137])^(a[178] & b[138])^(a[177] & b[139])^(a[176] & b[140])^(a[175] & b[141])^(a[174] & b[142])^(a[173] & b[143])^(a[172] & b[144])^(a[171] & b[145])^(a[170] & b[146])^(a[169] & b[147])^(a[168] & b[148])^(a[167] & b[149])^(a[166] & b[150])^(a[165] & b[151])^(a[164] & b[152])^(a[163] & b[153])^(a[162] & b[154])^(a[161] & b[155])^(a[160] & b[156])^(a[159] & b[157])^(a[158] & b[158])^(a[157] & b[159])^(a[156] & b[160])^(a[155] & b[161])^(a[154] & b[162])^(a[153] & b[163])^(a[152] & b[164])^(a[151] & b[165])^(a[150] & b[166])^(a[149] & b[167])^(a[148] & b[168])^(a[147] & b[169])^(a[146] & b[170])^(a[145] & b[171])^(a[144] & b[172])^(a[143] & b[173])^(a[142] & b[174])^(a[141] & b[175])^(a[140] & b[176])^(a[139] & b[177])^(a[138] & b[178])^(a[137] & b[179])^(a[136] & b[180])^(a[135] & b[181])^(a[134] & b[182])^(a[133] & b[183])^(a[132] & b[184])^(a[131] & b[185])^(a[130] & b[186])^(a[129] & b[187])^(a[128] & b[188])^(a[127] & b[189])^(a[126] & b[190])^(a[125] & b[191])^(a[124] & b[192])^(a[123] & b[193])^(a[122] & b[194])^(a[121] & b[195])^(a[120] & b[196])^(a[119] & b[197])^(a[118] & b[198])^(a[117] & b[199])^(a[116] & b[200])^(a[115] & b[201])^(a[114] & b[202])^(a[113] & b[203])^(a[112] & b[204])^(a[111] & b[205])^(a[110] & b[206])^(a[109] & b[207])^(a[108] & b[208])^(a[107] & b[209])^(a[106] & b[210])^(a[105] & b[211])^(a[104] & b[212])^(a[103] & b[213])^(a[102] & b[214])^(a[101] & b[215])^(a[100] & b[216])^(a[99] & b[217])^(a[98] & b[218])^(a[97] & b[219])^(a[96] & b[220])^(a[95] & b[221])^(a[94] & b[222])^(a[93] & b[223])^(a[92] & b[224])^(a[91] & b[225])^(a[90] & b[226])^(a[89] & b[227])^(a[88] & b[228])^(a[87] & b[229])^(a[86] & b[230])^(a[85] & b[231])^(a[84] & b[232]);
assign y[317] = (a[232] & b[85])^(a[231] & b[86])^(a[230] & b[87])^(a[229] & b[88])^(a[228] & b[89])^(a[227] & b[90])^(a[226] & b[91])^(a[225] & b[92])^(a[224] & b[93])^(a[223] & b[94])^(a[222] & b[95])^(a[221] & b[96])^(a[220] & b[97])^(a[219] & b[98])^(a[218] & b[99])^(a[217] & b[100])^(a[216] & b[101])^(a[215] & b[102])^(a[214] & b[103])^(a[213] & b[104])^(a[212] & b[105])^(a[211] & b[106])^(a[210] & b[107])^(a[209] & b[108])^(a[208] & b[109])^(a[207] & b[110])^(a[206] & b[111])^(a[205] & b[112])^(a[204] & b[113])^(a[203] & b[114])^(a[202] & b[115])^(a[201] & b[116])^(a[200] & b[117])^(a[199] & b[118])^(a[198] & b[119])^(a[197] & b[120])^(a[196] & b[121])^(a[195] & b[122])^(a[194] & b[123])^(a[193] & b[124])^(a[192] & b[125])^(a[191] & b[126])^(a[190] & b[127])^(a[189] & b[128])^(a[188] & b[129])^(a[187] & b[130])^(a[186] & b[131])^(a[185] & b[132])^(a[184] & b[133])^(a[183] & b[134])^(a[182] & b[135])^(a[181] & b[136])^(a[180] & b[137])^(a[179] & b[138])^(a[178] & b[139])^(a[177] & b[140])^(a[176] & b[141])^(a[175] & b[142])^(a[174] & b[143])^(a[173] & b[144])^(a[172] & b[145])^(a[171] & b[146])^(a[170] & b[147])^(a[169] & b[148])^(a[168] & b[149])^(a[167] & b[150])^(a[166] & b[151])^(a[165] & b[152])^(a[164] & b[153])^(a[163] & b[154])^(a[162] & b[155])^(a[161] & b[156])^(a[160] & b[157])^(a[159] & b[158])^(a[158] & b[159])^(a[157] & b[160])^(a[156] & b[161])^(a[155] & b[162])^(a[154] & b[163])^(a[153] & b[164])^(a[152] & b[165])^(a[151] & b[166])^(a[150] & b[167])^(a[149] & b[168])^(a[148] & b[169])^(a[147] & b[170])^(a[146] & b[171])^(a[145] & b[172])^(a[144] & b[173])^(a[143] & b[174])^(a[142] & b[175])^(a[141] & b[176])^(a[140] & b[177])^(a[139] & b[178])^(a[138] & b[179])^(a[137] & b[180])^(a[136] & b[181])^(a[135] & b[182])^(a[134] & b[183])^(a[133] & b[184])^(a[132] & b[185])^(a[131] & b[186])^(a[130] & b[187])^(a[129] & b[188])^(a[128] & b[189])^(a[127] & b[190])^(a[126] & b[191])^(a[125] & b[192])^(a[124] & b[193])^(a[123] & b[194])^(a[122] & b[195])^(a[121] & b[196])^(a[120] & b[197])^(a[119] & b[198])^(a[118] & b[199])^(a[117] & b[200])^(a[116] & b[201])^(a[115] & b[202])^(a[114] & b[203])^(a[113] & b[204])^(a[112] & b[205])^(a[111] & b[206])^(a[110] & b[207])^(a[109] & b[208])^(a[108] & b[209])^(a[107] & b[210])^(a[106] & b[211])^(a[105] & b[212])^(a[104] & b[213])^(a[103] & b[214])^(a[102] & b[215])^(a[101] & b[216])^(a[100] & b[217])^(a[99] & b[218])^(a[98] & b[219])^(a[97] & b[220])^(a[96] & b[221])^(a[95] & b[222])^(a[94] & b[223])^(a[93] & b[224])^(a[92] & b[225])^(a[91] & b[226])^(a[90] & b[227])^(a[89] & b[228])^(a[88] & b[229])^(a[87] & b[230])^(a[86] & b[231])^(a[85] & b[232]);
assign y[318] = (a[232] & b[86])^(a[231] & b[87])^(a[230] & b[88])^(a[229] & b[89])^(a[228] & b[90])^(a[227] & b[91])^(a[226] & b[92])^(a[225] & b[93])^(a[224] & b[94])^(a[223] & b[95])^(a[222] & b[96])^(a[221] & b[97])^(a[220] & b[98])^(a[219] & b[99])^(a[218] & b[100])^(a[217] & b[101])^(a[216] & b[102])^(a[215] & b[103])^(a[214] & b[104])^(a[213] & b[105])^(a[212] & b[106])^(a[211] & b[107])^(a[210] & b[108])^(a[209] & b[109])^(a[208] & b[110])^(a[207] & b[111])^(a[206] & b[112])^(a[205] & b[113])^(a[204] & b[114])^(a[203] & b[115])^(a[202] & b[116])^(a[201] & b[117])^(a[200] & b[118])^(a[199] & b[119])^(a[198] & b[120])^(a[197] & b[121])^(a[196] & b[122])^(a[195] & b[123])^(a[194] & b[124])^(a[193] & b[125])^(a[192] & b[126])^(a[191] & b[127])^(a[190] & b[128])^(a[189] & b[129])^(a[188] & b[130])^(a[187] & b[131])^(a[186] & b[132])^(a[185] & b[133])^(a[184] & b[134])^(a[183] & b[135])^(a[182] & b[136])^(a[181] & b[137])^(a[180] & b[138])^(a[179] & b[139])^(a[178] & b[140])^(a[177] & b[141])^(a[176] & b[142])^(a[175] & b[143])^(a[174] & b[144])^(a[173] & b[145])^(a[172] & b[146])^(a[171] & b[147])^(a[170] & b[148])^(a[169] & b[149])^(a[168] & b[150])^(a[167] & b[151])^(a[166] & b[152])^(a[165] & b[153])^(a[164] & b[154])^(a[163] & b[155])^(a[162] & b[156])^(a[161] & b[157])^(a[160] & b[158])^(a[159] & b[159])^(a[158] & b[160])^(a[157] & b[161])^(a[156] & b[162])^(a[155] & b[163])^(a[154] & b[164])^(a[153] & b[165])^(a[152] & b[166])^(a[151] & b[167])^(a[150] & b[168])^(a[149] & b[169])^(a[148] & b[170])^(a[147] & b[171])^(a[146] & b[172])^(a[145] & b[173])^(a[144] & b[174])^(a[143] & b[175])^(a[142] & b[176])^(a[141] & b[177])^(a[140] & b[178])^(a[139] & b[179])^(a[138] & b[180])^(a[137] & b[181])^(a[136] & b[182])^(a[135] & b[183])^(a[134] & b[184])^(a[133] & b[185])^(a[132] & b[186])^(a[131] & b[187])^(a[130] & b[188])^(a[129] & b[189])^(a[128] & b[190])^(a[127] & b[191])^(a[126] & b[192])^(a[125] & b[193])^(a[124] & b[194])^(a[123] & b[195])^(a[122] & b[196])^(a[121] & b[197])^(a[120] & b[198])^(a[119] & b[199])^(a[118] & b[200])^(a[117] & b[201])^(a[116] & b[202])^(a[115] & b[203])^(a[114] & b[204])^(a[113] & b[205])^(a[112] & b[206])^(a[111] & b[207])^(a[110] & b[208])^(a[109] & b[209])^(a[108] & b[210])^(a[107] & b[211])^(a[106] & b[212])^(a[105] & b[213])^(a[104] & b[214])^(a[103] & b[215])^(a[102] & b[216])^(a[101] & b[217])^(a[100] & b[218])^(a[99] & b[219])^(a[98] & b[220])^(a[97] & b[221])^(a[96] & b[222])^(a[95] & b[223])^(a[94] & b[224])^(a[93] & b[225])^(a[92] & b[226])^(a[91] & b[227])^(a[90] & b[228])^(a[89] & b[229])^(a[88] & b[230])^(a[87] & b[231])^(a[86] & b[232]);
assign y[319] = (a[232] & b[87])^(a[231] & b[88])^(a[230] & b[89])^(a[229] & b[90])^(a[228] & b[91])^(a[227] & b[92])^(a[226] & b[93])^(a[225] & b[94])^(a[224] & b[95])^(a[223] & b[96])^(a[222] & b[97])^(a[221] & b[98])^(a[220] & b[99])^(a[219] & b[100])^(a[218] & b[101])^(a[217] & b[102])^(a[216] & b[103])^(a[215] & b[104])^(a[214] & b[105])^(a[213] & b[106])^(a[212] & b[107])^(a[211] & b[108])^(a[210] & b[109])^(a[209] & b[110])^(a[208] & b[111])^(a[207] & b[112])^(a[206] & b[113])^(a[205] & b[114])^(a[204] & b[115])^(a[203] & b[116])^(a[202] & b[117])^(a[201] & b[118])^(a[200] & b[119])^(a[199] & b[120])^(a[198] & b[121])^(a[197] & b[122])^(a[196] & b[123])^(a[195] & b[124])^(a[194] & b[125])^(a[193] & b[126])^(a[192] & b[127])^(a[191] & b[128])^(a[190] & b[129])^(a[189] & b[130])^(a[188] & b[131])^(a[187] & b[132])^(a[186] & b[133])^(a[185] & b[134])^(a[184] & b[135])^(a[183] & b[136])^(a[182] & b[137])^(a[181] & b[138])^(a[180] & b[139])^(a[179] & b[140])^(a[178] & b[141])^(a[177] & b[142])^(a[176] & b[143])^(a[175] & b[144])^(a[174] & b[145])^(a[173] & b[146])^(a[172] & b[147])^(a[171] & b[148])^(a[170] & b[149])^(a[169] & b[150])^(a[168] & b[151])^(a[167] & b[152])^(a[166] & b[153])^(a[165] & b[154])^(a[164] & b[155])^(a[163] & b[156])^(a[162] & b[157])^(a[161] & b[158])^(a[160] & b[159])^(a[159] & b[160])^(a[158] & b[161])^(a[157] & b[162])^(a[156] & b[163])^(a[155] & b[164])^(a[154] & b[165])^(a[153] & b[166])^(a[152] & b[167])^(a[151] & b[168])^(a[150] & b[169])^(a[149] & b[170])^(a[148] & b[171])^(a[147] & b[172])^(a[146] & b[173])^(a[145] & b[174])^(a[144] & b[175])^(a[143] & b[176])^(a[142] & b[177])^(a[141] & b[178])^(a[140] & b[179])^(a[139] & b[180])^(a[138] & b[181])^(a[137] & b[182])^(a[136] & b[183])^(a[135] & b[184])^(a[134] & b[185])^(a[133] & b[186])^(a[132] & b[187])^(a[131] & b[188])^(a[130] & b[189])^(a[129] & b[190])^(a[128] & b[191])^(a[127] & b[192])^(a[126] & b[193])^(a[125] & b[194])^(a[124] & b[195])^(a[123] & b[196])^(a[122] & b[197])^(a[121] & b[198])^(a[120] & b[199])^(a[119] & b[200])^(a[118] & b[201])^(a[117] & b[202])^(a[116] & b[203])^(a[115] & b[204])^(a[114] & b[205])^(a[113] & b[206])^(a[112] & b[207])^(a[111] & b[208])^(a[110] & b[209])^(a[109] & b[210])^(a[108] & b[211])^(a[107] & b[212])^(a[106] & b[213])^(a[105] & b[214])^(a[104] & b[215])^(a[103] & b[216])^(a[102] & b[217])^(a[101] & b[218])^(a[100] & b[219])^(a[99] & b[220])^(a[98] & b[221])^(a[97] & b[222])^(a[96] & b[223])^(a[95] & b[224])^(a[94] & b[225])^(a[93] & b[226])^(a[92] & b[227])^(a[91] & b[228])^(a[90] & b[229])^(a[89] & b[230])^(a[88] & b[231])^(a[87] & b[232]);
assign y[320] = (a[232] & b[88])^(a[231] & b[89])^(a[230] & b[90])^(a[229] & b[91])^(a[228] & b[92])^(a[227] & b[93])^(a[226] & b[94])^(a[225] & b[95])^(a[224] & b[96])^(a[223] & b[97])^(a[222] & b[98])^(a[221] & b[99])^(a[220] & b[100])^(a[219] & b[101])^(a[218] & b[102])^(a[217] & b[103])^(a[216] & b[104])^(a[215] & b[105])^(a[214] & b[106])^(a[213] & b[107])^(a[212] & b[108])^(a[211] & b[109])^(a[210] & b[110])^(a[209] & b[111])^(a[208] & b[112])^(a[207] & b[113])^(a[206] & b[114])^(a[205] & b[115])^(a[204] & b[116])^(a[203] & b[117])^(a[202] & b[118])^(a[201] & b[119])^(a[200] & b[120])^(a[199] & b[121])^(a[198] & b[122])^(a[197] & b[123])^(a[196] & b[124])^(a[195] & b[125])^(a[194] & b[126])^(a[193] & b[127])^(a[192] & b[128])^(a[191] & b[129])^(a[190] & b[130])^(a[189] & b[131])^(a[188] & b[132])^(a[187] & b[133])^(a[186] & b[134])^(a[185] & b[135])^(a[184] & b[136])^(a[183] & b[137])^(a[182] & b[138])^(a[181] & b[139])^(a[180] & b[140])^(a[179] & b[141])^(a[178] & b[142])^(a[177] & b[143])^(a[176] & b[144])^(a[175] & b[145])^(a[174] & b[146])^(a[173] & b[147])^(a[172] & b[148])^(a[171] & b[149])^(a[170] & b[150])^(a[169] & b[151])^(a[168] & b[152])^(a[167] & b[153])^(a[166] & b[154])^(a[165] & b[155])^(a[164] & b[156])^(a[163] & b[157])^(a[162] & b[158])^(a[161] & b[159])^(a[160] & b[160])^(a[159] & b[161])^(a[158] & b[162])^(a[157] & b[163])^(a[156] & b[164])^(a[155] & b[165])^(a[154] & b[166])^(a[153] & b[167])^(a[152] & b[168])^(a[151] & b[169])^(a[150] & b[170])^(a[149] & b[171])^(a[148] & b[172])^(a[147] & b[173])^(a[146] & b[174])^(a[145] & b[175])^(a[144] & b[176])^(a[143] & b[177])^(a[142] & b[178])^(a[141] & b[179])^(a[140] & b[180])^(a[139] & b[181])^(a[138] & b[182])^(a[137] & b[183])^(a[136] & b[184])^(a[135] & b[185])^(a[134] & b[186])^(a[133] & b[187])^(a[132] & b[188])^(a[131] & b[189])^(a[130] & b[190])^(a[129] & b[191])^(a[128] & b[192])^(a[127] & b[193])^(a[126] & b[194])^(a[125] & b[195])^(a[124] & b[196])^(a[123] & b[197])^(a[122] & b[198])^(a[121] & b[199])^(a[120] & b[200])^(a[119] & b[201])^(a[118] & b[202])^(a[117] & b[203])^(a[116] & b[204])^(a[115] & b[205])^(a[114] & b[206])^(a[113] & b[207])^(a[112] & b[208])^(a[111] & b[209])^(a[110] & b[210])^(a[109] & b[211])^(a[108] & b[212])^(a[107] & b[213])^(a[106] & b[214])^(a[105] & b[215])^(a[104] & b[216])^(a[103] & b[217])^(a[102] & b[218])^(a[101] & b[219])^(a[100] & b[220])^(a[99] & b[221])^(a[98] & b[222])^(a[97] & b[223])^(a[96] & b[224])^(a[95] & b[225])^(a[94] & b[226])^(a[93] & b[227])^(a[92] & b[228])^(a[91] & b[229])^(a[90] & b[230])^(a[89] & b[231])^(a[88] & b[232]);
assign y[321] = (a[232] & b[89])^(a[231] & b[90])^(a[230] & b[91])^(a[229] & b[92])^(a[228] & b[93])^(a[227] & b[94])^(a[226] & b[95])^(a[225] & b[96])^(a[224] & b[97])^(a[223] & b[98])^(a[222] & b[99])^(a[221] & b[100])^(a[220] & b[101])^(a[219] & b[102])^(a[218] & b[103])^(a[217] & b[104])^(a[216] & b[105])^(a[215] & b[106])^(a[214] & b[107])^(a[213] & b[108])^(a[212] & b[109])^(a[211] & b[110])^(a[210] & b[111])^(a[209] & b[112])^(a[208] & b[113])^(a[207] & b[114])^(a[206] & b[115])^(a[205] & b[116])^(a[204] & b[117])^(a[203] & b[118])^(a[202] & b[119])^(a[201] & b[120])^(a[200] & b[121])^(a[199] & b[122])^(a[198] & b[123])^(a[197] & b[124])^(a[196] & b[125])^(a[195] & b[126])^(a[194] & b[127])^(a[193] & b[128])^(a[192] & b[129])^(a[191] & b[130])^(a[190] & b[131])^(a[189] & b[132])^(a[188] & b[133])^(a[187] & b[134])^(a[186] & b[135])^(a[185] & b[136])^(a[184] & b[137])^(a[183] & b[138])^(a[182] & b[139])^(a[181] & b[140])^(a[180] & b[141])^(a[179] & b[142])^(a[178] & b[143])^(a[177] & b[144])^(a[176] & b[145])^(a[175] & b[146])^(a[174] & b[147])^(a[173] & b[148])^(a[172] & b[149])^(a[171] & b[150])^(a[170] & b[151])^(a[169] & b[152])^(a[168] & b[153])^(a[167] & b[154])^(a[166] & b[155])^(a[165] & b[156])^(a[164] & b[157])^(a[163] & b[158])^(a[162] & b[159])^(a[161] & b[160])^(a[160] & b[161])^(a[159] & b[162])^(a[158] & b[163])^(a[157] & b[164])^(a[156] & b[165])^(a[155] & b[166])^(a[154] & b[167])^(a[153] & b[168])^(a[152] & b[169])^(a[151] & b[170])^(a[150] & b[171])^(a[149] & b[172])^(a[148] & b[173])^(a[147] & b[174])^(a[146] & b[175])^(a[145] & b[176])^(a[144] & b[177])^(a[143] & b[178])^(a[142] & b[179])^(a[141] & b[180])^(a[140] & b[181])^(a[139] & b[182])^(a[138] & b[183])^(a[137] & b[184])^(a[136] & b[185])^(a[135] & b[186])^(a[134] & b[187])^(a[133] & b[188])^(a[132] & b[189])^(a[131] & b[190])^(a[130] & b[191])^(a[129] & b[192])^(a[128] & b[193])^(a[127] & b[194])^(a[126] & b[195])^(a[125] & b[196])^(a[124] & b[197])^(a[123] & b[198])^(a[122] & b[199])^(a[121] & b[200])^(a[120] & b[201])^(a[119] & b[202])^(a[118] & b[203])^(a[117] & b[204])^(a[116] & b[205])^(a[115] & b[206])^(a[114] & b[207])^(a[113] & b[208])^(a[112] & b[209])^(a[111] & b[210])^(a[110] & b[211])^(a[109] & b[212])^(a[108] & b[213])^(a[107] & b[214])^(a[106] & b[215])^(a[105] & b[216])^(a[104] & b[217])^(a[103] & b[218])^(a[102] & b[219])^(a[101] & b[220])^(a[100] & b[221])^(a[99] & b[222])^(a[98] & b[223])^(a[97] & b[224])^(a[96] & b[225])^(a[95] & b[226])^(a[94] & b[227])^(a[93] & b[228])^(a[92] & b[229])^(a[91] & b[230])^(a[90] & b[231])^(a[89] & b[232]);
assign y[322] = (a[232] & b[90])^(a[231] & b[91])^(a[230] & b[92])^(a[229] & b[93])^(a[228] & b[94])^(a[227] & b[95])^(a[226] & b[96])^(a[225] & b[97])^(a[224] & b[98])^(a[223] & b[99])^(a[222] & b[100])^(a[221] & b[101])^(a[220] & b[102])^(a[219] & b[103])^(a[218] & b[104])^(a[217] & b[105])^(a[216] & b[106])^(a[215] & b[107])^(a[214] & b[108])^(a[213] & b[109])^(a[212] & b[110])^(a[211] & b[111])^(a[210] & b[112])^(a[209] & b[113])^(a[208] & b[114])^(a[207] & b[115])^(a[206] & b[116])^(a[205] & b[117])^(a[204] & b[118])^(a[203] & b[119])^(a[202] & b[120])^(a[201] & b[121])^(a[200] & b[122])^(a[199] & b[123])^(a[198] & b[124])^(a[197] & b[125])^(a[196] & b[126])^(a[195] & b[127])^(a[194] & b[128])^(a[193] & b[129])^(a[192] & b[130])^(a[191] & b[131])^(a[190] & b[132])^(a[189] & b[133])^(a[188] & b[134])^(a[187] & b[135])^(a[186] & b[136])^(a[185] & b[137])^(a[184] & b[138])^(a[183] & b[139])^(a[182] & b[140])^(a[181] & b[141])^(a[180] & b[142])^(a[179] & b[143])^(a[178] & b[144])^(a[177] & b[145])^(a[176] & b[146])^(a[175] & b[147])^(a[174] & b[148])^(a[173] & b[149])^(a[172] & b[150])^(a[171] & b[151])^(a[170] & b[152])^(a[169] & b[153])^(a[168] & b[154])^(a[167] & b[155])^(a[166] & b[156])^(a[165] & b[157])^(a[164] & b[158])^(a[163] & b[159])^(a[162] & b[160])^(a[161] & b[161])^(a[160] & b[162])^(a[159] & b[163])^(a[158] & b[164])^(a[157] & b[165])^(a[156] & b[166])^(a[155] & b[167])^(a[154] & b[168])^(a[153] & b[169])^(a[152] & b[170])^(a[151] & b[171])^(a[150] & b[172])^(a[149] & b[173])^(a[148] & b[174])^(a[147] & b[175])^(a[146] & b[176])^(a[145] & b[177])^(a[144] & b[178])^(a[143] & b[179])^(a[142] & b[180])^(a[141] & b[181])^(a[140] & b[182])^(a[139] & b[183])^(a[138] & b[184])^(a[137] & b[185])^(a[136] & b[186])^(a[135] & b[187])^(a[134] & b[188])^(a[133] & b[189])^(a[132] & b[190])^(a[131] & b[191])^(a[130] & b[192])^(a[129] & b[193])^(a[128] & b[194])^(a[127] & b[195])^(a[126] & b[196])^(a[125] & b[197])^(a[124] & b[198])^(a[123] & b[199])^(a[122] & b[200])^(a[121] & b[201])^(a[120] & b[202])^(a[119] & b[203])^(a[118] & b[204])^(a[117] & b[205])^(a[116] & b[206])^(a[115] & b[207])^(a[114] & b[208])^(a[113] & b[209])^(a[112] & b[210])^(a[111] & b[211])^(a[110] & b[212])^(a[109] & b[213])^(a[108] & b[214])^(a[107] & b[215])^(a[106] & b[216])^(a[105] & b[217])^(a[104] & b[218])^(a[103] & b[219])^(a[102] & b[220])^(a[101] & b[221])^(a[100] & b[222])^(a[99] & b[223])^(a[98] & b[224])^(a[97] & b[225])^(a[96] & b[226])^(a[95] & b[227])^(a[94] & b[228])^(a[93] & b[229])^(a[92] & b[230])^(a[91] & b[231])^(a[90] & b[232]);
assign y[323] = (a[232] & b[91])^(a[231] & b[92])^(a[230] & b[93])^(a[229] & b[94])^(a[228] & b[95])^(a[227] & b[96])^(a[226] & b[97])^(a[225] & b[98])^(a[224] & b[99])^(a[223] & b[100])^(a[222] & b[101])^(a[221] & b[102])^(a[220] & b[103])^(a[219] & b[104])^(a[218] & b[105])^(a[217] & b[106])^(a[216] & b[107])^(a[215] & b[108])^(a[214] & b[109])^(a[213] & b[110])^(a[212] & b[111])^(a[211] & b[112])^(a[210] & b[113])^(a[209] & b[114])^(a[208] & b[115])^(a[207] & b[116])^(a[206] & b[117])^(a[205] & b[118])^(a[204] & b[119])^(a[203] & b[120])^(a[202] & b[121])^(a[201] & b[122])^(a[200] & b[123])^(a[199] & b[124])^(a[198] & b[125])^(a[197] & b[126])^(a[196] & b[127])^(a[195] & b[128])^(a[194] & b[129])^(a[193] & b[130])^(a[192] & b[131])^(a[191] & b[132])^(a[190] & b[133])^(a[189] & b[134])^(a[188] & b[135])^(a[187] & b[136])^(a[186] & b[137])^(a[185] & b[138])^(a[184] & b[139])^(a[183] & b[140])^(a[182] & b[141])^(a[181] & b[142])^(a[180] & b[143])^(a[179] & b[144])^(a[178] & b[145])^(a[177] & b[146])^(a[176] & b[147])^(a[175] & b[148])^(a[174] & b[149])^(a[173] & b[150])^(a[172] & b[151])^(a[171] & b[152])^(a[170] & b[153])^(a[169] & b[154])^(a[168] & b[155])^(a[167] & b[156])^(a[166] & b[157])^(a[165] & b[158])^(a[164] & b[159])^(a[163] & b[160])^(a[162] & b[161])^(a[161] & b[162])^(a[160] & b[163])^(a[159] & b[164])^(a[158] & b[165])^(a[157] & b[166])^(a[156] & b[167])^(a[155] & b[168])^(a[154] & b[169])^(a[153] & b[170])^(a[152] & b[171])^(a[151] & b[172])^(a[150] & b[173])^(a[149] & b[174])^(a[148] & b[175])^(a[147] & b[176])^(a[146] & b[177])^(a[145] & b[178])^(a[144] & b[179])^(a[143] & b[180])^(a[142] & b[181])^(a[141] & b[182])^(a[140] & b[183])^(a[139] & b[184])^(a[138] & b[185])^(a[137] & b[186])^(a[136] & b[187])^(a[135] & b[188])^(a[134] & b[189])^(a[133] & b[190])^(a[132] & b[191])^(a[131] & b[192])^(a[130] & b[193])^(a[129] & b[194])^(a[128] & b[195])^(a[127] & b[196])^(a[126] & b[197])^(a[125] & b[198])^(a[124] & b[199])^(a[123] & b[200])^(a[122] & b[201])^(a[121] & b[202])^(a[120] & b[203])^(a[119] & b[204])^(a[118] & b[205])^(a[117] & b[206])^(a[116] & b[207])^(a[115] & b[208])^(a[114] & b[209])^(a[113] & b[210])^(a[112] & b[211])^(a[111] & b[212])^(a[110] & b[213])^(a[109] & b[214])^(a[108] & b[215])^(a[107] & b[216])^(a[106] & b[217])^(a[105] & b[218])^(a[104] & b[219])^(a[103] & b[220])^(a[102] & b[221])^(a[101] & b[222])^(a[100] & b[223])^(a[99] & b[224])^(a[98] & b[225])^(a[97] & b[226])^(a[96] & b[227])^(a[95] & b[228])^(a[94] & b[229])^(a[93] & b[230])^(a[92] & b[231])^(a[91] & b[232]);
assign y[324] = (a[232] & b[92])^(a[231] & b[93])^(a[230] & b[94])^(a[229] & b[95])^(a[228] & b[96])^(a[227] & b[97])^(a[226] & b[98])^(a[225] & b[99])^(a[224] & b[100])^(a[223] & b[101])^(a[222] & b[102])^(a[221] & b[103])^(a[220] & b[104])^(a[219] & b[105])^(a[218] & b[106])^(a[217] & b[107])^(a[216] & b[108])^(a[215] & b[109])^(a[214] & b[110])^(a[213] & b[111])^(a[212] & b[112])^(a[211] & b[113])^(a[210] & b[114])^(a[209] & b[115])^(a[208] & b[116])^(a[207] & b[117])^(a[206] & b[118])^(a[205] & b[119])^(a[204] & b[120])^(a[203] & b[121])^(a[202] & b[122])^(a[201] & b[123])^(a[200] & b[124])^(a[199] & b[125])^(a[198] & b[126])^(a[197] & b[127])^(a[196] & b[128])^(a[195] & b[129])^(a[194] & b[130])^(a[193] & b[131])^(a[192] & b[132])^(a[191] & b[133])^(a[190] & b[134])^(a[189] & b[135])^(a[188] & b[136])^(a[187] & b[137])^(a[186] & b[138])^(a[185] & b[139])^(a[184] & b[140])^(a[183] & b[141])^(a[182] & b[142])^(a[181] & b[143])^(a[180] & b[144])^(a[179] & b[145])^(a[178] & b[146])^(a[177] & b[147])^(a[176] & b[148])^(a[175] & b[149])^(a[174] & b[150])^(a[173] & b[151])^(a[172] & b[152])^(a[171] & b[153])^(a[170] & b[154])^(a[169] & b[155])^(a[168] & b[156])^(a[167] & b[157])^(a[166] & b[158])^(a[165] & b[159])^(a[164] & b[160])^(a[163] & b[161])^(a[162] & b[162])^(a[161] & b[163])^(a[160] & b[164])^(a[159] & b[165])^(a[158] & b[166])^(a[157] & b[167])^(a[156] & b[168])^(a[155] & b[169])^(a[154] & b[170])^(a[153] & b[171])^(a[152] & b[172])^(a[151] & b[173])^(a[150] & b[174])^(a[149] & b[175])^(a[148] & b[176])^(a[147] & b[177])^(a[146] & b[178])^(a[145] & b[179])^(a[144] & b[180])^(a[143] & b[181])^(a[142] & b[182])^(a[141] & b[183])^(a[140] & b[184])^(a[139] & b[185])^(a[138] & b[186])^(a[137] & b[187])^(a[136] & b[188])^(a[135] & b[189])^(a[134] & b[190])^(a[133] & b[191])^(a[132] & b[192])^(a[131] & b[193])^(a[130] & b[194])^(a[129] & b[195])^(a[128] & b[196])^(a[127] & b[197])^(a[126] & b[198])^(a[125] & b[199])^(a[124] & b[200])^(a[123] & b[201])^(a[122] & b[202])^(a[121] & b[203])^(a[120] & b[204])^(a[119] & b[205])^(a[118] & b[206])^(a[117] & b[207])^(a[116] & b[208])^(a[115] & b[209])^(a[114] & b[210])^(a[113] & b[211])^(a[112] & b[212])^(a[111] & b[213])^(a[110] & b[214])^(a[109] & b[215])^(a[108] & b[216])^(a[107] & b[217])^(a[106] & b[218])^(a[105] & b[219])^(a[104] & b[220])^(a[103] & b[221])^(a[102] & b[222])^(a[101] & b[223])^(a[100] & b[224])^(a[99] & b[225])^(a[98] & b[226])^(a[97] & b[227])^(a[96] & b[228])^(a[95] & b[229])^(a[94] & b[230])^(a[93] & b[231])^(a[92] & b[232]);
assign y[325] = (a[232] & b[93])^(a[231] & b[94])^(a[230] & b[95])^(a[229] & b[96])^(a[228] & b[97])^(a[227] & b[98])^(a[226] & b[99])^(a[225] & b[100])^(a[224] & b[101])^(a[223] & b[102])^(a[222] & b[103])^(a[221] & b[104])^(a[220] & b[105])^(a[219] & b[106])^(a[218] & b[107])^(a[217] & b[108])^(a[216] & b[109])^(a[215] & b[110])^(a[214] & b[111])^(a[213] & b[112])^(a[212] & b[113])^(a[211] & b[114])^(a[210] & b[115])^(a[209] & b[116])^(a[208] & b[117])^(a[207] & b[118])^(a[206] & b[119])^(a[205] & b[120])^(a[204] & b[121])^(a[203] & b[122])^(a[202] & b[123])^(a[201] & b[124])^(a[200] & b[125])^(a[199] & b[126])^(a[198] & b[127])^(a[197] & b[128])^(a[196] & b[129])^(a[195] & b[130])^(a[194] & b[131])^(a[193] & b[132])^(a[192] & b[133])^(a[191] & b[134])^(a[190] & b[135])^(a[189] & b[136])^(a[188] & b[137])^(a[187] & b[138])^(a[186] & b[139])^(a[185] & b[140])^(a[184] & b[141])^(a[183] & b[142])^(a[182] & b[143])^(a[181] & b[144])^(a[180] & b[145])^(a[179] & b[146])^(a[178] & b[147])^(a[177] & b[148])^(a[176] & b[149])^(a[175] & b[150])^(a[174] & b[151])^(a[173] & b[152])^(a[172] & b[153])^(a[171] & b[154])^(a[170] & b[155])^(a[169] & b[156])^(a[168] & b[157])^(a[167] & b[158])^(a[166] & b[159])^(a[165] & b[160])^(a[164] & b[161])^(a[163] & b[162])^(a[162] & b[163])^(a[161] & b[164])^(a[160] & b[165])^(a[159] & b[166])^(a[158] & b[167])^(a[157] & b[168])^(a[156] & b[169])^(a[155] & b[170])^(a[154] & b[171])^(a[153] & b[172])^(a[152] & b[173])^(a[151] & b[174])^(a[150] & b[175])^(a[149] & b[176])^(a[148] & b[177])^(a[147] & b[178])^(a[146] & b[179])^(a[145] & b[180])^(a[144] & b[181])^(a[143] & b[182])^(a[142] & b[183])^(a[141] & b[184])^(a[140] & b[185])^(a[139] & b[186])^(a[138] & b[187])^(a[137] & b[188])^(a[136] & b[189])^(a[135] & b[190])^(a[134] & b[191])^(a[133] & b[192])^(a[132] & b[193])^(a[131] & b[194])^(a[130] & b[195])^(a[129] & b[196])^(a[128] & b[197])^(a[127] & b[198])^(a[126] & b[199])^(a[125] & b[200])^(a[124] & b[201])^(a[123] & b[202])^(a[122] & b[203])^(a[121] & b[204])^(a[120] & b[205])^(a[119] & b[206])^(a[118] & b[207])^(a[117] & b[208])^(a[116] & b[209])^(a[115] & b[210])^(a[114] & b[211])^(a[113] & b[212])^(a[112] & b[213])^(a[111] & b[214])^(a[110] & b[215])^(a[109] & b[216])^(a[108] & b[217])^(a[107] & b[218])^(a[106] & b[219])^(a[105] & b[220])^(a[104] & b[221])^(a[103] & b[222])^(a[102] & b[223])^(a[101] & b[224])^(a[100] & b[225])^(a[99] & b[226])^(a[98] & b[227])^(a[97] & b[228])^(a[96] & b[229])^(a[95] & b[230])^(a[94] & b[231])^(a[93] & b[232]);
assign y[326] = (a[232] & b[94])^(a[231] & b[95])^(a[230] & b[96])^(a[229] & b[97])^(a[228] & b[98])^(a[227] & b[99])^(a[226] & b[100])^(a[225] & b[101])^(a[224] & b[102])^(a[223] & b[103])^(a[222] & b[104])^(a[221] & b[105])^(a[220] & b[106])^(a[219] & b[107])^(a[218] & b[108])^(a[217] & b[109])^(a[216] & b[110])^(a[215] & b[111])^(a[214] & b[112])^(a[213] & b[113])^(a[212] & b[114])^(a[211] & b[115])^(a[210] & b[116])^(a[209] & b[117])^(a[208] & b[118])^(a[207] & b[119])^(a[206] & b[120])^(a[205] & b[121])^(a[204] & b[122])^(a[203] & b[123])^(a[202] & b[124])^(a[201] & b[125])^(a[200] & b[126])^(a[199] & b[127])^(a[198] & b[128])^(a[197] & b[129])^(a[196] & b[130])^(a[195] & b[131])^(a[194] & b[132])^(a[193] & b[133])^(a[192] & b[134])^(a[191] & b[135])^(a[190] & b[136])^(a[189] & b[137])^(a[188] & b[138])^(a[187] & b[139])^(a[186] & b[140])^(a[185] & b[141])^(a[184] & b[142])^(a[183] & b[143])^(a[182] & b[144])^(a[181] & b[145])^(a[180] & b[146])^(a[179] & b[147])^(a[178] & b[148])^(a[177] & b[149])^(a[176] & b[150])^(a[175] & b[151])^(a[174] & b[152])^(a[173] & b[153])^(a[172] & b[154])^(a[171] & b[155])^(a[170] & b[156])^(a[169] & b[157])^(a[168] & b[158])^(a[167] & b[159])^(a[166] & b[160])^(a[165] & b[161])^(a[164] & b[162])^(a[163] & b[163])^(a[162] & b[164])^(a[161] & b[165])^(a[160] & b[166])^(a[159] & b[167])^(a[158] & b[168])^(a[157] & b[169])^(a[156] & b[170])^(a[155] & b[171])^(a[154] & b[172])^(a[153] & b[173])^(a[152] & b[174])^(a[151] & b[175])^(a[150] & b[176])^(a[149] & b[177])^(a[148] & b[178])^(a[147] & b[179])^(a[146] & b[180])^(a[145] & b[181])^(a[144] & b[182])^(a[143] & b[183])^(a[142] & b[184])^(a[141] & b[185])^(a[140] & b[186])^(a[139] & b[187])^(a[138] & b[188])^(a[137] & b[189])^(a[136] & b[190])^(a[135] & b[191])^(a[134] & b[192])^(a[133] & b[193])^(a[132] & b[194])^(a[131] & b[195])^(a[130] & b[196])^(a[129] & b[197])^(a[128] & b[198])^(a[127] & b[199])^(a[126] & b[200])^(a[125] & b[201])^(a[124] & b[202])^(a[123] & b[203])^(a[122] & b[204])^(a[121] & b[205])^(a[120] & b[206])^(a[119] & b[207])^(a[118] & b[208])^(a[117] & b[209])^(a[116] & b[210])^(a[115] & b[211])^(a[114] & b[212])^(a[113] & b[213])^(a[112] & b[214])^(a[111] & b[215])^(a[110] & b[216])^(a[109] & b[217])^(a[108] & b[218])^(a[107] & b[219])^(a[106] & b[220])^(a[105] & b[221])^(a[104] & b[222])^(a[103] & b[223])^(a[102] & b[224])^(a[101] & b[225])^(a[100] & b[226])^(a[99] & b[227])^(a[98] & b[228])^(a[97] & b[229])^(a[96] & b[230])^(a[95] & b[231])^(a[94] & b[232]);
assign y[327] = (a[232] & b[95])^(a[231] & b[96])^(a[230] & b[97])^(a[229] & b[98])^(a[228] & b[99])^(a[227] & b[100])^(a[226] & b[101])^(a[225] & b[102])^(a[224] & b[103])^(a[223] & b[104])^(a[222] & b[105])^(a[221] & b[106])^(a[220] & b[107])^(a[219] & b[108])^(a[218] & b[109])^(a[217] & b[110])^(a[216] & b[111])^(a[215] & b[112])^(a[214] & b[113])^(a[213] & b[114])^(a[212] & b[115])^(a[211] & b[116])^(a[210] & b[117])^(a[209] & b[118])^(a[208] & b[119])^(a[207] & b[120])^(a[206] & b[121])^(a[205] & b[122])^(a[204] & b[123])^(a[203] & b[124])^(a[202] & b[125])^(a[201] & b[126])^(a[200] & b[127])^(a[199] & b[128])^(a[198] & b[129])^(a[197] & b[130])^(a[196] & b[131])^(a[195] & b[132])^(a[194] & b[133])^(a[193] & b[134])^(a[192] & b[135])^(a[191] & b[136])^(a[190] & b[137])^(a[189] & b[138])^(a[188] & b[139])^(a[187] & b[140])^(a[186] & b[141])^(a[185] & b[142])^(a[184] & b[143])^(a[183] & b[144])^(a[182] & b[145])^(a[181] & b[146])^(a[180] & b[147])^(a[179] & b[148])^(a[178] & b[149])^(a[177] & b[150])^(a[176] & b[151])^(a[175] & b[152])^(a[174] & b[153])^(a[173] & b[154])^(a[172] & b[155])^(a[171] & b[156])^(a[170] & b[157])^(a[169] & b[158])^(a[168] & b[159])^(a[167] & b[160])^(a[166] & b[161])^(a[165] & b[162])^(a[164] & b[163])^(a[163] & b[164])^(a[162] & b[165])^(a[161] & b[166])^(a[160] & b[167])^(a[159] & b[168])^(a[158] & b[169])^(a[157] & b[170])^(a[156] & b[171])^(a[155] & b[172])^(a[154] & b[173])^(a[153] & b[174])^(a[152] & b[175])^(a[151] & b[176])^(a[150] & b[177])^(a[149] & b[178])^(a[148] & b[179])^(a[147] & b[180])^(a[146] & b[181])^(a[145] & b[182])^(a[144] & b[183])^(a[143] & b[184])^(a[142] & b[185])^(a[141] & b[186])^(a[140] & b[187])^(a[139] & b[188])^(a[138] & b[189])^(a[137] & b[190])^(a[136] & b[191])^(a[135] & b[192])^(a[134] & b[193])^(a[133] & b[194])^(a[132] & b[195])^(a[131] & b[196])^(a[130] & b[197])^(a[129] & b[198])^(a[128] & b[199])^(a[127] & b[200])^(a[126] & b[201])^(a[125] & b[202])^(a[124] & b[203])^(a[123] & b[204])^(a[122] & b[205])^(a[121] & b[206])^(a[120] & b[207])^(a[119] & b[208])^(a[118] & b[209])^(a[117] & b[210])^(a[116] & b[211])^(a[115] & b[212])^(a[114] & b[213])^(a[113] & b[214])^(a[112] & b[215])^(a[111] & b[216])^(a[110] & b[217])^(a[109] & b[218])^(a[108] & b[219])^(a[107] & b[220])^(a[106] & b[221])^(a[105] & b[222])^(a[104] & b[223])^(a[103] & b[224])^(a[102] & b[225])^(a[101] & b[226])^(a[100] & b[227])^(a[99] & b[228])^(a[98] & b[229])^(a[97] & b[230])^(a[96] & b[231])^(a[95] & b[232]);
assign y[328] = (a[232] & b[96])^(a[231] & b[97])^(a[230] & b[98])^(a[229] & b[99])^(a[228] & b[100])^(a[227] & b[101])^(a[226] & b[102])^(a[225] & b[103])^(a[224] & b[104])^(a[223] & b[105])^(a[222] & b[106])^(a[221] & b[107])^(a[220] & b[108])^(a[219] & b[109])^(a[218] & b[110])^(a[217] & b[111])^(a[216] & b[112])^(a[215] & b[113])^(a[214] & b[114])^(a[213] & b[115])^(a[212] & b[116])^(a[211] & b[117])^(a[210] & b[118])^(a[209] & b[119])^(a[208] & b[120])^(a[207] & b[121])^(a[206] & b[122])^(a[205] & b[123])^(a[204] & b[124])^(a[203] & b[125])^(a[202] & b[126])^(a[201] & b[127])^(a[200] & b[128])^(a[199] & b[129])^(a[198] & b[130])^(a[197] & b[131])^(a[196] & b[132])^(a[195] & b[133])^(a[194] & b[134])^(a[193] & b[135])^(a[192] & b[136])^(a[191] & b[137])^(a[190] & b[138])^(a[189] & b[139])^(a[188] & b[140])^(a[187] & b[141])^(a[186] & b[142])^(a[185] & b[143])^(a[184] & b[144])^(a[183] & b[145])^(a[182] & b[146])^(a[181] & b[147])^(a[180] & b[148])^(a[179] & b[149])^(a[178] & b[150])^(a[177] & b[151])^(a[176] & b[152])^(a[175] & b[153])^(a[174] & b[154])^(a[173] & b[155])^(a[172] & b[156])^(a[171] & b[157])^(a[170] & b[158])^(a[169] & b[159])^(a[168] & b[160])^(a[167] & b[161])^(a[166] & b[162])^(a[165] & b[163])^(a[164] & b[164])^(a[163] & b[165])^(a[162] & b[166])^(a[161] & b[167])^(a[160] & b[168])^(a[159] & b[169])^(a[158] & b[170])^(a[157] & b[171])^(a[156] & b[172])^(a[155] & b[173])^(a[154] & b[174])^(a[153] & b[175])^(a[152] & b[176])^(a[151] & b[177])^(a[150] & b[178])^(a[149] & b[179])^(a[148] & b[180])^(a[147] & b[181])^(a[146] & b[182])^(a[145] & b[183])^(a[144] & b[184])^(a[143] & b[185])^(a[142] & b[186])^(a[141] & b[187])^(a[140] & b[188])^(a[139] & b[189])^(a[138] & b[190])^(a[137] & b[191])^(a[136] & b[192])^(a[135] & b[193])^(a[134] & b[194])^(a[133] & b[195])^(a[132] & b[196])^(a[131] & b[197])^(a[130] & b[198])^(a[129] & b[199])^(a[128] & b[200])^(a[127] & b[201])^(a[126] & b[202])^(a[125] & b[203])^(a[124] & b[204])^(a[123] & b[205])^(a[122] & b[206])^(a[121] & b[207])^(a[120] & b[208])^(a[119] & b[209])^(a[118] & b[210])^(a[117] & b[211])^(a[116] & b[212])^(a[115] & b[213])^(a[114] & b[214])^(a[113] & b[215])^(a[112] & b[216])^(a[111] & b[217])^(a[110] & b[218])^(a[109] & b[219])^(a[108] & b[220])^(a[107] & b[221])^(a[106] & b[222])^(a[105] & b[223])^(a[104] & b[224])^(a[103] & b[225])^(a[102] & b[226])^(a[101] & b[227])^(a[100] & b[228])^(a[99] & b[229])^(a[98] & b[230])^(a[97] & b[231])^(a[96] & b[232]);
assign y[329] = (a[232] & b[97])^(a[231] & b[98])^(a[230] & b[99])^(a[229] & b[100])^(a[228] & b[101])^(a[227] & b[102])^(a[226] & b[103])^(a[225] & b[104])^(a[224] & b[105])^(a[223] & b[106])^(a[222] & b[107])^(a[221] & b[108])^(a[220] & b[109])^(a[219] & b[110])^(a[218] & b[111])^(a[217] & b[112])^(a[216] & b[113])^(a[215] & b[114])^(a[214] & b[115])^(a[213] & b[116])^(a[212] & b[117])^(a[211] & b[118])^(a[210] & b[119])^(a[209] & b[120])^(a[208] & b[121])^(a[207] & b[122])^(a[206] & b[123])^(a[205] & b[124])^(a[204] & b[125])^(a[203] & b[126])^(a[202] & b[127])^(a[201] & b[128])^(a[200] & b[129])^(a[199] & b[130])^(a[198] & b[131])^(a[197] & b[132])^(a[196] & b[133])^(a[195] & b[134])^(a[194] & b[135])^(a[193] & b[136])^(a[192] & b[137])^(a[191] & b[138])^(a[190] & b[139])^(a[189] & b[140])^(a[188] & b[141])^(a[187] & b[142])^(a[186] & b[143])^(a[185] & b[144])^(a[184] & b[145])^(a[183] & b[146])^(a[182] & b[147])^(a[181] & b[148])^(a[180] & b[149])^(a[179] & b[150])^(a[178] & b[151])^(a[177] & b[152])^(a[176] & b[153])^(a[175] & b[154])^(a[174] & b[155])^(a[173] & b[156])^(a[172] & b[157])^(a[171] & b[158])^(a[170] & b[159])^(a[169] & b[160])^(a[168] & b[161])^(a[167] & b[162])^(a[166] & b[163])^(a[165] & b[164])^(a[164] & b[165])^(a[163] & b[166])^(a[162] & b[167])^(a[161] & b[168])^(a[160] & b[169])^(a[159] & b[170])^(a[158] & b[171])^(a[157] & b[172])^(a[156] & b[173])^(a[155] & b[174])^(a[154] & b[175])^(a[153] & b[176])^(a[152] & b[177])^(a[151] & b[178])^(a[150] & b[179])^(a[149] & b[180])^(a[148] & b[181])^(a[147] & b[182])^(a[146] & b[183])^(a[145] & b[184])^(a[144] & b[185])^(a[143] & b[186])^(a[142] & b[187])^(a[141] & b[188])^(a[140] & b[189])^(a[139] & b[190])^(a[138] & b[191])^(a[137] & b[192])^(a[136] & b[193])^(a[135] & b[194])^(a[134] & b[195])^(a[133] & b[196])^(a[132] & b[197])^(a[131] & b[198])^(a[130] & b[199])^(a[129] & b[200])^(a[128] & b[201])^(a[127] & b[202])^(a[126] & b[203])^(a[125] & b[204])^(a[124] & b[205])^(a[123] & b[206])^(a[122] & b[207])^(a[121] & b[208])^(a[120] & b[209])^(a[119] & b[210])^(a[118] & b[211])^(a[117] & b[212])^(a[116] & b[213])^(a[115] & b[214])^(a[114] & b[215])^(a[113] & b[216])^(a[112] & b[217])^(a[111] & b[218])^(a[110] & b[219])^(a[109] & b[220])^(a[108] & b[221])^(a[107] & b[222])^(a[106] & b[223])^(a[105] & b[224])^(a[104] & b[225])^(a[103] & b[226])^(a[102] & b[227])^(a[101] & b[228])^(a[100] & b[229])^(a[99] & b[230])^(a[98] & b[231])^(a[97] & b[232]);
assign y[330] = (a[232] & b[98])^(a[231] & b[99])^(a[230] & b[100])^(a[229] & b[101])^(a[228] & b[102])^(a[227] & b[103])^(a[226] & b[104])^(a[225] & b[105])^(a[224] & b[106])^(a[223] & b[107])^(a[222] & b[108])^(a[221] & b[109])^(a[220] & b[110])^(a[219] & b[111])^(a[218] & b[112])^(a[217] & b[113])^(a[216] & b[114])^(a[215] & b[115])^(a[214] & b[116])^(a[213] & b[117])^(a[212] & b[118])^(a[211] & b[119])^(a[210] & b[120])^(a[209] & b[121])^(a[208] & b[122])^(a[207] & b[123])^(a[206] & b[124])^(a[205] & b[125])^(a[204] & b[126])^(a[203] & b[127])^(a[202] & b[128])^(a[201] & b[129])^(a[200] & b[130])^(a[199] & b[131])^(a[198] & b[132])^(a[197] & b[133])^(a[196] & b[134])^(a[195] & b[135])^(a[194] & b[136])^(a[193] & b[137])^(a[192] & b[138])^(a[191] & b[139])^(a[190] & b[140])^(a[189] & b[141])^(a[188] & b[142])^(a[187] & b[143])^(a[186] & b[144])^(a[185] & b[145])^(a[184] & b[146])^(a[183] & b[147])^(a[182] & b[148])^(a[181] & b[149])^(a[180] & b[150])^(a[179] & b[151])^(a[178] & b[152])^(a[177] & b[153])^(a[176] & b[154])^(a[175] & b[155])^(a[174] & b[156])^(a[173] & b[157])^(a[172] & b[158])^(a[171] & b[159])^(a[170] & b[160])^(a[169] & b[161])^(a[168] & b[162])^(a[167] & b[163])^(a[166] & b[164])^(a[165] & b[165])^(a[164] & b[166])^(a[163] & b[167])^(a[162] & b[168])^(a[161] & b[169])^(a[160] & b[170])^(a[159] & b[171])^(a[158] & b[172])^(a[157] & b[173])^(a[156] & b[174])^(a[155] & b[175])^(a[154] & b[176])^(a[153] & b[177])^(a[152] & b[178])^(a[151] & b[179])^(a[150] & b[180])^(a[149] & b[181])^(a[148] & b[182])^(a[147] & b[183])^(a[146] & b[184])^(a[145] & b[185])^(a[144] & b[186])^(a[143] & b[187])^(a[142] & b[188])^(a[141] & b[189])^(a[140] & b[190])^(a[139] & b[191])^(a[138] & b[192])^(a[137] & b[193])^(a[136] & b[194])^(a[135] & b[195])^(a[134] & b[196])^(a[133] & b[197])^(a[132] & b[198])^(a[131] & b[199])^(a[130] & b[200])^(a[129] & b[201])^(a[128] & b[202])^(a[127] & b[203])^(a[126] & b[204])^(a[125] & b[205])^(a[124] & b[206])^(a[123] & b[207])^(a[122] & b[208])^(a[121] & b[209])^(a[120] & b[210])^(a[119] & b[211])^(a[118] & b[212])^(a[117] & b[213])^(a[116] & b[214])^(a[115] & b[215])^(a[114] & b[216])^(a[113] & b[217])^(a[112] & b[218])^(a[111] & b[219])^(a[110] & b[220])^(a[109] & b[221])^(a[108] & b[222])^(a[107] & b[223])^(a[106] & b[224])^(a[105] & b[225])^(a[104] & b[226])^(a[103] & b[227])^(a[102] & b[228])^(a[101] & b[229])^(a[100] & b[230])^(a[99] & b[231])^(a[98] & b[232]);
assign y[331] = (a[232] & b[99])^(a[231] & b[100])^(a[230] & b[101])^(a[229] & b[102])^(a[228] & b[103])^(a[227] & b[104])^(a[226] & b[105])^(a[225] & b[106])^(a[224] & b[107])^(a[223] & b[108])^(a[222] & b[109])^(a[221] & b[110])^(a[220] & b[111])^(a[219] & b[112])^(a[218] & b[113])^(a[217] & b[114])^(a[216] & b[115])^(a[215] & b[116])^(a[214] & b[117])^(a[213] & b[118])^(a[212] & b[119])^(a[211] & b[120])^(a[210] & b[121])^(a[209] & b[122])^(a[208] & b[123])^(a[207] & b[124])^(a[206] & b[125])^(a[205] & b[126])^(a[204] & b[127])^(a[203] & b[128])^(a[202] & b[129])^(a[201] & b[130])^(a[200] & b[131])^(a[199] & b[132])^(a[198] & b[133])^(a[197] & b[134])^(a[196] & b[135])^(a[195] & b[136])^(a[194] & b[137])^(a[193] & b[138])^(a[192] & b[139])^(a[191] & b[140])^(a[190] & b[141])^(a[189] & b[142])^(a[188] & b[143])^(a[187] & b[144])^(a[186] & b[145])^(a[185] & b[146])^(a[184] & b[147])^(a[183] & b[148])^(a[182] & b[149])^(a[181] & b[150])^(a[180] & b[151])^(a[179] & b[152])^(a[178] & b[153])^(a[177] & b[154])^(a[176] & b[155])^(a[175] & b[156])^(a[174] & b[157])^(a[173] & b[158])^(a[172] & b[159])^(a[171] & b[160])^(a[170] & b[161])^(a[169] & b[162])^(a[168] & b[163])^(a[167] & b[164])^(a[166] & b[165])^(a[165] & b[166])^(a[164] & b[167])^(a[163] & b[168])^(a[162] & b[169])^(a[161] & b[170])^(a[160] & b[171])^(a[159] & b[172])^(a[158] & b[173])^(a[157] & b[174])^(a[156] & b[175])^(a[155] & b[176])^(a[154] & b[177])^(a[153] & b[178])^(a[152] & b[179])^(a[151] & b[180])^(a[150] & b[181])^(a[149] & b[182])^(a[148] & b[183])^(a[147] & b[184])^(a[146] & b[185])^(a[145] & b[186])^(a[144] & b[187])^(a[143] & b[188])^(a[142] & b[189])^(a[141] & b[190])^(a[140] & b[191])^(a[139] & b[192])^(a[138] & b[193])^(a[137] & b[194])^(a[136] & b[195])^(a[135] & b[196])^(a[134] & b[197])^(a[133] & b[198])^(a[132] & b[199])^(a[131] & b[200])^(a[130] & b[201])^(a[129] & b[202])^(a[128] & b[203])^(a[127] & b[204])^(a[126] & b[205])^(a[125] & b[206])^(a[124] & b[207])^(a[123] & b[208])^(a[122] & b[209])^(a[121] & b[210])^(a[120] & b[211])^(a[119] & b[212])^(a[118] & b[213])^(a[117] & b[214])^(a[116] & b[215])^(a[115] & b[216])^(a[114] & b[217])^(a[113] & b[218])^(a[112] & b[219])^(a[111] & b[220])^(a[110] & b[221])^(a[109] & b[222])^(a[108] & b[223])^(a[107] & b[224])^(a[106] & b[225])^(a[105] & b[226])^(a[104] & b[227])^(a[103] & b[228])^(a[102] & b[229])^(a[101] & b[230])^(a[100] & b[231])^(a[99] & b[232]);
assign y[332] = (a[232] & b[100])^(a[231] & b[101])^(a[230] & b[102])^(a[229] & b[103])^(a[228] & b[104])^(a[227] & b[105])^(a[226] & b[106])^(a[225] & b[107])^(a[224] & b[108])^(a[223] & b[109])^(a[222] & b[110])^(a[221] & b[111])^(a[220] & b[112])^(a[219] & b[113])^(a[218] & b[114])^(a[217] & b[115])^(a[216] & b[116])^(a[215] & b[117])^(a[214] & b[118])^(a[213] & b[119])^(a[212] & b[120])^(a[211] & b[121])^(a[210] & b[122])^(a[209] & b[123])^(a[208] & b[124])^(a[207] & b[125])^(a[206] & b[126])^(a[205] & b[127])^(a[204] & b[128])^(a[203] & b[129])^(a[202] & b[130])^(a[201] & b[131])^(a[200] & b[132])^(a[199] & b[133])^(a[198] & b[134])^(a[197] & b[135])^(a[196] & b[136])^(a[195] & b[137])^(a[194] & b[138])^(a[193] & b[139])^(a[192] & b[140])^(a[191] & b[141])^(a[190] & b[142])^(a[189] & b[143])^(a[188] & b[144])^(a[187] & b[145])^(a[186] & b[146])^(a[185] & b[147])^(a[184] & b[148])^(a[183] & b[149])^(a[182] & b[150])^(a[181] & b[151])^(a[180] & b[152])^(a[179] & b[153])^(a[178] & b[154])^(a[177] & b[155])^(a[176] & b[156])^(a[175] & b[157])^(a[174] & b[158])^(a[173] & b[159])^(a[172] & b[160])^(a[171] & b[161])^(a[170] & b[162])^(a[169] & b[163])^(a[168] & b[164])^(a[167] & b[165])^(a[166] & b[166])^(a[165] & b[167])^(a[164] & b[168])^(a[163] & b[169])^(a[162] & b[170])^(a[161] & b[171])^(a[160] & b[172])^(a[159] & b[173])^(a[158] & b[174])^(a[157] & b[175])^(a[156] & b[176])^(a[155] & b[177])^(a[154] & b[178])^(a[153] & b[179])^(a[152] & b[180])^(a[151] & b[181])^(a[150] & b[182])^(a[149] & b[183])^(a[148] & b[184])^(a[147] & b[185])^(a[146] & b[186])^(a[145] & b[187])^(a[144] & b[188])^(a[143] & b[189])^(a[142] & b[190])^(a[141] & b[191])^(a[140] & b[192])^(a[139] & b[193])^(a[138] & b[194])^(a[137] & b[195])^(a[136] & b[196])^(a[135] & b[197])^(a[134] & b[198])^(a[133] & b[199])^(a[132] & b[200])^(a[131] & b[201])^(a[130] & b[202])^(a[129] & b[203])^(a[128] & b[204])^(a[127] & b[205])^(a[126] & b[206])^(a[125] & b[207])^(a[124] & b[208])^(a[123] & b[209])^(a[122] & b[210])^(a[121] & b[211])^(a[120] & b[212])^(a[119] & b[213])^(a[118] & b[214])^(a[117] & b[215])^(a[116] & b[216])^(a[115] & b[217])^(a[114] & b[218])^(a[113] & b[219])^(a[112] & b[220])^(a[111] & b[221])^(a[110] & b[222])^(a[109] & b[223])^(a[108] & b[224])^(a[107] & b[225])^(a[106] & b[226])^(a[105] & b[227])^(a[104] & b[228])^(a[103] & b[229])^(a[102] & b[230])^(a[101] & b[231])^(a[100] & b[232]);
assign y[333] = (a[232] & b[101])^(a[231] & b[102])^(a[230] & b[103])^(a[229] & b[104])^(a[228] & b[105])^(a[227] & b[106])^(a[226] & b[107])^(a[225] & b[108])^(a[224] & b[109])^(a[223] & b[110])^(a[222] & b[111])^(a[221] & b[112])^(a[220] & b[113])^(a[219] & b[114])^(a[218] & b[115])^(a[217] & b[116])^(a[216] & b[117])^(a[215] & b[118])^(a[214] & b[119])^(a[213] & b[120])^(a[212] & b[121])^(a[211] & b[122])^(a[210] & b[123])^(a[209] & b[124])^(a[208] & b[125])^(a[207] & b[126])^(a[206] & b[127])^(a[205] & b[128])^(a[204] & b[129])^(a[203] & b[130])^(a[202] & b[131])^(a[201] & b[132])^(a[200] & b[133])^(a[199] & b[134])^(a[198] & b[135])^(a[197] & b[136])^(a[196] & b[137])^(a[195] & b[138])^(a[194] & b[139])^(a[193] & b[140])^(a[192] & b[141])^(a[191] & b[142])^(a[190] & b[143])^(a[189] & b[144])^(a[188] & b[145])^(a[187] & b[146])^(a[186] & b[147])^(a[185] & b[148])^(a[184] & b[149])^(a[183] & b[150])^(a[182] & b[151])^(a[181] & b[152])^(a[180] & b[153])^(a[179] & b[154])^(a[178] & b[155])^(a[177] & b[156])^(a[176] & b[157])^(a[175] & b[158])^(a[174] & b[159])^(a[173] & b[160])^(a[172] & b[161])^(a[171] & b[162])^(a[170] & b[163])^(a[169] & b[164])^(a[168] & b[165])^(a[167] & b[166])^(a[166] & b[167])^(a[165] & b[168])^(a[164] & b[169])^(a[163] & b[170])^(a[162] & b[171])^(a[161] & b[172])^(a[160] & b[173])^(a[159] & b[174])^(a[158] & b[175])^(a[157] & b[176])^(a[156] & b[177])^(a[155] & b[178])^(a[154] & b[179])^(a[153] & b[180])^(a[152] & b[181])^(a[151] & b[182])^(a[150] & b[183])^(a[149] & b[184])^(a[148] & b[185])^(a[147] & b[186])^(a[146] & b[187])^(a[145] & b[188])^(a[144] & b[189])^(a[143] & b[190])^(a[142] & b[191])^(a[141] & b[192])^(a[140] & b[193])^(a[139] & b[194])^(a[138] & b[195])^(a[137] & b[196])^(a[136] & b[197])^(a[135] & b[198])^(a[134] & b[199])^(a[133] & b[200])^(a[132] & b[201])^(a[131] & b[202])^(a[130] & b[203])^(a[129] & b[204])^(a[128] & b[205])^(a[127] & b[206])^(a[126] & b[207])^(a[125] & b[208])^(a[124] & b[209])^(a[123] & b[210])^(a[122] & b[211])^(a[121] & b[212])^(a[120] & b[213])^(a[119] & b[214])^(a[118] & b[215])^(a[117] & b[216])^(a[116] & b[217])^(a[115] & b[218])^(a[114] & b[219])^(a[113] & b[220])^(a[112] & b[221])^(a[111] & b[222])^(a[110] & b[223])^(a[109] & b[224])^(a[108] & b[225])^(a[107] & b[226])^(a[106] & b[227])^(a[105] & b[228])^(a[104] & b[229])^(a[103] & b[230])^(a[102] & b[231])^(a[101] & b[232]);
assign y[334] = (a[232] & b[102])^(a[231] & b[103])^(a[230] & b[104])^(a[229] & b[105])^(a[228] & b[106])^(a[227] & b[107])^(a[226] & b[108])^(a[225] & b[109])^(a[224] & b[110])^(a[223] & b[111])^(a[222] & b[112])^(a[221] & b[113])^(a[220] & b[114])^(a[219] & b[115])^(a[218] & b[116])^(a[217] & b[117])^(a[216] & b[118])^(a[215] & b[119])^(a[214] & b[120])^(a[213] & b[121])^(a[212] & b[122])^(a[211] & b[123])^(a[210] & b[124])^(a[209] & b[125])^(a[208] & b[126])^(a[207] & b[127])^(a[206] & b[128])^(a[205] & b[129])^(a[204] & b[130])^(a[203] & b[131])^(a[202] & b[132])^(a[201] & b[133])^(a[200] & b[134])^(a[199] & b[135])^(a[198] & b[136])^(a[197] & b[137])^(a[196] & b[138])^(a[195] & b[139])^(a[194] & b[140])^(a[193] & b[141])^(a[192] & b[142])^(a[191] & b[143])^(a[190] & b[144])^(a[189] & b[145])^(a[188] & b[146])^(a[187] & b[147])^(a[186] & b[148])^(a[185] & b[149])^(a[184] & b[150])^(a[183] & b[151])^(a[182] & b[152])^(a[181] & b[153])^(a[180] & b[154])^(a[179] & b[155])^(a[178] & b[156])^(a[177] & b[157])^(a[176] & b[158])^(a[175] & b[159])^(a[174] & b[160])^(a[173] & b[161])^(a[172] & b[162])^(a[171] & b[163])^(a[170] & b[164])^(a[169] & b[165])^(a[168] & b[166])^(a[167] & b[167])^(a[166] & b[168])^(a[165] & b[169])^(a[164] & b[170])^(a[163] & b[171])^(a[162] & b[172])^(a[161] & b[173])^(a[160] & b[174])^(a[159] & b[175])^(a[158] & b[176])^(a[157] & b[177])^(a[156] & b[178])^(a[155] & b[179])^(a[154] & b[180])^(a[153] & b[181])^(a[152] & b[182])^(a[151] & b[183])^(a[150] & b[184])^(a[149] & b[185])^(a[148] & b[186])^(a[147] & b[187])^(a[146] & b[188])^(a[145] & b[189])^(a[144] & b[190])^(a[143] & b[191])^(a[142] & b[192])^(a[141] & b[193])^(a[140] & b[194])^(a[139] & b[195])^(a[138] & b[196])^(a[137] & b[197])^(a[136] & b[198])^(a[135] & b[199])^(a[134] & b[200])^(a[133] & b[201])^(a[132] & b[202])^(a[131] & b[203])^(a[130] & b[204])^(a[129] & b[205])^(a[128] & b[206])^(a[127] & b[207])^(a[126] & b[208])^(a[125] & b[209])^(a[124] & b[210])^(a[123] & b[211])^(a[122] & b[212])^(a[121] & b[213])^(a[120] & b[214])^(a[119] & b[215])^(a[118] & b[216])^(a[117] & b[217])^(a[116] & b[218])^(a[115] & b[219])^(a[114] & b[220])^(a[113] & b[221])^(a[112] & b[222])^(a[111] & b[223])^(a[110] & b[224])^(a[109] & b[225])^(a[108] & b[226])^(a[107] & b[227])^(a[106] & b[228])^(a[105] & b[229])^(a[104] & b[230])^(a[103] & b[231])^(a[102] & b[232]);
assign y[335] = (a[232] & b[103])^(a[231] & b[104])^(a[230] & b[105])^(a[229] & b[106])^(a[228] & b[107])^(a[227] & b[108])^(a[226] & b[109])^(a[225] & b[110])^(a[224] & b[111])^(a[223] & b[112])^(a[222] & b[113])^(a[221] & b[114])^(a[220] & b[115])^(a[219] & b[116])^(a[218] & b[117])^(a[217] & b[118])^(a[216] & b[119])^(a[215] & b[120])^(a[214] & b[121])^(a[213] & b[122])^(a[212] & b[123])^(a[211] & b[124])^(a[210] & b[125])^(a[209] & b[126])^(a[208] & b[127])^(a[207] & b[128])^(a[206] & b[129])^(a[205] & b[130])^(a[204] & b[131])^(a[203] & b[132])^(a[202] & b[133])^(a[201] & b[134])^(a[200] & b[135])^(a[199] & b[136])^(a[198] & b[137])^(a[197] & b[138])^(a[196] & b[139])^(a[195] & b[140])^(a[194] & b[141])^(a[193] & b[142])^(a[192] & b[143])^(a[191] & b[144])^(a[190] & b[145])^(a[189] & b[146])^(a[188] & b[147])^(a[187] & b[148])^(a[186] & b[149])^(a[185] & b[150])^(a[184] & b[151])^(a[183] & b[152])^(a[182] & b[153])^(a[181] & b[154])^(a[180] & b[155])^(a[179] & b[156])^(a[178] & b[157])^(a[177] & b[158])^(a[176] & b[159])^(a[175] & b[160])^(a[174] & b[161])^(a[173] & b[162])^(a[172] & b[163])^(a[171] & b[164])^(a[170] & b[165])^(a[169] & b[166])^(a[168] & b[167])^(a[167] & b[168])^(a[166] & b[169])^(a[165] & b[170])^(a[164] & b[171])^(a[163] & b[172])^(a[162] & b[173])^(a[161] & b[174])^(a[160] & b[175])^(a[159] & b[176])^(a[158] & b[177])^(a[157] & b[178])^(a[156] & b[179])^(a[155] & b[180])^(a[154] & b[181])^(a[153] & b[182])^(a[152] & b[183])^(a[151] & b[184])^(a[150] & b[185])^(a[149] & b[186])^(a[148] & b[187])^(a[147] & b[188])^(a[146] & b[189])^(a[145] & b[190])^(a[144] & b[191])^(a[143] & b[192])^(a[142] & b[193])^(a[141] & b[194])^(a[140] & b[195])^(a[139] & b[196])^(a[138] & b[197])^(a[137] & b[198])^(a[136] & b[199])^(a[135] & b[200])^(a[134] & b[201])^(a[133] & b[202])^(a[132] & b[203])^(a[131] & b[204])^(a[130] & b[205])^(a[129] & b[206])^(a[128] & b[207])^(a[127] & b[208])^(a[126] & b[209])^(a[125] & b[210])^(a[124] & b[211])^(a[123] & b[212])^(a[122] & b[213])^(a[121] & b[214])^(a[120] & b[215])^(a[119] & b[216])^(a[118] & b[217])^(a[117] & b[218])^(a[116] & b[219])^(a[115] & b[220])^(a[114] & b[221])^(a[113] & b[222])^(a[112] & b[223])^(a[111] & b[224])^(a[110] & b[225])^(a[109] & b[226])^(a[108] & b[227])^(a[107] & b[228])^(a[106] & b[229])^(a[105] & b[230])^(a[104] & b[231])^(a[103] & b[232]);
assign y[336] = (a[232] & b[104])^(a[231] & b[105])^(a[230] & b[106])^(a[229] & b[107])^(a[228] & b[108])^(a[227] & b[109])^(a[226] & b[110])^(a[225] & b[111])^(a[224] & b[112])^(a[223] & b[113])^(a[222] & b[114])^(a[221] & b[115])^(a[220] & b[116])^(a[219] & b[117])^(a[218] & b[118])^(a[217] & b[119])^(a[216] & b[120])^(a[215] & b[121])^(a[214] & b[122])^(a[213] & b[123])^(a[212] & b[124])^(a[211] & b[125])^(a[210] & b[126])^(a[209] & b[127])^(a[208] & b[128])^(a[207] & b[129])^(a[206] & b[130])^(a[205] & b[131])^(a[204] & b[132])^(a[203] & b[133])^(a[202] & b[134])^(a[201] & b[135])^(a[200] & b[136])^(a[199] & b[137])^(a[198] & b[138])^(a[197] & b[139])^(a[196] & b[140])^(a[195] & b[141])^(a[194] & b[142])^(a[193] & b[143])^(a[192] & b[144])^(a[191] & b[145])^(a[190] & b[146])^(a[189] & b[147])^(a[188] & b[148])^(a[187] & b[149])^(a[186] & b[150])^(a[185] & b[151])^(a[184] & b[152])^(a[183] & b[153])^(a[182] & b[154])^(a[181] & b[155])^(a[180] & b[156])^(a[179] & b[157])^(a[178] & b[158])^(a[177] & b[159])^(a[176] & b[160])^(a[175] & b[161])^(a[174] & b[162])^(a[173] & b[163])^(a[172] & b[164])^(a[171] & b[165])^(a[170] & b[166])^(a[169] & b[167])^(a[168] & b[168])^(a[167] & b[169])^(a[166] & b[170])^(a[165] & b[171])^(a[164] & b[172])^(a[163] & b[173])^(a[162] & b[174])^(a[161] & b[175])^(a[160] & b[176])^(a[159] & b[177])^(a[158] & b[178])^(a[157] & b[179])^(a[156] & b[180])^(a[155] & b[181])^(a[154] & b[182])^(a[153] & b[183])^(a[152] & b[184])^(a[151] & b[185])^(a[150] & b[186])^(a[149] & b[187])^(a[148] & b[188])^(a[147] & b[189])^(a[146] & b[190])^(a[145] & b[191])^(a[144] & b[192])^(a[143] & b[193])^(a[142] & b[194])^(a[141] & b[195])^(a[140] & b[196])^(a[139] & b[197])^(a[138] & b[198])^(a[137] & b[199])^(a[136] & b[200])^(a[135] & b[201])^(a[134] & b[202])^(a[133] & b[203])^(a[132] & b[204])^(a[131] & b[205])^(a[130] & b[206])^(a[129] & b[207])^(a[128] & b[208])^(a[127] & b[209])^(a[126] & b[210])^(a[125] & b[211])^(a[124] & b[212])^(a[123] & b[213])^(a[122] & b[214])^(a[121] & b[215])^(a[120] & b[216])^(a[119] & b[217])^(a[118] & b[218])^(a[117] & b[219])^(a[116] & b[220])^(a[115] & b[221])^(a[114] & b[222])^(a[113] & b[223])^(a[112] & b[224])^(a[111] & b[225])^(a[110] & b[226])^(a[109] & b[227])^(a[108] & b[228])^(a[107] & b[229])^(a[106] & b[230])^(a[105] & b[231])^(a[104] & b[232]);
assign y[337] = (a[232] & b[105])^(a[231] & b[106])^(a[230] & b[107])^(a[229] & b[108])^(a[228] & b[109])^(a[227] & b[110])^(a[226] & b[111])^(a[225] & b[112])^(a[224] & b[113])^(a[223] & b[114])^(a[222] & b[115])^(a[221] & b[116])^(a[220] & b[117])^(a[219] & b[118])^(a[218] & b[119])^(a[217] & b[120])^(a[216] & b[121])^(a[215] & b[122])^(a[214] & b[123])^(a[213] & b[124])^(a[212] & b[125])^(a[211] & b[126])^(a[210] & b[127])^(a[209] & b[128])^(a[208] & b[129])^(a[207] & b[130])^(a[206] & b[131])^(a[205] & b[132])^(a[204] & b[133])^(a[203] & b[134])^(a[202] & b[135])^(a[201] & b[136])^(a[200] & b[137])^(a[199] & b[138])^(a[198] & b[139])^(a[197] & b[140])^(a[196] & b[141])^(a[195] & b[142])^(a[194] & b[143])^(a[193] & b[144])^(a[192] & b[145])^(a[191] & b[146])^(a[190] & b[147])^(a[189] & b[148])^(a[188] & b[149])^(a[187] & b[150])^(a[186] & b[151])^(a[185] & b[152])^(a[184] & b[153])^(a[183] & b[154])^(a[182] & b[155])^(a[181] & b[156])^(a[180] & b[157])^(a[179] & b[158])^(a[178] & b[159])^(a[177] & b[160])^(a[176] & b[161])^(a[175] & b[162])^(a[174] & b[163])^(a[173] & b[164])^(a[172] & b[165])^(a[171] & b[166])^(a[170] & b[167])^(a[169] & b[168])^(a[168] & b[169])^(a[167] & b[170])^(a[166] & b[171])^(a[165] & b[172])^(a[164] & b[173])^(a[163] & b[174])^(a[162] & b[175])^(a[161] & b[176])^(a[160] & b[177])^(a[159] & b[178])^(a[158] & b[179])^(a[157] & b[180])^(a[156] & b[181])^(a[155] & b[182])^(a[154] & b[183])^(a[153] & b[184])^(a[152] & b[185])^(a[151] & b[186])^(a[150] & b[187])^(a[149] & b[188])^(a[148] & b[189])^(a[147] & b[190])^(a[146] & b[191])^(a[145] & b[192])^(a[144] & b[193])^(a[143] & b[194])^(a[142] & b[195])^(a[141] & b[196])^(a[140] & b[197])^(a[139] & b[198])^(a[138] & b[199])^(a[137] & b[200])^(a[136] & b[201])^(a[135] & b[202])^(a[134] & b[203])^(a[133] & b[204])^(a[132] & b[205])^(a[131] & b[206])^(a[130] & b[207])^(a[129] & b[208])^(a[128] & b[209])^(a[127] & b[210])^(a[126] & b[211])^(a[125] & b[212])^(a[124] & b[213])^(a[123] & b[214])^(a[122] & b[215])^(a[121] & b[216])^(a[120] & b[217])^(a[119] & b[218])^(a[118] & b[219])^(a[117] & b[220])^(a[116] & b[221])^(a[115] & b[222])^(a[114] & b[223])^(a[113] & b[224])^(a[112] & b[225])^(a[111] & b[226])^(a[110] & b[227])^(a[109] & b[228])^(a[108] & b[229])^(a[107] & b[230])^(a[106] & b[231])^(a[105] & b[232]);
assign y[338] = (a[232] & b[106])^(a[231] & b[107])^(a[230] & b[108])^(a[229] & b[109])^(a[228] & b[110])^(a[227] & b[111])^(a[226] & b[112])^(a[225] & b[113])^(a[224] & b[114])^(a[223] & b[115])^(a[222] & b[116])^(a[221] & b[117])^(a[220] & b[118])^(a[219] & b[119])^(a[218] & b[120])^(a[217] & b[121])^(a[216] & b[122])^(a[215] & b[123])^(a[214] & b[124])^(a[213] & b[125])^(a[212] & b[126])^(a[211] & b[127])^(a[210] & b[128])^(a[209] & b[129])^(a[208] & b[130])^(a[207] & b[131])^(a[206] & b[132])^(a[205] & b[133])^(a[204] & b[134])^(a[203] & b[135])^(a[202] & b[136])^(a[201] & b[137])^(a[200] & b[138])^(a[199] & b[139])^(a[198] & b[140])^(a[197] & b[141])^(a[196] & b[142])^(a[195] & b[143])^(a[194] & b[144])^(a[193] & b[145])^(a[192] & b[146])^(a[191] & b[147])^(a[190] & b[148])^(a[189] & b[149])^(a[188] & b[150])^(a[187] & b[151])^(a[186] & b[152])^(a[185] & b[153])^(a[184] & b[154])^(a[183] & b[155])^(a[182] & b[156])^(a[181] & b[157])^(a[180] & b[158])^(a[179] & b[159])^(a[178] & b[160])^(a[177] & b[161])^(a[176] & b[162])^(a[175] & b[163])^(a[174] & b[164])^(a[173] & b[165])^(a[172] & b[166])^(a[171] & b[167])^(a[170] & b[168])^(a[169] & b[169])^(a[168] & b[170])^(a[167] & b[171])^(a[166] & b[172])^(a[165] & b[173])^(a[164] & b[174])^(a[163] & b[175])^(a[162] & b[176])^(a[161] & b[177])^(a[160] & b[178])^(a[159] & b[179])^(a[158] & b[180])^(a[157] & b[181])^(a[156] & b[182])^(a[155] & b[183])^(a[154] & b[184])^(a[153] & b[185])^(a[152] & b[186])^(a[151] & b[187])^(a[150] & b[188])^(a[149] & b[189])^(a[148] & b[190])^(a[147] & b[191])^(a[146] & b[192])^(a[145] & b[193])^(a[144] & b[194])^(a[143] & b[195])^(a[142] & b[196])^(a[141] & b[197])^(a[140] & b[198])^(a[139] & b[199])^(a[138] & b[200])^(a[137] & b[201])^(a[136] & b[202])^(a[135] & b[203])^(a[134] & b[204])^(a[133] & b[205])^(a[132] & b[206])^(a[131] & b[207])^(a[130] & b[208])^(a[129] & b[209])^(a[128] & b[210])^(a[127] & b[211])^(a[126] & b[212])^(a[125] & b[213])^(a[124] & b[214])^(a[123] & b[215])^(a[122] & b[216])^(a[121] & b[217])^(a[120] & b[218])^(a[119] & b[219])^(a[118] & b[220])^(a[117] & b[221])^(a[116] & b[222])^(a[115] & b[223])^(a[114] & b[224])^(a[113] & b[225])^(a[112] & b[226])^(a[111] & b[227])^(a[110] & b[228])^(a[109] & b[229])^(a[108] & b[230])^(a[107] & b[231])^(a[106] & b[232]);
assign y[339] = (a[232] & b[107])^(a[231] & b[108])^(a[230] & b[109])^(a[229] & b[110])^(a[228] & b[111])^(a[227] & b[112])^(a[226] & b[113])^(a[225] & b[114])^(a[224] & b[115])^(a[223] & b[116])^(a[222] & b[117])^(a[221] & b[118])^(a[220] & b[119])^(a[219] & b[120])^(a[218] & b[121])^(a[217] & b[122])^(a[216] & b[123])^(a[215] & b[124])^(a[214] & b[125])^(a[213] & b[126])^(a[212] & b[127])^(a[211] & b[128])^(a[210] & b[129])^(a[209] & b[130])^(a[208] & b[131])^(a[207] & b[132])^(a[206] & b[133])^(a[205] & b[134])^(a[204] & b[135])^(a[203] & b[136])^(a[202] & b[137])^(a[201] & b[138])^(a[200] & b[139])^(a[199] & b[140])^(a[198] & b[141])^(a[197] & b[142])^(a[196] & b[143])^(a[195] & b[144])^(a[194] & b[145])^(a[193] & b[146])^(a[192] & b[147])^(a[191] & b[148])^(a[190] & b[149])^(a[189] & b[150])^(a[188] & b[151])^(a[187] & b[152])^(a[186] & b[153])^(a[185] & b[154])^(a[184] & b[155])^(a[183] & b[156])^(a[182] & b[157])^(a[181] & b[158])^(a[180] & b[159])^(a[179] & b[160])^(a[178] & b[161])^(a[177] & b[162])^(a[176] & b[163])^(a[175] & b[164])^(a[174] & b[165])^(a[173] & b[166])^(a[172] & b[167])^(a[171] & b[168])^(a[170] & b[169])^(a[169] & b[170])^(a[168] & b[171])^(a[167] & b[172])^(a[166] & b[173])^(a[165] & b[174])^(a[164] & b[175])^(a[163] & b[176])^(a[162] & b[177])^(a[161] & b[178])^(a[160] & b[179])^(a[159] & b[180])^(a[158] & b[181])^(a[157] & b[182])^(a[156] & b[183])^(a[155] & b[184])^(a[154] & b[185])^(a[153] & b[186])^(a[152] & b[187])^(a[151] & b[188])^(a[150] & b[189])^(a[149] & b[190])^(a[148] & b[191])^(a[147] & b[192])^(a[146] & b[193])^(a[145] & b[194])^(a[144] & b[195])^(a[143] & b[196])^(a[142] & b[197])^(a[141] & b[198])^(a[140] & b[199])^(a[139] & b[200])^(a[138] & b[201])^(a[137] & b[202])^(a[136] & b[203])^(a[135] & b[204])^(a[134] & b[205])^(a[133] & b[206])^(a[132] & b[207])^(a[131] & b[208])^(a[130] & b[209])^(a[129] & b[210])^(a[128] & b[211])^(a[127] & b[212])^(a[126] & b[213])^(a[125] & b[214])^(a[124] & b[215])^(a[123] & b[216])^(a[122] & b[217])^(a[121] & b[218])^(a[120] & b[219])^(a[119] & b[220])^(a[118] & b[221])^(a[117] & b[222])^(a[116] & b[223])^(a[115] & b[224])^(a[114] & b[225])^(a[113] & b[226])^(a[112] & b[227])^(a[111] & b[228])^(a[110] & b[229])^(a[109] & b[230])^(a[108] & b[231])^(a[107] & b[232]);
assign y[340] = (a[232] & b[108])^(a[231] & b[109])^(a[230] & b[110])^(a[229] & b[111])^(a[228] & b[112])^(a[227] & b[113])^(a[226] & b[114])^(a[225] & b[115])^(a[224] & b[116])^(a[223] & b[117])^(a[222] & b[118])^(a[221] & b[119])^(a[220] & b[120])^(a[219] & b[121])^(a[218] & b[122])^(a[217] & b[123])^(a[216] & b[124])^(a[215] & b[125])^(a[214] & b[126])^(a[213] & b[127])^(a[212] & b[128])^(a[211] & b[129])^(a[210] & b[130])^(a[209] & b[131])^(a[208] & b[132])^(a[207] & b[133])^(a[206] & b[134])^(a[205] & b[135])^(a[204] & b[136])^(a[203] & b[137])^(a[202] & b[138])^(a[201] & b[139])^(a[200] & b[140])^(a[199] & b[141])^(a[198] & b[142])^(a[197] & b[143])^(a[196] & b[144])^(a[195] & b[145])^(a[194] & b[146])^(a[193] & b[147])^(a[192] & b[148])^(a[191] & b[149])^(a[190] & b[150])^(a[189] & b[151])^(a[188] & b[152])^(a[187] & b[153])^(a[186] & b[154])^(a[185] & b[155])^(a[184] & b[156])^(a[183] & b[157])^(a[182] & b[158])^(a[181] & b[159])^(a[180] & b[160])^(a[179] & b[161])^(a[178] & b[162])^(a[177] & b[163])^(a[176] & b[164])^(a[175] & b[165])^(a[174] & b[166])^(a[173] & b[167])^(a[172] & b[168])^(a[171] & b[169])^(a[170] & b[170])^(a[169] & b[171])^(a[168] & b[172])^(a[167] & b[173])^(a[166] & b[174])^(a[165] & b[175])^(a[164] & b[176])^(a[163] & b[177])^(a[162] & b[178])^(a[161] & b[179])^(a[160] & b[180])^(a[159] & b[181])^(a[158] & b[182])^(a[157] & b[183])^(a[156] & b[184])^(a[155] & b[185])^(a[154] & b[186])^(a[153] & b[187])^(a[152] & b[188])^(a[151] & b[189])^(a[150] & b[190])^(a[149] & b[191])^(a[148] & b[192])^(a[147] & b[193])^(a[146] & b[194])^(a[145] & b[195])^(a[144] & b[196])^(a[143] & b[197])^(a[142] & b[198])^(a[141] & b[199])^(a[140] & b[200])^(a[139] & b[201])^(a[138] & b[202])^(a[137] & b[203])^(a[136] & b[204])^(a[135] & b[205])^(a[134] & b[206])^(a[133] & b[207])^(a[132] & b[208])^(a[131] & b[209])^(a[130] & b[210])^(a[129] & b[211])^(a[128] & b[212])^(a[127] & b[213])^(a[126] & b[214])^(a[125] & b[215])^(a[124] & b[216])^(a[123] & b[217])^(a[122] & b[218])^(a[121] & b[219])^(a[120] & b[220])^(a[119] & b[221])^(a[118] & b[222])^(a[117] & b[223])^(a[116] & b[224])^(a[115] & b[225])^(a[114] & b[226])^(a[113] & b[227])^(a[112] & b[228])^(a[111] & b[229])^(a[110] & b[230])^(a[109] & b[231])^(a[108] & b[232]);
assign y[341] = (a[232] & b[109])^(a[231] & b[110])^(a[230] & b[111])^(a[229] & b[112])^(a[228] & b[113])^(a[227] & b[114])^(a[226] & b[115])^(a[225] & b[116])^(a[224] & b[117])^(a[223] & b[118])^(a[222] & b[119])^(a[221] & b[120])^(a[220] & b[121])^(a[219] & b[122])^(a[218] & b[123])^(a[217] & b[124])^(a[216] & b[125])^(a[215] & b[126])^(a[214] & b[127])^(a[213] & b[128])^(a[212] & b[129])^(a[211] & b[130])^(a[210] & b[131])^(a[209] & b[132])^(a[208] & b[133])^(a[207] & b[134])^(a[206] & b[135])^(a[205] & b[136])^(a[204] & b[137])^(a[203] & b[138])^(a[202] & b[139])^(a[201] & b[140])^(a[200] & b[141])^(a[199] & b[142])^(a[198] & b[143])^(a[197] & b[144])^(a[196] & b[145])^(a[195] & b[146])^(a[194] & b[147])^(a[193] & b[148])^(a[192] & b[149])^(a[191] & b[150])^(a[190] & b[151])^(a[189] & b[152])^(a[188] & b[153])^(a[187] & b[154])^(a[186] & b[155])^(a[185] & b[156])^(a[184] & b[157])^(a[183] & b[158])^(a[182] & b[159])^(a[181] & b[160])^(a[180] & b[161])^(a[179] & b[162])^(a[178] & b[163])^(a[177] & b[164])^(a[176] & b[165])^(a[175] & b[166])^(a[174] & b[167])^(a[173] & b[168])^(a[172] & b[169])^(a[171] & b[170])^(a[170] & b[171])^(a[169] & b[172])^(a[168] & b[173])^(a[167] & b[174])^(a[166] & b[175])^(a[165] & b[176])^(a[164] & b[177])^(a[163] & b[178])^(a[162] & b[179])^(a[161] & b[180])^(a[160] & b[181])^(a[159] & b[182])^(a[158] & b[183])^(a[157] & b[184])^(a[156] & b[185])^(a[155] & b[186])^(a[154] & b[187])^(a[153] & b[188])^(a[152] & b[189])^(a[151] & b[190])^(a[150] & b[191])^(a[149] & b[192])^(a[148] & b[193])^(a[147] & b[194])^(a[146] & b[195])^(a[145] & b[196])^(a[144] & b[197])^(a[143] & b[198])^(a[142] & b[199])^(a[141] & b[200])^(a[140] & b[201])^(a[139] & b[202])^(a[138] & b[203])^(a[137] & b[204])^(a[136] & b[205])^(a[135] & b[206])^(a[134] & b[207])^(a[133] & b[208])^(a[132] & b[209])^(a[131] & b[210])^(a[130] & b[211])^(a[129] & b[212])^(a[128] & b[213])^(a[127] & b[214])^(a[126] & b[215])^(a[125] & b[216])^(a[124] & b[217])^(a[123] & b[218])^(a[122] & b[219])^(a[121] & b[220])^(a[120] & b[221])^(a[119] & b[222])^(a[118] & b[223])^(a[117] & b[224])^(a[116] & b[225])^(a[115] & b[226])^(a[114] & b[227])^(a[113] & b[228])^(a[112] & b[229])^(a[111] & b[230])^(a[110] & b[231])^(a[109] & b[232]);
assign y[342] = (a[232] & b[110])^(a[231] & b[111])^(a[230] & b[112])^(a[229] & b[113])^(a[228] & b[114])^(a[227] & b[115])^(a[226] & b[116])^(a[225] & b[117])^(a[224] & b[118])^(a[223] & b[119])^(a[222] & b[120])^(a[221] & b[121])^(a[220] & b[122])^(a[219] & b[123])^(a[218] & b[124])^(a[217] & b[125])^(a[216] & b[126])^(a[215] & b[127])^(a[214] & b[128])^(a[213] & b[129])^(a[212] & b[130])^(a[211] & b[131])^(a[210] & b[132])^(a[209] & b[133])^(a[208] & b[134])^(a[207] & b[135])^(a[206] & b[136])^(a[205] & b[137])^(a[204] & b[138])^(a[203] & b[139])^(a[202] & b[140])^(a[201] & b[141])^(a[200] & b[142])^(a[199] & b[143])^(a[198] & b[144])^(a[197] & b[145])^(a[196] & b[146])^(a[195] & b[147])^(a[194] & b[148])^(a[193] & b[149])^(a[192] & b[150])^(a[191] & b[151])^(a[190] & b[152])^(a[189] & b[153])^(a[188] & b[154])^(a[187] & b[155])^(a[186] & b[156])^(a[185] & b[157])^(a[184] & b[158])^(a[183] & b[159])^(a[182] & b[160])^(a[181] & b[161])^(a[180] & b[162])^(a[179] & b[163])^(a[178] & b[164])^(a[177] & b[165])^(a[176] & b[166])^(a[175] & b[167])^(a[174] & b[168])^(a[173] & b[169])^(a[172] & b[170])^(a[171] & b[171])^(a[170] & b[172])^(a[169] & b[173])^(a[168] & b[174])^(a[167] & b[175])^(a[166] & b[176])^(a[165] & b[177])^(a[164] & b[178])^(a[163] & b[179])^(a[162] & b[180])^(a[161] & b[181])^(a[160] & b[182])^(a[159] & b[183])^(a[158] & b[184])^(a[157] & b[185])^(a[156] & b[186])^(a[155] & b[187])^(a[154] & b[188])^(a[153] & b[189])^(a[152] & b[190])^(a[151] & b[191])^(a[150] & b[192])^(a[149] & b[193])^(a[148] & b[194])^(a[147] & b[195])^(a[146] & b[196])^(a[145] & b[197])^(a[144] & b[198])^(a[143] & b[199])^(a[142] & b[200])^(a[141] & b[201])^(a[140] & b[202])^(a[139] & b[203])^(a[138] & b[204])^(a[137] & b[205])^(a[136] & b[206])^(a[135] & b[207])^(a[134] & b[208])^(a[133] & b[209])^(a[132] & b[210])^(a[131] & b[211])^(a[130] & b[212])^(a[129] & b[213])^(a[128] & b[214])^(a[127] & b[215])^(a[126] & b[216])^(a[125] & b[217])^(a[124] & b[218])^(a[123] & b[219])^(a[122] & b[220])^(a[121] & b[221])^(a[120] & b[222])^(a[119] & b[223])^(a[118] & b[224])^(a[117] & b[225])^(a[116] & b[226])^(a[115] & b[227])^(a[114] & b[228])^(a[113] & b[229])^(a[112] & b[230])^(a[111] & b[231])^(a[110] & b[232]);
assign y[343] = (a[232] & b[111])^(a[231] & b[112])^(a[230] & b[113])^(a[229] & b[114])^(a[228] & b[115])^(a[227] & b[116])^(a[226] & b[117])^(a[225] & b[118])^(a[224] & b[119])^(a[223] & b[120])^(a[222] & b[121])^(a[221] & b[122])^(a[220] & b[123])^(a[219] & b[124])^(a[218] & b[125])^(a[217] & b[126])^(a[216] & b[127])^(a[215] & b[128])^(a[214] & b[129])^(a[213] & b[130])^(a[212] & b[131])^(a[211] & b[132])^(a[210] & b[133])^(a[209] & b[134])^(a[208] & b[135])^(a[207] & b[136])^(a[206] & b[137])^(a[205] & b[138])^(a[204] & b[139])^(a[203] & b[140])^(a[202] & b[141])^(a[201] & b[142])^(a[200] & b[143])^(a[199] & b[144])^(a[198] & b[145])^(a[197] & b[146])^(a[196] & b[147])^(a[195] & b[148])^(a[194] & b[149])^(a[193] & b[150])^(a[192] & b[151])^(a[191] & b[152])^(a[190] & b[153])^(a[189] & b[154])^(a[188] & b[155])^(a[187] & b[156])^(a[186] & b[157])^(a[185] & b[158])^(a[184] & b[159])^(a[183] & b[160])^(a[182] & b[161])^(a[181] & b[162])^(a[180] & b[163])^(a[179] & b[164])^(a[178] & b[165])^(a[177] & b[166])^(a[176] & b[167])^(a[175] & b[168])^(a[174] & b[169])^(a[173] & b[170])^(a[172] & b[171])^(a[171] & b[172])^(a[170] & b[173])^(a[169] & b[174])^(a[168] & b[175])^(a[167] & b[176])^(a[166] & b[177])^(a[165] & b[178])^(a[164] & b[179])^(a[163] & b[180])^(a[162] & b[181])^(a[161] & b[182])^(a[160] & b[183])^(a[159] & b[184])^(a[158] & b[185])^(a[157] & b[186])^(a[156] & b[187])^(a[155] & b[188])^(a[154] & b[189])^(a[153] & b[190])^(a[152] & b[191])^(a[151] & b[192])^(a[150] & b[193])^(a[149] & b[194])^(a[148] & b[195])^(a[147] & b[196])^(a[146] & b[197])^(a[145] & b[198])^(a[144] & b[199])^(a[143] & b[200])^(a[142] & b[201])^(a[141] & b[202])^(a[140] & b[203])^(a[139] & b[204])^(a[138] & b[205])^(a[137] & b[206])^(a[136] & b[207])^(a[135] & b[208])^(a[134] & b[209])^(a[133] & b[210])^(a[132] & b[211])^(a[131] & b[212])^(a[130] & b[213])^(a[129] & b[214])^(a[128] & b[215])^(a[127] & b[216])^(a[126] & b[217])^(a[125] & b[218])^(a[124] & b[219])^(a[123] & b[220])^(a[122] & b[221])^(a[121] & b[222])^(a[120] & b[223])^(a[119] & b[224])^(a[118] & b[225])^(a[117] & b[226])^(a[116] & b[227])^(a[115] & b[228])^(a[114] & b[229])^(a[113] & b[230])^(a[112] & b[231])^(a[111] & b[232]);
assign y[344] = (a[232] & b[112])^(a[231] & b[113])^(a[230] & b[114])^(a[229] & b[115])^(a[228] & b[116])^(a[227] & b[117])^(a[226] & b[118])^(a[225] & b[119])^(a[224] & b[120])^(a[223] & b[121])^(a[222] & b[122])^(a[221] & b[123])^(a[220] & b[124])^(a[219] & b[125])^(a[218] & b[126])^(a[217] & b[127])^(a[216] & b[128])^(a[215] & b[129])^(a[214] & b[130])^(a[213] & b[131])^(a[212] & b[132])^(a[211] & b[133])^(a[210] & b[134])^(a[209] & b[135])^(a[208] & b[136])^(a[207] & b[137])^(a[206] & b[138])^(a[205] & b[139])^(a[204] & b[140])^(a[203] & b[141])^(a[202] & b[142])^(a[201] & b[143])^(a[200] & b[144])^(a[199] & b[145])^(a[198] & b[146])^(a[197] & b[147])^(a[196] & b[148])^(a[195] & b[149])^(a[194] & b[150])^(a[193] & b[151])^(a[192] & b[152])^(a[191] & b[153])^(a[190] & b[154])^(a[189] & b[155])^(a[188] & b[156])^(a[187] & b[157])^(a[186] & b[158])^(a[185] & b[159])^(a[184] & b[160])^(a[183] & b[161])^(a[182] & b[162])^(a[181] & b[163])^(a[180] & b[164])^(a[179] & b[165])^(a[178] & b[166])^(a[177] & b[167])^(a[176] & b[168])^(a[175] & b[169])^(a[174] & b[170])^(a[173] & b[171])^(a[172] & b[172])^(a[171] & b[173])^(a[170] & b[174])^(a[169] & b[175])^(a[168] & b[176])^(a[167] & b[177])^(a[166] & b[178])^(a[165] & b[179])^(a[164] & b[180])^(a[163] & b[181])^(a[162] & b[182])^(a[161] & b[183])^(a[160] & b[184])^(a[159] & b[185])^(a[158] & b[186])^(a[157] & b[187])^(a[156] & b[188])^(a[155] & b[189])^(a[154] & b[190])^(a[153] & b[191])^(a[152] & b[192])^(a[151] & b[193])^(a[150] & b[194])^(a[149] & b[195])^(a[148] & b[196])^(a[147] & b[197])^(a[146] & b[198])^(a[145] & b[199])^(a[144] & b[200])^(a[143] & b[201])^(a[142] & b[202])^(a[141] & b[203])^(a[140] & b[204])^(a[139] & b[205])^(a[138] & b[206])^(a[137] & b[207])^(a[136] & b[208])^(a[135] & b[209])^(a[134] & b[210])^(a[133] & b[211])^(a[132] & b[212])^(a[131] & b[213])^(a[130] & b[214])^(a[129] & b[215])^(a[128] & b[216])^(a[127] & b[217])^(a[126] & b[218])^(a[125] & b[219])^(a[124] & b[220])^(a[123] & b[221])^(a[122] & b[222])^(a[121] & b[223])^(a[120] & b[224])^(a[119] & b[225])^(a[118] & b[226])^(a[117] & b[227])^(a[116] & b[228])^(a[115] & b[229])^(a[114] & b[230])^(a[113] & b[231])^(a[112] & b[232]);
assign y[345] = (a[232] & b[113])^(a[231] & b[114])^(a[230] & b[115])^(a[229] & b[116])^(a[228] & b[117])^(a[227] & b[118])^(a[226] & b[119])^(a[225] & b[120])^(a[224] & b[121])^(a[223] & b[122])^(a[222] & b[123])^(a[221] & b[124])^(a[220] & b[125])^(a[219] & b[126])^(a[218] & b[127])^(a[217] & b[128])^(a[216] & b[129])^(a[215] & b[130])^(a[214] & b[131])^(a[213] & b[132])^(a[212] & b[133])^(a[211] & b[134])^(a[210] & b[135])^(a[209] & b[136])^(a[208] & b[137])^(a[207] & b[138])^(a[206] & b[139])^(a[205] & b[140])^(a[204] & b[141])^(a[203] & b[142])^(a[202] & b[143])^(a[201] & b[144])^(a[200] & b[145])^(a[199] & b[146])^(a[198] & b[147])^(a[197] & b[148])^(a[196] & b[149])^(a[195] & b[150])^(a[194] & b[151])^(a[193] & b[152])^(a[192] & b[153])^(a[191] & b[154])^(a[190] & b[155])^(a[189] & b[156])^(a[188] & b[157])^(a[187] & b[158])^(a[186] & b[159])^(a[185] & b[160])^(a[184] & b[161])^(a[183] & b[162])^(a[182] & b[163])^(a[181] & b[164])^(a[180] & b[165])^(a[179] & b[166])^(a[178] & b[167])^(a[177] & b[168])^(a[176] & b[169])^(a[175] & b[170])^(a[174] & b[171])^(a[173] & b[172])^(a[172] & b[173])^(a[171] & b[174])^(a[170] & b[175])^(a[169] & b[176])^(a[168] & b[177])^(a[167] & b[178])^(a[166] & b[179])^(a[165] & b[180])^(a[164] & b[181])^(a[163] & b[182])^(a[162] & b[183])^(a[161] & b[184])^(a[160] & b[185])^(a[159] & b[186])^(a[158] & b[187])^(a[157] & b[188])^(a[156] & b[189])^(a[155] & b[190])^(a[154] & b[191])^(a[153] & b[192])^(a[152] & b[193])^(a[151] & b[194])^(a[150] & b[195])^(a[149] & b[196])^(a[148] & b[197])^(a[147] & b[198])^(a[146] & b[199])^(a[145] & b[200])^(a[144] & b[201])^(a[143] & b[202])^(a[142] & b[203])^(a[141] & b[204])^(a[140] & b[205])^(a[139] & b[206])^(a[138] & b[207])^(a[137] & b[208])^(a[136] & b[209])^(a[135] & b[210])^(a[134] & b[211])^(a[133] & b[212])^(a[132] & b[213])^(a[131] & b[214])^(a[130] & b[215])^(a[129] & b[216])^(a[128] & b[217])^(a[127] & b[218])^(a[126] & b[219])^(a[125] & b[220])^(a[124] & b[221])^(a[123] & b[222])^(a[122] & b[223])^(a[121] & b[224])^(a[120] & b[225])^(a[119] & b[226])^(a[118] & b[227])^(a[117] & b[228])^(a[116] & b[229])^(a[115] & b[230])^(a[114] & b[231])^(a[113] & b[232]);
assign y[346] = (a[232] & b[114])^(a[231] & b[115])^(a[230] & b[116])^(a[229] & b[117])^(a[228] & b[118])^(a[227] & b[119])^(a[226] & b[120])^(a[225] & b[121])^(a[224] & b[122])^(a[223] & b[123])^(a[222] & b[124])^(a[221] & b[125])^(a[220] & b[126])^(a[219] & b[127])^(a[218] & b[128])^(a[217] & b[129])^(a[216] & b[130])^(a[215] & b[131])^(a[214] & b[132])^(a[213] & b[133])^(a[212] & b[134])^(a[211] & b[135])^(a[210] & b[136])^(a[209] & b[137])^(a[208] & b[138])^(a[207] & b[139])^(a[206] & b[140])^(a[205] & b[141])^(a[204] & b[142])^(a[203] & b[143])^(a[202] & b[144])^(a[201] & b[145])^(a[200] & b[146])^(a[199] & b[147])^(a[198] & b[148])^(a[197] & b[149])^(a[196] & b[150])^(a[195] & b[151])^(a[194] & b[152])^(a[193] & b[153])^(a[192] & b[154])^(a[191] & b[155])^(a[190] & b[156])^(a[189] & b[157])^(a[188] & b[158])^(a[187] & b[159])^(a[186] & b[160])^(a[185] & b[161])^(a[184] & b[162])^(a[183] & b[163])^(a[182] & b[164])^(a[181] & b[165])^(a[180] & b[166])^(a[179] & b[167])^(a[178] & b[168])^(a[177] & b[169])^(a[176] & b[170])^(a[175] & b[171])^(a[174] & b[172])^(a[173] & b[173])^(a[172] & b[174])^(a[171] & b[175])^(a[170] & b[176])^(a[169] & b[177])^(a[168] & b[178])^(a[167] & b[179])^(a[166] & b[180])^(a[165] & b[181])^(a[164] & b[182])^(a[163] & b[183])^(a[162] & b[184])^(a[161] & b[185])^(a[160] & b[186])^(a[159] & b[187])^(a[158] & b[188])^(a[157] & b[189])^(a[156] & b[190])^(a[155] & b[191])^(a[154] & b[192])^(a[153] & b[193])^(a[152] & b[194])^(a[151] & b[195])^(a[150] & b[196])^(a[149] & b[197])^(a[148] & b[198])^(a[147] & b[199])^(a[146] & b[200])^(a[145] & b[201])^(a[144] & b[202])^(a[143] & b[203])^(a[142] & b[204])^(a[141] & b[205])^(a[140] & b[206])^(a[139] & b[207])^(a[138] & b[208])^(a[137] & b[209])^(a[136] & b[210])^(a[135] & b[211])^(a[134] & b[212])^(a[133] & b[213])^(a[132] & b[214])^(a[131] & b[215])^(a[130] & b[216])^(a[129] & b[217])^(a[128] & b[218])^(a[127] & b[219])^(a[126] & b[220])^(a[125] & b[221])^(a[124] & b[222])^(a[123] & b[223])^(a[122] & b[224])^(a[121] & b[225])^(a[120] & b[226])^(a[119] & b[227])^(a[118] & b[228])^(a[117] & b[229])^(a[116] & b[230])^(a[115] & b[231])^(a[114] & b[232]);
assign y[347] = (a[232] & b[115])^(a[231] & b[116])^(a[230] & b[117])^(a[229] & b[118])^(a[228] & b[119])^(a[227] & b[120])^(a[226] & b[121])^(a[225] & b[122])^(a[224] & b[123])^(a[223] & b[124])^(a[222] & b[125])^(a[221] & b[126])^(a[220] & b[127])^(a[219] & b[128])^(a[218] & b[129])^(a[217] & b[130])^(a[216] & b[131])^(a[215] & b[132])^(a[214] & b[133])^(a[213] & b[134])^(a[212] & b[135])^(a[211] & b[136])^(a[210] & b[137])^(a[209] & b[138])^(a[208] & b[139])^(a[207] & b[140])^(a[206] & b[141])^(a[205] & b[142])^(a[204] & b[143])^(a[203] & b[144])^(a[202] & b[145])^(a[201] & b[146])^(a[200] & b[147])^(a[199] & b[148])^(a[198] & b[149])^(a[197] & b[150])^(a[196] & b[151])^(a[195] & b[152])^(a[194] & b[153])^(a[193] & b[154])^(a[192] & b[155])^(a[191] & b[156])^(a[190] & b[157])^(a[189] & b[158])^(a[188] & b[159])^(a[187] & b[160])^(a[186] & b[161])^(a[185] & b[162])^(a[184] & b[163])^(a[183] & b[164])^(a[182] & b[165])^(a[181] & b[166])^(a[180] & b[167])^(a[179] & b[168])^(a[178] & b[169])^(a[177] & b[170])^(a[176] & b[171])^(a[175] & b[172])^(a[174] & b[173])^(a[173] & b[174])^(a[172] & b[175])^(a[171] & b[176])^(a[170] & b[177])^(a[169] & b[178])^(a[168] & b[179])^(a[167] & b[180])^(a[166] & b[181])^(a[165] & b[182])^(a[164] & b[183])^(a[163] & b[184])^(a[162] & b[185])^(a[161] & b[186])^(a[160] & b[187])^(a[159] & b[188])^(a[158] & b[189])^(a[157] & b[190])^(a[156] & b[191])^(a[155] & b[192])^(a[154] & b[193])^(a[153] & b[194])^(a[152] & b[195])^(a[151] & b[196])^(a[150] & b[197])^(a[149] & b[198])^(a[148] & b[199])^(a[147] & b[200])^(a[146] & b[201])^(a[145] & b[202])^(a[144] & b[203])^(a[143] & b[204])^(a[142] & b[205])^(a[141] & b[206])^(a[140] & b[207])^(a[139] & b[208])^(a[138] & b[209])^(a[137] & b[210])^(a[136] & b[211])^(a[135] & b[212])^(a[134] & b[213])^(a[133] & b[214])^(a[132] & b[215])^(a[131] & b[216])^(a[130] & b[217])^(a[129] & b[218])^(a[128] & b[219])^(a[127] & b[220])^(a[126] & b[221])^(a[125] & b[222])^(a[124] & b[223])^(a[123] & b[224])^(a[122] & b[225])^(a[121] & b[226])^(a[120] & b[227])^(a[119] & b[228])^(a[118] & b[229])^(a[117] & b[230])^(a[116] & b[231])^(a[115] & b[232]);
assign y[348] = (a[232] & b[116])^(a[231] & b[117])^(a[230] & b[118])^(a[229] & b[119])^(a[228] & b[120])^(a[227] & b[121])^(a[226] & b[122])^(a[225] & b[123])^(a[224] & b[124])^(a[223] & b[125])^(a[222] & b[126])^(a[221] & b[127])^(a[220] & b[128])^(a[219] & b[129])^(a[218] & b[130])^(a[217] & b[131])^(a[216] & b[132])^(a[215] & b[133])^(a[214] & b[134])^(a[213] & b[135])^(a[212] & b[136])^(a[211] & b[137])^(a[210] & b[138])^(a[209] & b[139])^(a[208] & b[140])^(a[207] & b[141])^(a[206] & b[142])^(a[205] & b[143])^(a[204] & b[144])^(a[203] & b[145])^(a[202] & b[146])^(a[201] & b[147])^(a[200] & b[148])^(a[199] & b[149])^(a[198] & b[150])^(a[197] & b[151])^(a[196] & b[152])^(a[195] & b[153])^(a[194] & b[154])^(a[193] & b[155])^(a[192] & b[156])^(a[191] & b[157])^(a[190] & b[158])^(a[189] & b[159])^(a[188] & b[160])^(a[187] & b[161])^(a[186] & b[162])^(a[185] & b[163])^(a[184] & b[164])^(a[183] & b[165])^(a[182] & b[166])^(a[181] & b[167])^(a[180] & b[168])^(a[179] & b[169])^(a[178] & b[170])^(a[177] & b[171])^(a[176] & b[172])^(a[175] & b[173])^(a[174] & b[174])^(a[173] & b[175])^(a[172] & b[176])^(a[171] & b[177])^(a[170] & b[178])^(a[169] & b[179])^(a[168] & b[180])^(a[167] & b[181])^(a[166] & b[182])^(a[165] & b[183])^(a[164] & b[184])^(a[163] & b[185])^(a[162] & b[186])^(a[161] & b[187])^(a[160] & b[188])^(a[159] & b[189])^(a[158] & b[190])^(a[157] & b[191])^(a[156] & b[192])^(a[155] & b[193])^(a[154] & b[194])^(a[153] & b[195])^(a[152] & b[196])^(a[151] & b[197])^(a[150] & b[198])^(a[149] & b[199])^(a[148] & b[200])^(a[147] & b[201])^(a[146] & b[202])^(a[145] & b[203])^(a[144] & b[204])^(a[143] & b[205])^(a[142] & b[206])^(a[141] & b[207])^(a[140] & b[208])^(a[139] & b[209])^(a[138] & b[210])^(a[137] & b[211])^(a[136] & b[212])^(a[135] & b[213])^(a[134] & b[214])^(a[133] & b[215])^(a[132] & b[216])^(a[131] & b[217])^(a[130] & b[218])^(a[129] & b[219])^(a[128] & b[220])^(a[127] & b[221])^(a[126] & b[222])^(a[125] & b[223])^(a[124] & b[224])^(a[123] & b[225])^(a[122] & b[226])^(a[121] & b[227])^(a[120] & b[228])^(a[119] & b[229])^(a[118] & b[230])^(a[117] & b[231])^(a[116] & b[232]);
assign y[349] = (a[232] & b[117])^(a[231] & b[118])^(a[230] & b[119])^(a[229] & b[120])^(a[228] & b[121])^(a[227] & b[122])^(a[226] & b[123])^(a[225] & b[124])^(a[224] & b[125])^(a[223] & b[126])^(a[222] & b[127])^(a[221] & b[128])^(a[220] & b[129])^(a[219] & b[130])^(a[218] & b[131])^(a[217] & b[132])^(a[216] & b[133])^(a[215] & b[134])^(a[214] & b[135])^(a[213] & b[136])^(a[212] & b[137])^(a[211] & b[138])^(a[210] & b[139])^(a[209] & b[140])^(a[208] & b[141])^(a[207] & b[142])^(a[206] & b[143])^(a[205] & b[144])^(a[204] & b[145])^(a[203] & b[146])^(a[202] & b[147])^(a[201] & b[148])^(a[200] & b[149])^(a[199] & b[150])^(a[198] & b[151])^(a[197] & b[152])^(a[196] & b[153])^(a[195] & b[154])^(a[194] & b[155])^(a[193] & b[156])^(a[192] & b[157])^(a[191] & b[158])^(a[190] & b[159])^(a[189] & b[160])^(a[188] & b[161])^(a[187] & b[162])^(a[186] & b[163])^(a[185] & b[164])^(a[184] & b[165])^(a[183] & b[166])^(a[182] & b[167])^(a[181] & b[168])^(a[180] & b[169])^(a[179] & b[170])^(a[178] & b[171])^(a[177] & b[172])^(a[176] & b[173])^(a[175] & b[174])^(a[174] & b[175])^(a[173] & b[176])^(a[172] & b[177])^(a[171] & b[178])^(a[170] & b[179])^(a[169] & b[180])^(a[168] & b[181])^(a[167] & b[182])^(a[166] & b[183])^(a[165] & b[184])^(a[164] & b[185])^(a[163] & b[186])^(a[162] & b[187])^(a[161] & b[188])^(a[160] & b[189])^(a[159] & b[190])^(a[158] & b[191])^(a[157] & b[192])^(a[156] & b[193])^(a[155] & b[194])^(a[154] & b[195])^(a[153] & b[196])^(a[152] & b[197])^(a[151] & b[198])^(a[150] & b[199])^(a[149] & b[200])^(a[148] & b[201])^(a[147] & b[202])^(a[146] & b[203])^(a[145] & b[204])^(a[144] & b[205])^(a[143] & b[206])^(a[142] & b[207])^(a[141] & b[208])^(a[140] & b[209])^(a[139] & b[210])^(a[138] & b[211])^(a[137] & b[212])^(a[136] & b[213])^(a[135] & b[214])^(a[134] & b[215])^(a[133] & b[216])^(a[132] & b[217])^(a[131] & b[218])^(a[130] & b[219])^(a[129] & b[220])^(a[128] & b[221])^(a[127] & b[222])^(a[126] & b[223])^(a[125] & b[224])^(a[124] & b[225])^(a[123] & b[226])^(a[122] & b[227])^(a[121] & b[228])^(a[120] & b[229])^(a[119] & b[230])^(a[118] & b[231])^(a[117] & b[232]);
assign y[350] = (a[232] & b[118])^(a[231] & b[119])^(a[230] & b[120])^(a[229] & b[121])^(a[228] & b[122])^(a[227] & b[123])^(a[226] & b[124])^(a[225] & b[125])^(a[224] & b[126])^(a[223] & b[127])^(a[222] & b[128])^(a[221] & b[129])^(a[220] & b[130])^(a[219] & b[131])^(a[218] & b[132])^(a[217] & b[133])^(a[216] & b[134])^(a[215] & b[135])^(a[214] & b[136])^(a[213] & b[137])^(a[212] & b[138])^(a[211] & b[139])^(a[210] & b[140])^(a[209] & b[141])^(a[208] & b[142])^(a[207] & b[143])^(a[206] & b[144])^(a[205] & b[145])^(a[204] & b[146])^(a[203] & b[147])^(a[202] & b[148])^(a[201] & b[149])^(a[200] & b[150])^(a[199] & b[151])^(a[198] & b[152])^(a[197] & b[153])^(a[196] & b[154])^(a[195] & b[155])^(a[194] & b[156])^(a[193] & b[157])^(a[192] & b[158])^(a[191] & b[159])^(a[190] & b[160])^(a[189] & b[161])^(a[188] & b[162])^(a[187] & b[163])^(a[186] & b[164])^(a[185] & b[165])^(a[184] & b[166])^(a[183] & b[167])^(a[182] & b[168])^(a[181] & b[169])^(a[180] & b[170])^(a[179] & b[171])^(a[178] & b[172])^(a[177] & b[173])^(a[176] & b[174])^(a[175] & b[175])^(a[174] & b[176])^(a[173] & b[177])^(a[172] & b[178])^(a[171] & b[179])^(a[170] & b[180])^(a[169] & b[181])^(a[168] & b[182])^(a[167] & b[183])^(a[166] & b[184])^(a[165] & b[185])^(a[164] & b[186])^(a[163] & b[187])^(a[162] & b[188])^(a[161] & b[189])^(a[160] & b[190])^(a[159] & b[191])^(a[158] & b[192])^(a[157] & b[193])^(a[156] & b[194])^(a[155] & b[195])^(a[154] & b[196])^(a[153] & b[197])^(a[152] & b[198])^(a[151] & b[199])^(a[150] & b[200])^(a[149] & b[201])^(a[148] & b[202])^(a[147] & b[203])^(a[146] & b[204])^(a[145] & b[205])^(a[144] & b[206])^(a[143] & b[207])^(a[142] & b[208])^(a[141] & b[209])^(a[140] & b[210])^(a[139] & b[211])^(a[138] & b[212])^(a[137] & b[213])^(a[136] & b[214])^(a[135] & b[215])^(a[134] & b[216])^(a[133] & b[217])^(a[132] & b[218])^(a[131] & b[219])^(a[130] & b[220])^(a[129] & b[221])^(a[128] & b[222])^(a[127] & b[223])^(a[126] & b[224])^(a[125] & b[225])^(a[124] & b[226])^(a[123] & b[227])^(a[122] & b[228])^(a[121] & b[229])^(a[120] & b[230])^(a[119] & b[231])^(a[118] & b[232]);
assign y[351] = (a[232] & b[119])^(a[231] & b[120])^(a[230] & b[121])^(a[229] & b[122])^(a[228] & b[123])^(a[227] & b[124])^(a[226] & b[125])^(a[225] & b[126])^(a[224] & b[127])^(a[223] & b[128])^(a[222] & b[129])^(a[221] & b[130])^(a[220] & b[131])^(a[219] & b[132])^(a[218] & b[133])^(a[217] & b[134])^(a[216] & b[135])^(a[215] & b[136])^(a[214] & b[137])^(a[213] & b[138])^(a[212] & b[139])^(a[211] & b[140])^(a[210] & b[141])^(a[209] & b[142])^(a[208] & b[143])^(a[207] & b[144])^(a[206] & b[145])^(a[205] & b[146])^(a[204] & b[147])^(a[203] & b[148])^(a[202] & b[149])^(a[201] & b[150])^(a[200] & b[151])^(a[199] & b[152])^(a[198] & b[153])^(a[197] & b[154])^(a[196] & b[155])^(a[195] & b[156])^(a[194] & b[157])^(a[193] & b[158])^(a[192] & b[159])^(a[191] & b[160])^(a[190] & b[161])^(a[189] & b[162])^(a[188] & b[163])^(a[187] & b[164])^(a[186] & b[165])^(a[185] & b[166])^(a[184] & b[167])^(a[183] & b[168])^(a[182] & b[169])^(a[181] & b[170])^(a[180] & b[171])^(a[179] & b[172])^(a[178] & b[173])^(a[177] & b[174])^(a[176] & b[175])^(a[175] & b[176])^(a[174] & b[177])^(a[173] & b[178])^(a[172] & b[179])^(a[171] & b[180])^(a[170] & b[181])^(a[169] & b[182])^(a[168] & b[183])^(a[167] & b[184])^(a[166] & b[185])^(a[165] & b[186])^(a[164] & b[187])^(a[163] & b[188])^(a[162] & b[189])^(a[161] & b[190])^(a[160] & b[191])^(a[159] & b[192])^(a[158] & b[193])^(a[157] & b[194])^(a[156] & b[195])^(a[155] & b[196])^(a[154] & b[197])^(a[153] & b[198])^(a[152] & b[199])^(a[151] & b[200])^(a[150] & b[201])^(a[149] & b[202])^(a[148] & b[203])^(a[147] & b[204])^(a[146] & b[205])^(a[145] & b[206])^(a[144] & b[207])^(a[143] & b[208])^(a[142] & b[209])^(a[141] & b[210])^(a[140] & b[211])^(a[139] & b[212])^(a[138] & b[213])^(a[137] & b[214])^(a[136] & b[215])^(a[135] & b[216])^(a[134] & b[217])^(a[133] & b[218])^(a[132] & b[219])^(a[131] & b[220])^(a[130] & b[221])^(a[129] & b[222])^(a[128] & b[223])^(a[127] & b[224])^(a[126] & b[225])^(a[125] & b[226])^(a[124] & b[227])^(a[123] & b[228])^(a[122] & b[229])^(a[121] & b[230])^(a[120] & b[231])^(a[119] & b[232]);
assign y[352] = (a[232] & b[120])^(a[231] & b[121])^(a[230] & b[122])^(a[229] & b[123])^(a[228] & b[124])^(a[227] & b[125])^(a[226] & b[126])^(a[225] & b[127])^(a[224] & b[128])^(a[223] & b[129])^(a[222] & b[130])^(a[221] & b[131])^(a[220] & b[132])^(a[219] & b[133])^(a[218] & b[134])^(a[217] & b[135])^(a[216] & b[136])^(a[215] & b[137])^(a[214] & b[138])^(a[213] & b[139])^(a[212] & b[140])^(a[211] & b[141])^(a[210] & b[142])^(a[209] & b[143])^(a[208] & b[144])^(a[207] & b[145])^(a[206] & b[146])^(a[205] & b[147])^(a[204] & b[148])^(a[203] & b[149])^(a[202] & b[150])^(a[201] & b[151])^(a[200] & b[152])^(a[199] & b[153])^(a[198] & b[154])^(a[197] & b[155])^(a[196] & b[156])^(a[195] & b[157])^(a[194] & b[158])^(a[193] & b[159])^(a[192] & b[160])^(a[191] & b[161])^(a[190] & b[162])^(a[189] & b[163])^(a[188] & b[164])^(a[187] & b[165])^(a[186] & b[166])^(a[185] & b[167])^(a[184] & b[168])^(a[183] & b[169])^(a[182] & b[170])^(a[181] & b[171])^(a[180] & b[172])^(a[179] & b[173])^(a[178] & b[174])^(a[177] & b[175])^(a[176] & b[176])^(a[175] & b[177])^(a[174] & b[178])^(a[173] & b[179])^(a[172] & b[180])^(a[171] & b[181])^(a[170] & b[182])^(a[169] & b[183])^(a[168] & b[184])^(a[167] & b[185])^(a[166] & b[186])^(a[165] & b[187])^(a[164] & b[188])^(a[163] & b[189])^(a[162] & b[190])^(a[161] & b[191])^(a[160] & b[192])^(a[159] & b[193])^(a[158] & b[194])^(a[157] & b[195])^(a[156] & b[196])^(a[155] & b[197])^(a[154] & b[198])^(a[153] & b[199])^(a[152] & b[200])^(a[151] & b[201])^(a[150] & b[202])^(a[149] & b[203])^(a[148] & b[204])^(a[147] & b[205])^(a[146] & b[206])^(a[145] & b[207])^(a[144] & b[208])^(a[143] & b[209])^(a[142] & b[210])^(a[141] & b[211])^(a[140] & b[212])^(a[139] & b[213])^(a[138] & b[214])^(a[137] & b[215])^(a[136] & b[216])^(a[135] & b[217])^(a[134] & b[218])^(a[133] & b[219])^(a[132] & b[220])^(a[131] & b[221])^(a[130] & b[222])^(a[129] & b[223])^(a[128] & b[224])^(a[127] & b[225])^(a[126] & b[226])^(a[125] & b[227])^(a[124] & b[228])^(a[123] & b[229])^(a[122] & b[230])^(a[121] & b[231])^(a[120] & b[232]);
assign y[353] = (a[232] & b[121])^(a[231] & b[122])^(a[230] & b[123])^(a[229] & b[124])^(a[228] & b[125])^(a[227] & b[126])^(a[226] & b[127])^(a[225] & b[128])^(a[224] & b[129])^(a[223] & b[130])^(a[222] & b[131])^(a[221] & b[132])^(a[220] & b[133])^(a[219] & b[134])^(a[218] & b[135])^(a[217] & b[136])^(a[216] & b[137])^(a[215] & b[138])^(a[214] & b[139])^(a[213] & b[140])^(a[212] & b[141])^(a[211] & b[142])^(a[210] & b[143])^(a[209] & b[144])^(a[208] & b[145])^(a[207] & b[146])^(a[206] & b[147])^(a[205] & b[148])^(a[204] & b[149])^(a[203] & b[150])^(a[202] & b[151])^(a[201] & b[152])^(a[200] & b[153])^(a[199] & b[154])^(a[198] & b[155])^(a[197] & b[156])^(a[196] & b[157])^(a[195] & b[158])^(a[194] & b[159])^(a[193] & b[160])^(a[192] & b[161])^(a[191] & b[162])^(a[190] & b[163])^(a[189] & b[164])^(a[188] & b[165])^(a[187] & b[166])^(a[186] & b[167])^(a[185] & b[168])^(a[184] & b[169])^(a[183] & b[170])^(a[182] & b[171])^(a[181] & b[172])^(a[180] & b[173])^(a[179] & b[174])^(a[178] & b[175])^(a[177] & b[176])^(a[176] & b[177])^(a[175] & b[178])^(a[174] & b[179])^(a[173] & b[180])^(a[172] & b[181])^(a[171] & b[182])^(a[170] & b[183])^(a[169] & b[184])^(a[168] & b[185])^(a[167] & b[186])^(a[166] & b[187])^(a[165] & b[188])^(a[164] & b[189])^(a[163] & b[190])^(a[162] & b[191])^(a[161] & b[192])^(a[160] & b[193])^(a[159] & b[194])^(a[158] & b[195])^(a[157] & b[196])^(a[156] & b[197])^(a[155] & b[198])^(a[154] & b[199])^(a[153] & b[200])^(a[152] & b[201])^(a[151] & b[202])^(a[150] & b[203])^(a[149] & b[204])^(a[148] & b[205])^(a[147] & b[206])^(a[146] & b[207])^(a[145] & b[208])^(a[144] & b[209])^(a[143] & b[210])^(a[142] & b[211])^(a[141] & b[212])^(a[140] & b[213])^(a[139] & b[214])^(a[138] & b[215])^(a[137] & b[216])^(a[136] & b[217])^(a[135] & b[218])^(a[134] & b[219])^(a[133] & b[220])^(a[132] & b[221])^(a[131] & b[222])^(a[130] & b[223])^(a[129] & b[224])^(a[128] & b[225])^(a[127] & b[226])^(a[126] & b[227])^(a[125] & b[228])^(a[124] & b[229])^(a[123] & b[230])^(a[122] & b[231])^(a[121] & b[232]);
assign y[354] = (a[232] & b[122])^(a[231] & b[123])^(a[230] & b[124])^(a[229] & b[125])^(a[228] & b[126])^(a[227] & b[127])^(a[226] & b[128])^(a[225] & b[129])^(a[224] & b[130])^(a[223] & b[131])^(a[222] & b[132])^(a[221] & b[133])^(a[220] & b[134])^(a[219] & b[135])^(a[218] & b[136])^(a[217] & b[137])^(a[216] & b[138])^(a[215] & b[139])^(a[214] & b[140])^(a[213] & b[141])^(a[212] & b[142])^(a[211] & b[143])^(a[210] & b[144])^(a[209] & b[145])^(a[208] & b[146])^(a[207] & b[147])^(a[206] & b[148])^(a[205] & b[149])^(a[204] & b[150])^(a[203] & b[151])^(a[202] & b[152])^(a[201] & b[153])^(a[200] & b[154])^(a[199] & b[155])^(a[198] & b[156])^(a[197] & b[157])^(a[196] & b[158])^(a[195] & b[159])^(a[194] & b[160])^(a[193] & b[161])^(a[192] & b[162])^(a[191] & b[163])^(a[190] & b[164])^(a[189] & b[165])^(a[188] & b[166])^(a[187] & b[167])^(a[186] & b[168])^(a[185] & b[169])^(a[184] & b[170])^(a[183] & b[171])^(a[182] & b[172])^(a[181] & b[173])^(a[180] & b[174])^(a[179] & b[175])^(a[178] & b[176])^(a[177] & b[177])^(a[176] & b[178])^(a[175] & b[179])^(a[174] & b[180])^(a[173] & b[181])^(a[172] & b[182])^(a[171] & b[183])^(a[170] & b[184])^(a[169] & b[185])^(a[168] & b[186])^(a[167] & b[187])^(a[166] & b[188])^(a[165] & b[189])^(a[164] & b[190])^(a[163] & b[191])^(a[162] & b[192])^(a[161] & b[193])^(a[160] & b[194])^(a[159] & b[195])^(a[158] & b[196])^(a[157] & b[197])^(a[156] & b[198])^(a[155] & b[199])^(a[154] & b[200])^(a[153] & b[201])^(a[152] & b[202])^(a[151] & b[203])^(a[150] & b[204])^(a[149] & b[205])^(a[148] & b[206])^(a[147] & b[207])^(a[146] & b[208])^(a[145] & b[209])^(a[144] & b[210])^(a[143] & b[211])^(a[142] & b[212])^(a[141] & b[213])^(a[140] & b[214])^(a[139] & b[215])^(a[138] & b[216])^(a[137] & b[217])^(a[136] & b[218])^(a[135] & b[219])^(a[134] & b[220])^(a[133] & b[221])^(a[132] & b[222])^(a[131] & b[223])^(a[130] & b[224])^(a[129] & b[225])^(a[128] & b[226])^(a[127] & b[227])^(a[126] & b[228])^(a[125] & b[229])^(a[124] & b[230])^(a[123] & b[231])^(a[122] & b[232]);
assign y[355] = (a[232] & b[123])^(a[231] & b[124])^(a[230] & b[125])^(a[229] & b[126])^(a[228] & b[127])^(a[227] & b[128])^(a[226] & b[129])^(a[225] & b[130])^(a[224] & b[131])^(a[223] & b[132])^(a[222] & b[133])^(a[221] & b[134])^(a[220] & b[135])^(a[219] & b[136])^(a[218] & b[137])^(a[217] & b[138])^(a[216] & b[139])^(a[215] & b[140])^(a[214] & b[141])^(a[213] & b[142])^(a[212] & b[143])^(a[211] & b[144])^(a[210] & b[145])^(a[209] & b[146])^(a[208] & b[147])^(a[207] & b[148])^(a[206] & b[149])^(a[205] & b[150])^(a[204] & b[151])^(a[203] & b[152])^(a[202] & b[153])^(a[201] & b[154])^(a[200] & b[155])^(a[199] & b[156])^(a[198] & b[157])^(a[197] & b[158])^(a[196] & b[159])^(a[195] & b[160])^(a[194] & b[161])^(a[193] & b[162])^(a[192] & b[163])^(a[191] & b[164])^(a[190] & b[165])^(a[189] & b[166])^(a[188] & b[167])^(a[187] & b[168])^(a[186] & b[169])^(a[185] & b[170])^(a[184] & b[171])^(a[183] & b[172])^(a[182] & b[173])^(a[181] & b[174])^(a[180] & b[175])^(a[179] & b[176])^(a[178] & b[177])^(a[177] & b[178])^(a[176] & b[179])^(a[175] & b[180])^(a[174] & b[181])^(a[173] & b[182])^(a[172] & b[183])^(a[171] & b[184])^(a[170] & b[185])^(a[169] & b[186])^(a[168] & b[187])^(a[167] & b[188])^(a[166] & b[189])^(a[165] & b[190])^(a[164] & b[191])^(a[163] & b[192])^(a[162] & b[193])^(a[161] & b[194])^(a[160] & b[195])^(a[159] & b[196])^(a[158] & b[197])^(a[157] & b[198])^(a[156] & b[199])^(a[155] & b[200])^(a[154] & b[201])^(a[153] & b[202])^(a[152] & b[203])^(a[151] & b[204])^(a[150] & b[205])^(a[149] & b[206])^(a[148] & b[207])^(a[147] & b[208])^(a[146] & b[209])^(a[145] & b[210])^(a[144] & b[211])^(a[143] & b[212])^(a[142] & b[213])^(a[141] & b[214])^(a[140] & b[215])^(a[139] & b[216])^(a[138] & b[217])^(a[137] & b[218])^(a[136] & b[219])^(a[135] & b[220])^(a[134] & b[221])^(a[133] & b[222])^(a[132] & b[223])^(a[131] & b[224])^(a[130] & b[225])^(a[129] & b[226])^(a[128] & b[227])^(a[127] & b[228])^(a[126] & b[229])^(a[125] & b[230])^(a[124] & b[231])^(a[123] & b[232]);
assign y[356] = (a[232] & b[124])^(a[231] & b[125])^(a[230] & b[126])^(a[229] & b[127])^(a[228] & b[128])^(a[227] & b[129])^(a[226] & b[130])^(a[225] & b[131])^(a[224] & b[132])^(a[223] & b[133])^(a[222] & b[134])^(a[221] & b[135])^(a[220] & b[136])^(a[219] & b[137])^(a[218] & b[138])^(a[217] & b[139])^(a[216] & b[140])^(a[215] & b[141])^(a[214] & b[142])^(a[213] & b[143])^(a[212] & b[144])^(a[211] & b[145])^(a[210] & b[146])^(a[209] & b[147])^(a[208] & b[148])^(a[207] & b[149])^(a[206] & b[150])^(a[205] & b[151])^(a[204] & b[152])^(a[203] & b[153])^(a[202] & b[154])^(a[201] & b[155])^(a[200] & b[156])^(a[199] & b[157])^(a[198] & b[158])^(a[197] & b[159])^(a[196] & b[160])^(a[195] & b[161])^(a[194] & b[162])^(a[193] & b[163])^(a[192] & b[164])^(a[191] & b[165])^(a[190] & b[166])^(a[189] & b[167])^(a[188] & b[168])^(a[187] & b[169])^(a[186] & b[170])^(a[185] & b[171])^(a[184] & b[172])^(a[183] & b[173])^(a[182] & b[174])^(a[181] & b[175])^(a[180] & b[176])^(a[179] & b[177])^(a[178] & b[178])^(a[177] & b[179])^(a[176] & b[180])^(a[175] & b[181])^(a[174] & b[182])^(a[173] & b[183])^(a[172] & b[184])^(a[171] & b[185])^(a[170] & b[186])^(a[169] & b[187])^(a[168] & b[188])^(a[167] & b[189])^(a[166] & b[190])^(a[165] & b[191])^(a[164] & b[192])^(a[163] & b[193])^(a[162] & b[194])^(a[161] & b[195])^(a[160] & b[196])^(a[159] & b[197])^(a[158] & b[198])^(a[157] & b[199])^(a[156] & b[200])^(a[155] & b[201])^(a[154] & b[202])^(a[153] & b[203])^(a[152] & b[204])^(a[151] & b[205])^(a[150] & b[206])^(a[149] & b[207])^(a[148] & b[208])^(a[147] & b[209])^(a[146] & b[210])^(a[145] & b[211])^(a[144] & b[212])^(a[143] & b[213])^(a[142] & b[214])^(a[141] & b[215])^(a[140] & b[216])^(a[139] & b[217])^(a[138] & b[218])^(a[137] & b[219])^(a[136] & b[220])^(a[135] & b[221])^(a[134] & b[222])^(a[133] & b[223])^(a[132] & b[224])^(a[131] & b[225])^(a[130] & b[226])^(a[129] & b[227])^(a[128] & b[228])^(a[127] & b[229])^(a[126] & b[230])^(a[125] & b[231])^(a[124] & b[232]);
assign y[357] = (a[232] & b[125])^(a[231] & b[126])^(a[230] & b[127])^(a[229] & b[128])^(a[228] & b[129])^(a[227] & b[130])^(a[226] & b[131])^(a[225] & b[132])^(a[224] & b[133])^(a[223] & b[134])^(a[222] & b[135])^(a[221] & b[136])^(a[220] & b[137])^(a[219] & b[138])^(a[218] & b[139])^(a[217] & b[140])^(a[216] & b[141])^(a[215] & b[142])^(a[214] & b[143])^(a[213] & b[144])^(a[212] & b[145])^(a[211] & b[146])^(a[210] & b[147])^(a[209] & b[148])^(a[208] & b[149])^(a[207] & b[150])^(a[206] & b[151])^(a[205] & b[152])^(a[204] & b[153])^(a[203] & b[154])^(a[202] & b[155])^(a[201] & b[156])^(a[200] & b[157])^(a[199] & b[158])^(a[198] & b[159])^(a[197] & b[160])^(a[196] & b[161])^(a[195] & b[162])^(a[194] & b[163])^(a[193] & b[164])^(a[192] & b[165])^(a[191] & b[166])^(a[190] & b[167])^(a[189] & b[168])^(a[188] & b[169])^(a[187] & b[170])^(a[186] & b[171])^(a[185] & b[172])^(a[184] & b[173])^(a[183] & b[174])^(a[182] & b[175])^(a[181] & b[176])^(a[180] & b[177])^(a[179] & b[178])^(a[178] & b[179])^(a[177] & b[180])^(a[176] & b[181])^(a[175] & b[182])^(a[174] & b[183])^(a[173] & b[184])^(a[172] & b[185])^(a[171] & b[186])^(a[170] & b[187])^(a[169] & b[188])^(a[168] & b[189])^(a[167] & b[190])^(a[166] & b[191])^(a[165] & b[192])^(a[164] & b[193])^(a[163] & b[194])^(a[162] & b[195])^(a[161] & b[196])^(a[160] & b[197])^(a[159] & b[198])^(a[158] & b[199])^(a[157] & b[200])^(a[156] & b[201])^(a[155] & b[202])^(a[154] & b[203])^(a[153] & b[204])^(a[152] & b[205])^(a[151] & b[206])^(a[150] & b[207])^(a[149] & b[208])^(a[148] & b[209])^(a[147] & b[210])^(a[146] & b[211])^(a[145] & b[212])^(a[144] & b[213])^(a[143] & b[214])^(a[142] & b[215])^(a[141] & b[216])^(a[140] & b[217])^(a[139] & b[218])^(a[138] & b[219])^(a[137] & b[220])^(a[136] & b[221])^(a[135] & b[222])^(a[134] & b[223])^(a[133] & b[224])^(a[132] & b[225])^(a[131] & b[226])^(a[130] & b[227])^(a[129] & b[228])^(a[128] & b[229])^(a[127] & b[230])^(a[126] & b[231])^(a[125] & b[232]);
assign y[358] = (a[232] & b[126])^(a[231] & b[127])^(a[230] & b[128])^(a[229] & b[129])^(a[228] & b[130])^(a[227] & b[131])^(a[226] & b[132])^(a[225] & b[133])^(a[224] & b[134])^(a[223] & b[135])^(a[222] & b[136])^(a[221] & b[137])^(a[220] & b[138])^(a[219] & b[139])^(a[218] & b[140])^(a[217] & b[141])^(a[216] & b[142])^(a[215] & b[143])^(a[214] & b[144])^(a[213] & b[145])^(a[212] & b[146])^(a[211] & b[147])^(a[210] & b[148])^(a[209] & b[149])^(a[208] & b[150])^(a[207] & b[151])^(a[206] & b[152])^(a[205] & b[153])^(a[204] & b[154])^(a[203] & b[155])^(a[202] & b[156])^(a[201] & b[157])^(a[200] & b[158])^(a[199] & b[159])^(a[198] & b[160])^(a[197] & b[161])^(a[196] & b[162])^(a[195] & b[163])^(a[194] & b[164])^(a[193] & b[165])^(a[192] & b[166])^(a[191] & b[167])^(a[190] & b[168])^(a[189] & b[169])^(a[188] & b[170])^(a[187] & b[171])^(a[186] & b[172])^(a[185] & b[173])^(a[184] & b[174])^(a[183] & b[175])^(a[182] & b[176])^(a[181] & b[177])^(a[180] & b[178])^(a[179] & b[179])^(a[178] & b[180])^(a[177] & b[181])^(a[176] & b[182])^(a[175] & b[183])^(a[174] & b[184])^(a[173] & b[185])^(a[172] & b[186])^(a[171] & b[187])^(a[170] & b[188])^(a[169] & b[189])^(a[168] & b[190])^(a[167] & b[191])^(a[166] & b[192])^(a[165] & b[193])^(a[164] & b[194])^(a[163] & b[195])^(a[162] & b[196])^(a[161] & b[197])^(a[160] & b[198])^(a[159] & b[199])^(a[158] & b[200])^(a[157] & b[201])^(a[156] & b[202])^(a[155] & b[203])^(a[154] & b[204])^(a[153] & b[205])^(a[152] & b[206])^(a[151] & b[207])^(a[150] & b[208])^(a[149] & b[209])^(a[148] & b[210])^(a[147] & b[211])^(a[146] & b[212])^(a[145] & b[213])^(a[144] & b[214])^(a[143] & b[215])^(a[142] & b[216])^(a[141] & b[217])^(a[140] & b[218])^(a[139] & b[219])^(a[138] & b[220])^(a[137] & b[221])^(a[136] & b[222])^(a[135] & b[223])^(a[134] & b[224])^(a[133] & b[225])^(a[132] & b[226])^(a[131] & b[227])^(a[130] & b[228])^(a[129] & b[229])^(a[128] & b[230])^(a[127] & b[231])^(a[126] & b[232]);
assign y[359] = (a[232] & b[127])^(a[231] & b[128])^(a[230] & b[129])^(a[229] & b[130])^(a[228] & b[131])^(a[227] & b[132])^(a[226] & b[133])^(a[225] & b[134])^(a[224] & b[135])^(a[223] & b[136])^(a[222] & b[137])^(a[221] & b[138])^(a[220] & b[139])^(a[219] & b[140])^(a[218] & b[141])^(a[217] & b[142])^(a[216] & b[143])^(a[215] & b[144])^(a[214] & b[145])^(a[213] & b[146])^(a[212] & b[147])^(a[211] & b[148])^(a[210] & b[149])^(a[209] & b[150])^(a[208] & b[151])^(a[207] & b[152])^(a[206] & b[153])^(a[205] & b[154])^(a[204] & b[155])^(a[203] & b[156])^(a[202] & b[157])^(a[201] & b[158])^(a[200] & b[159])^(a[199] & b[160])^(a[198] & b[161])^(a[197] & b[162])^(a[196] & b[163])^(a[195] & b[164])^(a[194] & b[165])^(a[193] & b[166])^(a[192] & b[167])^(a[191] & b[168])^(a[190] & b[169])^(a[189] & b[170])^(a[188] & b[171])^(a[187] & b[172])^(a[186] & b[173])^(a[185] & b[174])^(a[184] & b[175])^(a[183] & b[176])^(a[182] & b[177])^(a[181] & b[178])^(a[180] & b[179])^(a[179] & b[180])^(a[178] & b[181])^(a[177] & b[182])^(a[176] & b[183])^(a[175] & b[184])^(a[174] & b[185])^(a[173] & b[186])^(a[172] & b[187])^(a[171] & b[188])^(a[170] & b[189])^(a[169] & b[190])^(a[168] & b[191])^(a[167] & b[192])^(a[166] & b[193])^(a[165] & b[194])^(a[164] & b[195])^(a[163] & b[196])^(a[162] & b[197])^(a[161] & b[198])^(a[160] & b[199])^(a[159] & b[200])^(a[158] & b[201])^(a[157] & b[202])^(a[156] & b[203])^(a[155] & b[204])^(a[154] & b[205])^(a[153] & b[206])^(a[152] & b[207])^(a[151] & b[208])^(a[150] & b[209])^(a[149] & b[210])^(a[148] & b[211])^(a[147] & b[212])^(a[146] & b[213])^(a[145] & b[214])^(a[144] & b[215])^(a[143] & b[216])^(a[142] & b[217])^(a[141] & b[218])^(a[140] & b[219])^(a[139] & b[220])^(a[138] & b[221])^(a[137] & b[222])^(a[136] & b[223])^(a[135] & b[224])^(a[134] & b[225])^(a[133] & b[226])^(a[132] & b[227])^(a[131] & b[228])^(a[130] & b[229])^(a[129] & b[230])^(a[128] & b[231])^(a[127] & b[232]);
assign y[360] = (a[232] & b[128])^(a[231] & b[129])^(a[230] & b[130])^(a[229] & b[131])^(a[228] & b[132])^(a[227] & b[133])^(a[226] & b[134])^(a[225] & b[135])^(a[224] & b[136])^(a[223] & b[137])^(a[222] & b[138])^(a[221] & b[139])^(a[220] & b[140])^(a[219] & b[141])^(a[218] & b[142])^(a[217] & b[143])^(a[216] & b[144])^(a[215] & b[145])^(a[214] & b[146])^(a[213] & b[147])^(a[212] & b[148])^(a[211] & b[149])^(a[210] & b[150])^(a[209] & b[151])^(a[208] & b[152])^(a[207] & b[153])^(a[206] & b[154])^(a[205] & b[155])^(a[204] & b[156])^(a[203] & b[157])^(a[202] & b[158])^(a[201] & b[159])^(a[200] & b[160])^(a[199] & b[161])^(a[198] & b[162])^(a[197] & b[163])^(a[196] & b[164])^(a[195] & b[165])^(a[194] & b[166])^(a[193] & b[167])^(a[192] & b[168])^(a[191] & b[169])^(a[190] & b[170])^(a[189] & b[171])^(a[188] & b[172])^(a[187] & b[173])^(a[186] & b[174])^(a[185] & b[175])^(a[184] & b[176])^(a[183] & b[177])^(a[182] & b[178])^(a[181] & b[179])^(a[180] & b[180])^(a[179] & b[181])^(a[178] & b[182])^(a[177] & b[183])^(a[176] & b[184])^(a[175] & b[185])^(a[174] & b[186])^(a[173] & b[187])^(a[172] & b[188])^(a[171] & b[189])^(a[170] & b[190])^(a[169] & b[191])^(a[168] & b[192])^(a[167] & b[193])^(a[166] & b[194])^(a[165] & b[195])^(a[164] & b[196])^(a[163] & b[197])^(a[162] & b[198])^(a[161] & b[199])^(a[160] & b[200])^(a[159] & b[201])^(a[158] & b[202])^(a[157] & b[203])^(a[156] & b[204])^(a[155] & b[205])^(a[154] & b[206])^(a[153] & b[207])^(a[152] & b[208])^(a[151] & b[209])^(a[150] & b[210])^(a[149] & b[211])^(a[148] & b[212])^(a[147] & b[213])^(a[146] & b[214])^(a[145] & b[215])^(a[144] & b[216])^(a[143] & b[217])^(a[142] & b[218])^(a[141] & b[219])^(a[140] & b[220])^(a[139] & b[221])^(a[138] & b[222])^(a[137] & b[223])^(a[136] & b[224])^(a[135] & b[225])^(a[134] & b[226])^(a[133] & b[227])^(a[132] & b[228])^(a[131] & b[229])^(a[130] & b[230])^(a[129] & b[231])^(a[128] & b[232]);
assign y[361] = (a[232] & b[129])^(a[231] & b[130])^(a[230] & b[131])^(a[229] & b[132])^(a[228] & b[133])^(a[227] & b[134])^(a[226] & b[135])^(a[225] & b[136])^(a[224] & b[137])^(a[223] & b[138])^(a[222] & b[139])^(a[221] & b[140])^(a[220] & b[141])^(a[219] & b[142])^(a[218] & b[143])^(a[217] & b[144])^(a[216] & b[145])^(a[215] & b[146])^(a[214] & b[147])^(a[213] & b[148])^(a[212] & b[149])^(a[211] & b[150])^(a[210] & b[151])^(a[209] & b[152])^(a[208] & b[153])^(a[207] & b[154])^(a[206] & b[155])^(a[205] & b[156])^(a[204] & b[157])^(a[203] & b[158])^(a[202] & b[159])^(a[201] & b[160])^(a[200] & b[161])^(a[199] & b[162])^(a[198] & b[163])^(a[197] & b[164])^(a[196] & b[165])^(a[195] & b[166])^(a[194] & b[167])^(a[193] & b[168])^(a[192] & b[169])^(a[191] & b[170])^(a[190] & b[171])^(a[189] & b[172])^(a[188] & b[173])^(a[187] & b[174])^(a[186] & b[175])^(a[185] & b[176])^(a[184] & b[177])^(a[183] & b[178])^(a[182] & b[179])^(a[181] & b[180])^(a[180] & b[181])^(a[179] & b[182])^(a[178] & b[183])^(a[177] & b[184])^(a[176] & b[185])^(a[175] & b[186])^(a[174] & b[187])^(a[173] & b[188])^(a[172] & b[189])^(a[171] & b[190])^(a[170] & b[191])^(a[169] & b[192])^(a[168] & b[193])^(a[167] & b[194])^(a[166] & b[195])^(a[165] & b[196])^(a[164] & b[197])^(a[163] & b[198])^(a[162] & b[199])^(a[161] & b[200])^(a[160] & b[201])^(a[159] & b[202])^(a[158] & b[203])^(a[157] & b[204])^(a[156] & b[205])^(a[155] & b[206])^(a[154] & b[207])^(a[153] & b[208])^(a[152] & b[209])^(a[151] & b[210])^(a[150] & b[211])^(a[149] & b[212])^(a[148] & b[213])^(a[147] & b[214])^(a[146] & b[215])^(a[145] & b[216])^(a[144] & b[217])^(a[143] & b[218])^(a[142] & b[219])^(a[141] & b[220])^(a[140] & b[221])^(a[139] & b[222])^(a[138] & b[223])^(a[137] & b[224])^(a[136] & b[225])^(a[135] & b[226])^(a[134] & b[227])^(a[133] & b[228])^(a[132] & b[229])^(a[131] & b[230])^(a[130] & b[231])^(a[129] & b[232]);
assign y[362] = (a[232] & b[130])^(a[231] & b[131])^(a[230] & b[132])^(a[229] & b[133])^(a[228] & b[134])^(a[227] & b[135])^(a[226] & b[136])^(a[225] & b[137])^(a[224] & b[138])^(a[223] & b[139])^(a[222] & b[140])^(a[221] & b[141])^(a[220] & b[142])^(a[219] & b[143])^(a[218] & b[144])^(a[217] & b[145])^(a[216] & b[146])^(a[215] & b[147])^(a[214] & b[148])^(a[213] & b[149])^(a[212] & b[150])^(a[211] & b[151])^(a[210] & b[152])^(a[209] & b[153])^(a[208] & b[154])^(a[207] & b[155])^(a[206] & b[156])^(a[205] & b[157])^(a[204] & b[158])^(a[203] & b[159])^(a[202] & b[160])^(a[201] & b[161])^(a[200] & b[162])^(a[199] & b[163])^(a[198] & b[164])^(a[197] & b[165])^(a[196] & b[166])^(a[195] & b[167])^(a[194] & b[168])^(a[193] & b[169])^(a[192] & b[170])^(a[191] & b[171])^(a[190] & b[172])^(a[189] & b[173])^(a[188] & b[174])^(a[187] & b[175])^(a[186] & b[176])^(a[185] & b[177])^(a[184] & b[178])^(a[183] & b[179])^(a[182] & b[180])^(a[181] & b[181])^(a[180] & b[182])^(a[179] & b[183])^(a[178] & b[184])^(a[177] & b[185])^(a[176] & b[186])^(a[175] & b[187])^(a[174] & b[188])^(a[173] & b[189])^(a[172] & b[190])^(a[171] & b[191])^(a[170] & b[192])^(a[169] & b[193])^(a[168] & b[194])^(a[167] & b[195])^(a[166] & b[196])^(a[165] & b[197])^(a[164] & b[198])^(a[163] & b[199])^(a[162] & b[200])^(a[161] & b[201])^(a[160] & b[202])^(a[159] & b[203])^(a[158] & b[204])^(a[157] & b[205])^(a[156] & b[206])^(a[155] & b[207])^(a[154] & b[208])^(a[153] & b[209])^(a[152] & b[210])^(a[151] & b[211])^(a[150] & b[212])^(a[149] & b[213])^(a[148] & b[214])^(a[147] & b[215])^(a[146] & b[216])^(a[145] & b[217])^(a[144] & b[218])^(a[143] & b[219])^(a[142] & b[220])^(a[141] & b[221])^(a[140] & b[222])^(a[139] & b[223])^(a[138] & b[224])^(a[137] & b[225])^(a[136] & b[226])^(a[135] & b[227])^(a[134] & b[228])^(a[133] & b[229])^(a[132] & b[230])^(a[131] & b[231])^(a[130] & b[232]);
assign y[363] = (a[232] & b[131])^(a[231] & b[132])^(a[230] & b[133])^(a[229] & b[134])^(a[228] & b[135])^(a[227] & b[136])^(a[226] & b[137])^(a[225] & b[138])^(a[224] & b[139])^(a[223] & b[140])^(a[222] & b[141])^(a[221] & b[142])^(a[220] & b[143])^(a[219] & b[144])^(a[218] & b[145])^(a[217] & b[146])^(a[216] & b[147])^(a[215] & b[148])^(a[214] & b[149])^(a[213] & b[150])^(a[212] & b[151])^(a[211] & b[152])^(a[210] & b[153])^(a[209] & b[154])^(a[208] & b[155])^(a[207] & b[156])^(a[206] & b[157])^(a[205] & b[158])^(a[204] & b[159])^(a[203] & b[160])^(a[202] & b[161])^(a[201] & b[162])^(a[200] & b[163])^(a[199] & b[164])^(a[198] & b[165])^(a[197] & b[166])^(a[196] & b[167])^(a[195] & b[168])^(a[194] & b[169])^(a[193] & b[170])^(a[192] & b[171])^(a[191] & b[172])^(a[190] & b[173])^(a[189] & b[174])^(a[188] & b[175])^(a[187] & b[176])^(a[186] & b[177])^(a[185] & b[178])^(a[184] & b[179])^(a[183] & b[180])^(a[182] & b[181])^(a[181] & b[182])^(a[180] & b[183])^(a[179] & b[184])^(a[178] & b[185])^(a[177] & b[186])^(a[176] & b[187])^(a[175] & b[188])^(a[174] & b[189])^(a[173] & b[190])^(a[172] & b[191])^(a[171] & b[192])^(a[170] & b[193])^(a[169] & b[194])^(a[168] & b[195])^(a[167] & b[196])^(a[166] & b[197])^(a[165] & b[198])^(a[164] & b[199])^(a[163] & b[200])^(a[162] & b[201])^(a[161] & b[202])^(a[160] & b[203])^(a[159] & b[204])^(a[158] & b[205])^(a[157] & b[206])^(a[156] & b[207])^(a[155] & b[208])^(a[154] & b[209])^(a[153] & b[210])^(a[152] & b[211])^(a[151] & b[212])^(a[150] & b[213])^(a[149] & b[214])^(a[148] & b[215])^(a[147] & b[216])^(a[146] & b[217])^(a[145] & b[218])^(a[144] & b[219])^(a[143] & b[220])^(a[142] & b[221])^(a[141] & b[222])^(a[140] & b[223])^(a[139] & b[224])^(a[138] & b[225])^(a[137] & b[226])^(a[136] & b[227])^(a[135] & b[228])^(a[134] & b[229])^(a[133] & b[230])^(a[132] & b[231])^(a[131] & b[232]);
assign y[364] = (a[232] & b[132])^(a[231] & b[133])^(a[230] & b[134])^(a[229] & b[135])^(a[228] & b[136])^(a[227] & b[137])^(a[226] & b[138])^(a[225] & b[139])^(a[224] & b[140])^(a[223] & b[141])^(a[222] & b[142])^(a[221] & b[143])^(a[220] & b[144])^(a[219] & b[145])^(a[218] & b[146])^(a[217] & b[147])^(a[216] & b[148])^(a[215] & b[149])^(a[214] & b[150])^(a[213] & b[151])^(a[212] & b[152])^(a[211] & b[153])^(a[210] & b[154])^(a[209] & b[155])^(a[208] & b[156])^(a[207] & b[157])^(a[206] & b[158])^(a[205] & b[159])^(a[204] & b[160])^(a[203] & b[161])^(a[202] & b[162])^(a[201] & b[163])^(a[200] & b[164])^(a[199] & b[165])^(a[198] & b[166])^(a[197] & b[167])^(a[196] & b[168])^(a[195] & b[169])^(a[194] & b[170])^(a[193] & b[171])^(a[192] & b[172])^(a[191] & b[173])^(a[190] & b[174])^(a[189] & b[175])^(a[188] & b[176])^(a[187] & b[177])^(a[186] & b[178])^(a[185] & b[179])^(a[184] & b[180])^(a[183] & b[181])^(a[182] & b[182])^(a[181] & b[183])^(a[180] & b[184])^(a[179] & b[185])^(a[178] & b[186])^(a[177] & b[187])^(a[176] & b[188])^(a[175] & b[189])^(a[174] & b[190])^(a[173] & b[191])^(a[172] & b[192])^(a[171] & b[193])^(a[170] & b[194])^(a[169] & b[195])^(a[168] & b[196])^(a[167] & b[197])^(a[166] & b[198])^(a[165] & b[199])^(a[164] & b[200])^(a[163] & b[201])^(a[162] & b[202])^(a[161] & b[203])^(a[160] & b[204])^(a[159] & b[205])^(a[158] & b[206])^(a[157] & b[207])^(a[156] & b[208])^(a[155] & b[209])^(a[154] & b[210])^(a[153] & b[211])^(a[152] & b[212])^(a[151] & b[213])^(a[150] & b[214])^(a[149] & b[215])^(a[148] & b[216])^(a[147] & b[217])^(a[146] & b[218])^(a[145] & b[219])^(a[144] & b[220])^(a[143] & b[221])^(a[142] & b[222])^(a[141] & b[223])^(a[140] & b[224])^(a[139] & b[225])^(a[138] & b[226])^(a[137] & b[227])^(a[136] & b[228])^(a[135] & b[229])^(a[134] & b[230])^(a[133] & b[231])^(a[132] & b[232]);
assign y[365] = (a[232] & b[133])^(a[231] & b[134])^(a[230] & b[135])^(a[229] & b[136])^(a[228] & b[137])^(a[227] & b[138])^(a[226] & b[139])^(a[225] & b[140])^(a[224] & b[141])^(a[223] & b[142])^(a[222] & b[143])^(a[221] & b[144])^(a[220] & b[145])^(a[219] & b[146])^(a[218] & b[147])^(a[217] & b[148])^(a[216] & b[149])^(a[215] & b[150])^(a[214] & b[151])^(a[213] & b[152])^(a[212] & b[153])^(a[211] & b[154])^(a[210] & b[155])^(a[209] & b[156])^(a[208] & b[157])^(a[207] & b[158])^(a[206] & b[159])^(a[205] & b[160])^(a[204] & b[161])^(a[203] & b[162])^(a[202] & b[163])^(a[201] & b[164])^(a[200] & b[165])^(a[199] & b[166])^(a[198] & b[167])^(a[197] & b[168])^(a[196] & b[169])^(a[195] & b[170])^(a[194] & b[171])^(a[193] & b[172])^(a[192] & b[173])^(a[191] & b[174])^(a[190] & b[175])^(a[189] & b[176])^(a[188] & b[177])^(a[187] & b[178])^(a[186] & b[179])^(a[185] & b[180])^(a[184] & b[181])^(a[183] & b[182])^(a[182] & b[183])^(a[181] & b[184])^(a[180] & b[185])^(a[179] & b[186])^(a[178] & b[187])^(a[177] & b[188])^(a[176] & b[189])^(a[175] & b[190])^(a[174] & b[191])^(a[173] & b[192])^(a[172] & b[193])^(a[171] & b[194])^(a[170] & b[195])^(a[169] & b[196])^(a[168] & b[197])^(a[167] & b[198])^(a[166] & b[199])^(a[165] & b[200])^(a[164] & b[201])^(a[163] & b[202])^(a[162] & b[203])^(a[161] & b[204])^(a[160] & b[205])^(a[159] & b[206])^(a[158] & b[207])^(a[157] & b[208])^(a[156] & b[209])^(a[155] & b[210])^(a[154] & b[211])^(a[153] & b[212])^(a[152] & b[213])^(a[151] & b[214])^(a[150] & b[215])^(a[149] & b[216])^(a[148] & b[217])^(a[147] & b[218])^(a[146] & b[219])^(a[145] & b[220])^(a[144] & b[221])^(a[143] & b[222])^(a[142] & b[223])^(a[141] & b[224])^(a[140] & b[225])^(a[139] & b[226])^(a[138] & b[227])^(a[137] & b[228])^(a[136] & b[229])^(a[135] & b[230])^(a[134] & b[231])^(a[133] & b[232]);
assign y[366] = (a[232] & b[134])^(a[231] & b[135])^(a[230] & b[136])^(a[229] & b[137])^(a[228] & b[138])^(a[227] & b[139])^(a[226] & b[140])^(a[225] & b[141])^(a[224] & b[142])^(a[223] & b[143])^(a[222] & b[144])^(a[221] & b[145])^(a[220] & b[146])^(a[219] & b[147])^(a[218] & b[148])^(a[217] & b[149])^(a[216] & b[150])^(a[215] & b[151])^(a[214] & b[152])^(a[213] & b[153])^(a[212] & b[154])^(a[211] & b[155])^(a[210] & b[156])^(a[209] & b[157])^(a[208] & b[158])^(a[207] & b[159])^(a[206] & b[160])^(a[205] & b[161])^(a[204] & b[162])^(a[203] & b[163])^(a[202] & b[164])^(a[201] & b[165])^(a[200] & b[166])^(a[199] & b[167])^(a[198] & b[168])^(a[197] & b[169])^(a[196] & b[170])^(a[195] & b[171])^(a[194] & b[172])^(a[193] & b[173])^(a[192] & b[174])^(a[191] & b[175])^(a[190] & b[176])^(a[189] & b[177])^(a[188] & b[178])^(a[187] & b[179])^(a[186] & b[180])^(a[185] & b[181])^(a[184] & b[182])^(a[183] & b[183])^(a[182] & b[184])^(a[181] & b[185])^(a[180] & b[186])^(a[179] & b[187])^(a[178] & b[188])^(a[177] & b[189])^(a[176] & b[190])^(a[175] & b[191])^(a[174] & b[192])^(a[173] & b[193])^(a[172] & b[194])^(a[171] & b[195])^(a[170] & b[196])^(a[169] & b[197])^(a[168] & b[198])^(a[167] & b[199])^(a[166] & b[200])^(a[165] & b[201])^(a[164] & b[202])^(a[163] & b[203])^(a[162] & b[204])^(a[161] & b[205])^(a[160] & b[206])^(a[159] & b[207])^(a[158] & b[208])^(a[157] & b[209])^(a[156] & b[210])^(a[155] & b[211])^(a[154] & b[212])^(a[153] & b[213])^(a[152] & b[214])^(a[151] & b[215])^(a[150] & b[216])^(a[149] & b[217])^(a[148] & b[218])^(a[147] & b[219])^(a[146] & b[220])^(a[145] & b[221])^(a[144] & b[222])^(a[143] & b[223])^(a[142] & b[224])^(a[141] & b[225])^(a[140] & b[226])^(a[139] & b[227])^(a[138] & b[228])^(a[137] & b[229])^(a[136] & b[230])^(a[135] & b[231])^(a[134] & b[232]);
assign y[367] = (a[232] & b[135])^(a[231] & b[136])^(a[230] & b[137])^(a[229] & b[138])^(a[228] & b[139])^(a[227] & b[140])^(a[226] & b[141])^(a[225] & b[142])^(a[224] & b[143])^(a[223] & b[144])^(a[222] & b[145])^(a[221] & b[146])^(a[220] & b[147])^(a[219] & b[148])^(a[218] & b[149])^(a[217] & b[150])^(a[216] & b[151])^(a[215] & b[152])^(a[214] & b[153])^(a[213] & b[154])^(a[212] & b[155])^(a[211] & b[156])^(a[210] & b[157])^(a[209] & b[158])^(a[208] & b[159])^(a[207] & b[160])^(a[206] & b[161])^(a[205] & b[162])^(a[204] & b[163])^(a[203] & b[164])^(a[202] & b[165])^(a[201] & b[166])^(a[200] & b[167])^(a[199] & b[168])^(a[198] & b[169])^(a[197] & b[170])^(a[196] & b[171])^(a[195] & b[172])^(a[194] & b[173])^(a[193] & b[174])^(a[192] & b[175])^(a[191] & b[176])^(a[190] & b[177])^(a[189] & b[178])^(a[188] & b[179])^(a[187] & b[180])^(a[186] & b[181])^(a[185] & b[182])^(a[184] & b[183])^(a[183] & b[184])^(a[182] & b[185])^(a[181] & b[186])^(a[180] & b[187])^(a[179] & b[188])^(a[178] & b[189])^(a[177] & b[190])^(a[176] & b[191])^(a[175] & b[192])^(a[174] & b[193])^(a[173] & b[194])^(a[172] & b[195])^(a[171] & b[196])^(a[170] & b[197])^(a[169] & b[198])^(a[168] & b[199])^(a[167] & b[200])^(a[166] & b[201])^(a[165] & b[202])^(a[164] & b[203])^(a[163] & b[204])^(a[162] & b[205])^(a[161] & b[206])^(a[160] & b[207])^(a[159] & b[208])^(a[158] & b[209])^(a[157] & b[210])^(a[156] & b[211])^(a[155] & b[212])^(a[154] & b[213])^(a[153] & b[214])^(a[152] & b[215])^(a[151] & b[216])^(a[150] & b[217])^(a[149] & b[218])^(a[148] & b[219])^(a[147] & b[220])^(a[146] & b[221])^(a[145] & b[222])^(a[144] & b[223])^(a[143] & b[224])^(a[142] & b[225])^(a[141] & b[226])^(a[140] & b[227])^(a[139] & b[228])^(a[138] & b[229])^(a[137] & b[230])^(a[136] & b[231])^(a[135] & b[232]);
assign y[368] = (a[232] & b[136])^(a[231] & b[137])^(a[230] & b[138])^(a[229] & b[139])^(a[228] & b[140])^(a[227] & b[141])^(a[226] & b[142])^(a[225] & b[143])^(a[224] & b[144])^(a[223] & b[145])^(a[222] & b[146])^(a[221] & b[147])^(a[220] & b[148])^(a[219] & b[149])^(a[218] & b[150])^(a[217] & b[151])^(a[216] & b[152])^(a[215] & b[153])^(a[214] & b[154])^(a[213] & b[155])^(a[212] & b[156])^(a[211] & b[157])^(a[210] & b[158])^(a[209] & b[159])^(a[208] & b[160])^(a[207] & b[161])^(a[206] & b[162])^(a[205] & b[163])^(a[204] & b[164])^(a[203] & b[165])^(a[202] & b[166])^(a[201] & b[167])^(a[200] & b[168])^(a[199] & b[169])^(a[198] & b[170])^(a[197] & b[171])^(a[196] & b[172])^(a[195] & b[173])^(a[194] & b[174])^(a[193] & b[175])^(a[192] & b[176])^(a[191] & b[177])^(a[190] & b[178])^(a[189] & b[179])^(a[188] & b[180])^(a[187] & b[181])^(a[186] & b[182])^(a[185] & b[183])^(a[184] & b[184])^(a[183] & b[185])^(a[182] & b[186])^(a[181] & b[187])^(a[180] & b[188])^(a[179] & b[189])^(a[178] & b[190])^(a[177] & b[191])^(a[176] & b[192])^(a[175] & b[193])^(a[174] & b[194])^(a[173] & b[195])^(a[172] & b[196])^(a[171] & b[197])^(a[170] & b[198])^(a[169] & b[199])^(a[168] & b[200])^(a[167] & b[201])^(a[166] & b[202])^(a[165] & b[203])^(a[164] & b[204])^(a[163] & b[205])^(a[162] & b[206])^(a[161] & b[207])^(a[160] & b[208])^(a[159] & b[209])^(a[158] & b[210])^(a[157] & b[211])^(a[156] & b[212])^(a[155] & b[213])^(a[154] & b[214])^(a[153] & b[215])^(a[152] & b[216])^(a[151] & b[217])^(a[150] & b[218])^(a[149] & b[219])^(a[148] & b[220])^(a[147] & b[221])^(a[146] & b[222])^(a[145] & b[223])^(a[144] & b[224])^(a[143] & b[225])^(a[142] & b[226])^(a[141] & b[227])^(a[140] & b[228])^(a[139] & b[229])^(a[138] & b[230])^(a[137] & b[231])^(a[136] & b[232]);
assign y[369] = (a[232] & b[137])^(a[231] & b[138])^(a[230] & b[139])^(a[229] & b[140])^(a[228] & b[141])^(a[227] & b[142])^(a[226] & b[143])^(a[225] & b[144])^(a[224] & b[145])^(a[223] & b[146])^(a[222] & b[147])^(a[221] & b[148])^(a[220] & b[149])^(a[219] & b[150])^(a[218] & b[151])^(a[217] & b[152])^(a[216] & b[153])^(a[215] & b[154])^(a[214] & b[155])^(a[213] & b[156])^(a[212] & b[157])^(a[211] & b[158])^(a[210] & b[159])^(a[209] & b[160])^(a[208] & b[161])^(a[207] & b[162])^(a[206] & b[163])^(a[205] & b[164])^(a[204] & b[165])^(a[203] & b[166])^(a[202] & b[167])^(a[201] & b[168])^(a[200] & b[169])^(a[199] & b[170])^(a[198] & b[171])^(a[197] & b[172])^(a[196] & b[173])^(a[195] & b[174])^(a[194] & b[175])^(a[193] & b[176])^(a[192] & b[177])^(a[191] & b[178])^(a[190] & b[179])^(a[189] & b[180])^(a[188] & b[181])^(a[187] & b[182])^(a[186] & b[183])^(a[185] & b[184])^(a[184] & b[185])^(a[183] & b[186])^(a[182] & b[187])^(a[181] & b[188])^(a[180] & b[189])^(a[179] & b[190])^(a[178] & b[191])^(a[177] & b[192])^(a[176] & b[193])^(a[175] & b[194])^(a[174] & b[195])^(a[173] & b[196])^(a[172] & b[197])^(a[171] & b[198])^(a[170] & b[199])^(a[169] & b[200])^(a[168] & b[201])^(a[167] & b[202])^(a[166] & b[203])^(a[165] & b[204])^(a[164] & b[205])^(a[163] & b[206])^(a[162] & b[207])^(a[161] & b[208])^(a[160] & b[209])^(a[159] & b[210])^(a[158] & b[211])^(a[157] & b[212])^(a[156] & b[213])^(a[155] & b[214])^(a[154] & b[215])^(a[153] & b[216])^(a[152] & b[217])^(a[151] & b[218])^(a[150] & b[219])^(a[149] & b[220])^(a[148] & b[221])^(a[147] & b[222])^(a[146] & b[223])^(a[145] & b[224])^(a[144] & b[225])^(a[143] & b[226])^(a[142] & b[227])^(a[141] & b[228])^(a[140] & b[229])^(a[139] & b[230])^(a[138] & b[231])^(a[137] & b[232]);
assign y[370] = (a[232] & b[138])^(a[231] & b[139])^(a[230] & b[140])^(a[229] & b[141])^(a[228] & b[142])^(a[227] & b[143])^(a[226] & b[144])^(a[225] & b[145])^(a[224] & b[146])^(a[223] & b[147])^(a[222] & b[148])^(a[221] & b[149])^(a[220] & b[150])^(a[219] & b[151])^(a[218] & b[152])^(a[217] & b[153])^(a[216] & b[154])^(a[215] & b[155])^(a[214] & b[156])^(a[213] & b[157])^(a[212] & b[158])^(a[211] & b[159])^(a[210] & b[160])^(a[209] & b[161])^(a[208] & b[162])^(a[207] & b[163])^(a[206] & b[164])^(a[205] & b[165])^(a[204] & b[166])^(a[203] & b[167])^(a[202] & b[168])^(a[201] & b[169])^(a[200] & b[170])^(a[199] & b[171])^(a[198] & b[172])^(a[197] & b[173])^(a[196] & b[174])^(a[195] & b[175])^(a[194] & b[176])^(a[193] & b[177])^(a[192] & b[178])^(a[191] & b[179])^(a[190] & b[180])^(a[189] & b[181])^(a[188] & b[182])^(a[187] & b[183])^(a[186] & b[184])^(a[185] & b[185])^(a[184] & b[186])^(a[183] & b[187])^(a[182] & b[188])^(a[181] & b[189])^(a[180] & b[190])^(a[179] & b[191])^(a[178] & b[192])^(a[177] & b[193])^(a[176] & b[194])^(a[175] & b[195])^(a[174] & b[196])^(a[173] & b[197])^(a[172] & b[198])^(a[171] & b[199])^(a[170] & b[200])^(a[169] & b[201])^(a[168] & b[202])^(a[167] & b[203])^(a[166] & b[204])^(a[165] & b[205])^(a[164] & b[206])^(a[163] & b[207])^(a[162] & b[208])^(a[161] & b[209])^(a[160] & b[210])^(a[159] & b[211])^(a[158] & b[212])^(a[157] & b[213])^(a[156] & b[214])^(a[155] & b[215])^(a[154] & b[216])^(a[153] & b[217])^(a[152] & b[218])^(a[151] & b[219])^(a[150] & b[220])^(a[149] & b[221])^(a[148] & b[222])^(a[147] & b[223])^(a[146] & b[224])^(a[145] & b[225])^(a[144] & b[226])^(a[143] & b[227])^(a[142] & b[228])^(a[141] & b[229])^(a[140] & b[230])^(a[139] & b[231])^(a[138] & b[232]);
assign y[371] = (a[232] & b[139])^(a[231] & b[140])^(a[230] & b[141])^(a[229] & b[142])^(a[228] & b[143])^(a[227] & b[144])^(a[226] & b[145])^(a[225] & b[146])^(a[224] & b[147])^(a[223] & b[148])^(a[222] & b[149])^(a[221] & b[150])^(a[220] & b[151])^(a[219] & b[152])^(a[218] & b[153])^(a[217] & b[154])^(a[216] & b[155])^(a[215] & b[156])^(a[214] & b[157])^(a[213] & b[158])^(a[212] & b[159])^(a[211] & b[160])^(a[210] & b[161])^(a[209] & b[162])^(a[208] & b[163])^(a[207] & b[164])^(a[206] & b[165])^(a[205] & b[166])^(a[204] & b[167])^(a[203] & b[168])^(a[202] & b[169])^(a[201] & b[170])^(a[200] & b[171])^(a[199] & b[172])^(a[198] & b[173])^(a[197] & b[174])^(a[196] & b[175])^(a[195] & b[176])^(a[194] & b[177])^(a[193] & b[178])^(a[192] & b[179])^(a[191] & b[180])^(a[190] & b[181])^(a[189] & b[182])^(a[188] & b[183])^(a[187] & b[184])^(a[186] & b[185])^(a[185] & b[186])^(a[184] & b[187])^(a[183] & b[188])^(a[182] & b[189])^(a[181] & b[190])^(a[180] & b[191])^(a[179] & b[192])^(a[178] & b[193])^(a[177] & b[194])^(a[176] & b[195])^(a[175] & b[196])^(a[174] & b[197])^(a[173] & b[198])^(a[172] & b[199])^(a[171] & b[200])^(a[170] & b[201])^(a[169] & b[202])^(a[168] & b[203])^(a[167] & b[204])^(a[166] & b[205])^(a[165] & b[206])^(a[164] & b[207])^(a[163] & b[208])^(a[162] & b[209])^(a[161] & b[210])^(a[160] & b[211])^(a[159] & b[212])^(a[158] & b[213])^(a[157] & b[214])^(a[156] & b[215])^(a[155] & b[216])^(a[154] & b[217])^(a[153] & b[218])^(a[152] & b[219])^(a[151] & b[220])^(a[150] & b[221])^(a[149] & b[222])^(a[148] & b[223])^(a[147] & b[224])^(a[146] & b[225])^(a[145] & b[226])^(a[144] & b[227])^(a[143] & b[228])^(a[142] & b[229])^(a[141] & b[230])^(a[140] & b[231])^(a[139] & b[232]);
assign y[372] = (a[232] & b[140])^(a[231] & b[141])^(a[230] & b[142])^(a[229] & b[143])^(a[228] & b[144])^(a[227] & b[145])^(a[226] & b[146])^(a[225] & b[147])^(a[224] & b[148])^(a[223] & b[149])^(a[222] & b[150])^(a[221] & b[151])^(a[220] & b[152])^(a[219] & b[153])^(a[218] & b[154])^(a[217] & b[155])^(a[216] & b[156])^(a[215] & b[157])^(a[214] & b[158])^(a[213] & b[159])^(a[212] & b[160])^(a[211] & b[161])^(a[210] & b[162])^(a[209] & b[163])^(a[208] & b[164])^(a[207] & b[165])^(a[206] & b[166])^(a[205] & b[167])^(a[204] & b[168])^(a[203] & b[169])^(a[202] & b[170])^(a[201] & b[171])^(a[200] & b[172])^(a[199] & b[173])^(a[198] & b[174])^(a[197] & b[175])^(a[196] & b[176])^(a[195] & b[177])^(a[194] & b[178])^(a[193] & b[179])^(a[192] & b[180])^(a[191] & b[181])^(a[190] & b[182])^(a[189] & b[183])^(a[188] & b[184])^(a[187] & b[185])^(a[186] & b[186])^(a[185] & b[187])^(a[184] & b[188])^(a[183] & b[189])^(a[182] & b[190])^(a[181] & b[191])^(a[180] & b[192])^(a[179] & b[193])^(a[178] & b[194])^(a[177] & b[195])^(a[176] & b[196])^(a[175] & b[197])^(a[174] & b[198])^(a[173] & b[199])^(a[172] & b[200])^(a[171] & b[201])^(a[170] & b[202])^(a[169] & b[203])^(a[168] & b[204])^(a[167] & b[205])^(a[166] & b[206])^(a[165] & b[207])^(a[164] & b[208])^(a[163] & b[209])^(a[162] & b[210])^(a[161] & b[211])^(a[160] & b[212])^(a[159] & b[213])^(a[158] & b[214])^(a[157] & b[215])^(a[156] & b[216])^(a[155] & b[217])^(a[154] & b[218])^(a[153] & b[219])^(a[152] & b[220])^(a[151] & b[221])^(a[150] & b[222])^(a[149] & b[223])^(a[148] & b[224])^(a[147] & b[225])^(a[146] & b[226])^(a[145] & b[227])^(a[144] & b[228])^(a[143] & b[229])^(a[142] & b[230])^(a[141] & b[231])^(a[140] & b[232]);
assign y[373] = (a[232] & b[141])^(a[231] & b[142])^(a[230] & b[143])^(a[229] & b[144])^(a[228] & b[145])^(a[227] & b[146])^(a[226] & b[147])^(a[225] & b[148])^(a[224] & b[149])^(a[223] & b[150])^(a[222] & b[151])^(a[221] & b[152])^(a[220] & b[153])^(a[219] & b[154])^(a[218] & b[155])^(a[217] & b[156])^(a[216] & b[157])^(a[215] & b[158])^(a[214] & b[159])^(a[213] & b[160])^(a[212] & b[161])^(a[211] & b[162])^(a[210] & b[163])^(a[209] & b[164])^(a[208] & b[165])^(a[207] & b[166])^(a[206] & b[167])^(a[205] & b[168])^(a[204] & b[169])^(a[203] & b[170])^(a[202] & b[171])^(a[201] & b[172])^(a[200] & b[173])^(a[199] & b[174])^(a[198] & b[175])^(a[197] & b[176])^(a[196] & b[177])^(a[195] & b[178])^(a[194] & b[179])^(a[193] & b[180])^(a[192] & b[181])^(a[191] & b[182])^(a[190] & b[183])^(a[189] & b[184])^(a[188] & b[185])^(a[187] & b[186])^(a[186] & b[187])^(a[185] & b[188])^(a[184] & b[189])^(a[183] & b[190])^(a[182] & b[191])^(a[181] & b[192])^(a[180] & b[193])^(a[179] & b[194])^(a[178] & b[195])^(a[177] & b[196])^(a[176] & b[197])^(a[175] & b[198])^(a[174] & b[199])^(a[173] & b[200])^(a[172] & b[201])^(a[171] & b[202])^(a[170] & b[203])^(a[169] & b[204])^(a[168] & b[205])^(a[167] & b[206])^(a[166] & b[207])^(a[165] & b[208])^(a[164] & b[209])^(a[163] & b[210])^(a[162] & b[211])^(a[161] & b[212])^(a[160] & b[213])^(a[159] & b[214])^(a[158] & b[215])^(a[157] & b[216])^(a[156] & b[217])^(a[155] & b[218])^(a[154] & b[219])^(a[153] & b[220])^(a[152] & b[221])^(a[151] & b[222])^(a[150] & b[223])^(a[149] & b[224])^(a[148] & b[225])^(a[147] & b[226])^(a[146] & b[227])^(a[145] & b[228])^(a[144] & b[229])^(a[143] & b[230])^(a[142] & b[231])^(a[141] & b[232]);
assign y[374] = (a[232] & b[142])^(a[231] & b[143])^(a[230] & b[144])^(a[229] & b[145])^(a[228] & b[146])^(a[227] & b[147])^(a[226] & b[148])^(a[225] & b[149])^(a[224] & b[150])^(a[223] & b[151])^(a[222] & b[152])^(a[221] & b[153])^(a[220] & b[154])^(a[219] & b[155])^(a[218] & b[156])^(a[217] & b[157])^(a[216] & b[158])^(a[215] & b[159])^(a[214] & b[160])^(a[213] & b[161])^(a[212] & b[162])^(a[211] & b[163])^(a[210] & b[164])^(a[209] & b[165])^(a[208] & b[166])^(a[207] & b[167])^(a[206] & b[168])^(a[205] & b[169])^(a[204] & b[170])^(a[203] & b[171])^(a[202] & b[172])^(a[201] & b[173])^(a[200] & b[174])^(a[199] & b[175])^(a[198] & b[176])^(a[197] & b[177])^(a[196] & b[178])^(a[195] & b[179])^(a[194] & b[180])^(a[193] & b[181])^(a[192] & b[182])^(a[191] & b[183])^(a[190] & b[184])^(a[189] & b[185])^(a[188] & b[186])^(a[187] & b[187])^(a[186] & b[188])^(a[185] & b[189])^(a[184] & b[190])^(a[183] & b[191])^(a[182] & b[192])^(a[181] & b[193])^(a[180] & b[194])^(a[179] & b[195])^(a[178] & b[196])^(a[177] & b[197])^(a[176] & b[198])^(a[175] & b[199])^(a[174] & b[200])^(a[173] & b[201])^(a[172] & b[202])^(a[171] & b[203])^(a[170] & b[204])^(a[169] & b[205])^(a[168] & b[206])^(a[167] & b[207])^(a[166] & b[208])^(a[165] & b[209])^(a[164] & b[210])^(a[163] & b[211])^(a[162] & b[212])^(a[161] & b[213])^(a[160] & b[214])^(a[159] & b[215])^(a[158] & b[216])^(a[157] & b[217])^(a[156] & b[218])^(a[155] & b[219])^(a[154] & b[220])^(a[153] & b[221])^(a[152] & b[222])^(a[151] & b[223])^(a[150] & b[224])^(a[149] & b[225])^(a[148] & b[226])^(a[147] & b[227])^(a[146] & b[228])^(a[145] & b[229])^(a[144] & b[230])^(a[143] & b[231])^(a[142] & b[232]);
assign y[375] = (a[232] & b[143])^(a[231] & b[144])^(a[230] & b[145])^(a[229] & b[146])^(a[228] & b[147])^(a[227] & b[148])^(a[226] & b[149])^(a[225] & b[150])^(a[224] & b[151])^(a[223] & b[152])^(a[222] & b[153])^(a[221] & b[154])^(a[220] & b[155])^(a[219] & b[156])^(a[218] & b[157])^(a[217] & b[158])^(a[216] & b[159])^(a[215] & b[160])^(a[214] & b[161])^(a[213] & b[162])^(a[212] & b[163])^(a[211] & b[164])^(a[210] & b[165])^(a[209] & b[166])^(a[208] & b[167])^(a[207] & b[168])^(a[206] & b[169])^(a[205] & b[170])^(a[204] & b[171])^(a[203] & b[172])^(a[202] & b[173])^(a[201] & b[174])^(a[200] & b[175])^(a[199] & b[176])^(a[198] & b[177])^(a[197] & b[178])^(a[196] & b[179])^(a[195] & b[180])^(a[194] & b[181])^(a[193] & b[182])^(a[192] & b[183])^(a[191] & b[184])^(a[190] & b[185])^(a[189] & b[186])^(a[188] & b[187])^(a[187] & b[188])^(a[186] & b[189])^(a[185] & b[190])^(a[184] & b[191])^(a[183] & b[192])^(a[182] & b[193])^(a[181] & b[194])^(a[180] & b[195])^(a[179] & b[196])^(a[178] & b[197])^(a[177] & b[198])^(a[176] & b[199])^(a[175] & b[200])^(a[174] & b[201])^(a[173] & b[202])^(a[172] & b[203])^(a[171] & b[204])^(a[170] & b[205])^(a[169] & b[206])^(a[168] & b[207])^(a[167] & b[208])^(a[166] & b[209])^(a[165] & b[210])^(a[164] & b[211])^(a[163] & b[212])^(a[162] & b[213])^(a[161] & b[214])^(a[160] & b[215])^(a[159] & b[216])^(a[158] & b[217])^(a[157] & b[218])^(a[156] & b[219])^(a[155] & b[220])^(a[154] & b[221])^(a[153] & b[222])^(a[152] & b[223])^(a[151] & b[224])^(a[150] & b[225])^(a[149] & b[226])^(a[148] & b[227])^(a[147] & b[228])^(a[146] & b[229])^(a[145] & b[230])^(a[144] & b[231])^(a[143] & b[232]);
assign y[376] = (a[232] & b[144])^(a[231] & b[145])^(a[230] & b[146])^(a[229] & b[147])^(a[228] & b[148])^(a[227] & b[149])^(a[226] & b[150])^(a[225] & b[151])^(a[224] & b[152])^(a[223] & b[153])^(a[222] & b[154])^(a[221] & b[155])^(a[220] & b[156])^(a[219] & b[157])^(a[218] & b[158])^(a[217] & b[159])^(a[216] & b[160])^(a[215] & b[161])^(a[214] & b[162])^(a[213] & b[163])^(a[212] & b[164])^(a[211] & b[165])^(a[210] & b[166])^(a[209] & b[167])^(a[208] & b[168])^(a[207] & b[169])^(a[206] & b[170])^(a[205] & b[171])^(a[204] & b[172])^(a[203] & b[173])^(a[202] & b[174])^(a[201] & b[175])^(a[200] & b[176])^(a[199] & b[177])^(a[198] & b[178])^(a[197] & b[179])^(a[196] & b[180])^(a[195] & b[181])^(a[194] & b[182])^(a[193] & b[183])^(a[192] & b[184])^(a[191] & b[185])^(a[190] & b[186])^(a[189] & b[187])^(a[188] & b[188])^(a[187] & b[189])^(a[186] & b[190])^(a[185] & b[191])^(a[184] & b[192])^(a[183] & b[193])^(a[182] & b[194])^(a[181] & b[195])^(a[180] & b[196])^(a[179] & b[197])^(a[178] & b[198])^(a[177] & b[199])^(a[176] & b[200])^(a[175] & b[201])^(a[174] & b[202])^(a[173] & b[203])^(a[172] & b[204])^(a[171] & b[205])^(a[170] & b[206])^(a[169] & b[207])^(a[168] & b[208])^(a[167] & b[209])^(a[166] & b[210])^(a[165] & b[211])^(a[164] & b[212])^(a[163] & b[213])^(a[162] & b[214])^(a[161] & b[215])^(a[160] & b[216])^(a[159] & b[217])^(a[158] & b[218])^(a[157] & b[219])^(a[156] & b[220])^(a[155] & b[221])^(a[154] & b[222])^(a[153] & b[223])^(a[152] & b[224])^(a[151] & b[225])^(a[150] & b[226])^(a[149] & b[227])^(a[148] & b[228])^(a[147] & b[229])^(a[146] & b[230])^(a[145] & b[231])^(a[144] & b[232]);
assign y[377] = (a[232] & b[145])^(a[231] & b[146])^(a[230] & b[147])^(a[229] & b[148])^(a[228] & b[149])^(a[227] & b[150])^(a[226] & b[151])^(a[225] & b[152])^(a[224] & b[153])^(a[223] & b[154])^(a[222] & b[155])^(a[221] & b[156])^(a[220] & b[157])^(a[219] & b[158])^(a[218] & b[159])^(a[217] & b[160])^(a[216] & b[161])^(a[215] & b[162])^(a[214] & b[163])^(a[213] & b[164])^(a[212] & b[165])^(a[211] & b[166])^(a[210] & b[167])^(a[209] & b[168])^(a[208] & b[169])^(a[207] & b[170])^(a[206] & b[171])^(a[205] & b[172])^(a[204] & b[173])^(a[203] & b[174])^(a[202] & b[175])^(a[201] & b[176])^(a[200] & b[177])^(a[199] & b[178])^(a[198] & b[179])^(a[197] & b[180])^(a[196] & b[181])^(a[195] & b[182])^(a[194] & b[183])^(a[193] & b[184])^(a[192] & b[185])^(a[191] & b[186])^(a[190] & b[187])^(a[189] & b[188])^(a[188] & b[189])^(a[187] & b[190])^(a[186] & b[191])^(a[185] & b[192])^(a[184] & b[193])^(a[183] & b[194])^(a[182] & b[195])^(a[181] & b[196])^(a[180] & b[197])^(a[179] & b[198])^(a[178] & b[199])^(a[177] & b[200])^(a[176] & b[201])^(a[175] & b[202])^(a[174] & b[203])^(a[173] & b[204])^(a[172] & b[205])^(a[171] & b[206])^(a[170] & b[207])^(a[169] & b[208])^(a[168] & b[209])^(a[167] & b[210])^(a[166] & b[211])^(a[165] & b[212])^(a[164] & b[213])^(a[163] & b[214])^(a[162] & b[215])^(a[161] & b[216])^(a[160] & b[217])^(a[159] & b[218])^(a[158] & b[219])^(a[157] & b[220])^(a[156] & b[221])^(a[155] & b[222])^(a[154] & b[223])^(a[153] & b[224])^(a[152] & b[225])^(a[151] & b[226])^(a[150] & b[227])^(a[149] & b[228])^(a[148] & b[229])^(a[147] & b[230])^(a[146] & b[231])^(a[145] & b[232]);
assign y[378] = (a[232] & b[146])^(a[231] & b[147])^(a[230] & b[148])^(a[229] & b[149])^(a[228] & b[150])^(a[227] & b[151])^(a[226] & b[152])^(a[225] & b[153])^(a[224] & b[154])^(a[223] & b[155])^(a[222] & b[156])^(a[221] & b[157])^(a[220] & b[158])^(a[219] & b[159])^(a[218] & b[160])^(a[217] & b[161])^(a[216] & b[162])^(a[215] & b[163])^(a[214] & b[164])^(a[213] & b[165])^(a[212] & b[166])^(a[211] & b[167])^(a[210] & b[168])^(a[209] & b[169])^(a[208] & b[170])^(a[207] & b[171])^(a[206] & b[172])^(a[205] & b[173])^(a[204] & b[174])^(a[203] & b[175])^(a[202] & b[176])^(a[201] & b[177])^(a[200] & b[178])^(a[199] & b[179])^(a[198] & b[180])^(a[197] & b[181])^(a[196] & b[182])^(a[195] & b[183])^(a[194] & b[184])^(a[193] & b[185])^(a[192] & b[186])^(a[191] & b[187])^(a[190] & b[188])^(a[189] & b[189])^(a[188] & b[190])^(a[187] & b[191])^(a[186] & b[192])^(a[185] & b[193])^(a[184] & b[194])^(a[183] & b[195])^(a[182] & b[196])^(a[181] & b[197])^(a[180] & b[198])^(a[179] & b[199])^(a[178] & b[200])^(a[177] & b[201])^(a[176] & b[202])^(a[175] & b[203])^(a[174] & b[204])^(a[173] & b[205])^(a[172] & b[206])^(a[171] & b[207])^(a[170] & b[208])^(a[169] & b[209])^(a[168] & b[210])^(a[167] & b[211])^(a[166] & b[212])^(a[165] & b[213])^(a[164] & b[214])^(a[163] & b[215])^(a[162] & b[216])^(a[161] & b[217])^(a[160] & b[218])^(a[159] & b[219])^(a[158] & b[220])^(a[157] & b[221])^(a[156] & b[222])^(a[155] & b[223])^(a[154] & b[224])^(a[153] & b[225])^(a[152] & b[226])^(a[151] & b[227])^(a[150] & b[228])^(a[149] & b[229])^(a[148] & b[230])^(a[147] & b[231])^(a[146] & b[232]);
assign y[379] = (a[232] & b[147])^(a[231] & b[148])^(a[230] & b[149])^(a[229] & b[150])^(a[228] & b[151])^(a[227] & b[152])^(a[226] & b[153])^(a[225] & b[154])^(a[224] & b[155])^(a[223] & b[156])^(a[222] & b[157])^(a[221] & b[158])^(a[220] & b[159])^(a[219] & b[160])^(a[218] & b[161])^(a[217] & b[162])^(a[216] & b[163])^(a[215] & b[164])^(a[214] & b[165])^(a[213] & b[166])^(a[212] & b[167])^(a[211] & b[168])^(a[210] & b[169])^(a[209] & b[170])^(a[208] & b[171])^(a[207] & b[172])^(a[206] & b[173])^(a[205] & b[174])^(a[204] & b[175])^(a[203] & b[176])^(a[202] & b[177])^(a[201] & b[178])^(a[200] & b[179])^(a[199] & b[180])^(a[198] & b[181])^(a[197] & b[182])^(a[196] & b[183])^(a[195] & b[184])^(a[194] & b[185])^(a[193] & b[186])^(a[192] & b[187])^(a[191] & b[188])^(a[190] & b[189])^(a[189] & b[190])^(a[188] & b[191])^(a[187] & b[192])^(a[186] & b[193])^(a[185] & b[194])^(a[184] & b[195])^(a[183] & b[196])^(a[182] & b[197])^(a[181] & b[198])^(a[180] & b[199])^(a[179] & b[200])^(a[178] & b[201])^(a[177] & b[202])^(a[176] & b[203])^(a[175] & b[204])^(a[174] & b[205])^(a[173] & b[206])^(a[172] & b[207])^(a[171] & b[208])^(a[170] & b[209])^(a[169] & b[210])^(a[168] & b[211])^(a[167] & b[212])^(a[166] & b[213])^(a[165] & b[214])^(a[164] & b[215])^(a[163] & b[216])^(a[162] & b[217])^(a[161] & b[218])^(a[160] & b[219])^(a[159] & b[220])^(a[158] & b[221])^(a[157] & b[222])^(a[156] & b[223])^(a[155] & b[224])^(a[154] & b[225])^(a[153] & b[226])^(a[152] & b[227])^(a[151] & b[228])^(a[150] & b[229])^(a[149] & b[230])^(a[148] & b[231])^(a[147] & b[232]);
assign y[380] = (a[232] & b[148])^(a[231] & b[149])^(a[230] & b[150])^(a[229] & b[151])^(a[228] & b[152])^(a[227] & b[153])^(a[226] & b[154])^(a[225] & b[155])^(a[224] & b[156])^(a[223] & b[157])^(a[222] & b[158])^(a[221] & b[159])^(a[220] & b[160])^(a[219] & b[161])^(a[218] & b[162])^(a[217] & b[163])^(a[216] & b[164])^(a[215] & b[165])^(a[214] & b[166])^(a[213] & b[167])^(a[212] & b[168])^(a[211] & b[169])^(a[210] & b[170])^(a[209] & b[171])^(a[208] & b[172])^(a[207] & b[173])^(a[206] & b[174])^(a[205] & b[175])^(a[204] & b[176])^(a[203] & b[177])^(a[202] & b[178])^(a[201] & b[179])^(a[200] & b[180])^(a[199] & b[181])^(a[198] & b[182])^(a[197] & b[183])^(a[196] & b[184])^(a[195] & b[185])^(a[194] & b[186])^(a[193] & b[187])^(a[192] & b[188])^(a[191] & b[189])^(a[190] & b[190])^(a[189] & b[191])^(a[188] & b[192])^(a[187] & b[193])^(a[186] & b[194])^(a[185] & b[195])^(a[184] & b[196])^(a[183] & b[197])^(a[182] & b[198])^(a[181] & b[199])^(a[180] & b[200])^(a[179] & b[201])^(a[178] & b[202])^(a[177] & b[203])^(a[176] & b[204])^(a[175] & b[205])^(a[174] & b[206])^(a[173] & b[207])^(a[172] & b[208])^(a[171] & b[209])^(a[170] & b[210])^(a[169] & b[211])^(a[168] & b[212])^(a[167] & b[213])^(a[166] & b[214])^(a[165] & b[215])^(a[164] & b[216])^(a[163] & b[217])^(a[162] & b[218])^(a[161] & b[219])^(a[160] & b[220])^(a[159] & b[221])^(a[158] & b[222])^(a[157] & b[223])^(a[156] & b[224])^(a[155] & b[225])^(a[154] & b[226])^(a[153] & b[227])^(a[152] & b[228])^(a[151] & b[229])^(a[150] & b[230])^(a[149] & b[231])^(a[148] & b[232]);
assign y[381] = (a[232] & b[149])^(a[231] & b[150])^(a[230] & b[151])^(a[229] & b[152])^(a[228] & b[153])^(a[227] & b[154])^(a[226] & b[155])^(a[225] & b[156])^(a[224] & b[157])^(a[223] & b[158])^(a[222] & b[159])^(a[221] & b[160])^(a[220] & b[161])^(a[219] & b[162])^(a[218] & b[163])^(a[217] & b[164])^(a[216] & b[165])^(a[215] & b[166])^(a[214] & b[167])^(a[213] & b[168])^(a[212] & b[169])^(a[211] & b[170])^(a[210] & b[171])^(a[209] & b[172])^(a[208] & b[173])^(a[207] & b[174])^(a[206] & b[175])^(a[205] & b[176])^(a[204] & b[177])^(a[203] & b[178])^(a[202] & b[179])^(a[201] & b[180])^(a[200] & b[181])^(a[199] & b[182])^(a[198] & b[183])^(a[197] & b[184])^(a[196] & b[185])^(a[195] & b[186])^(a[194] & b[187])^(a[193] & b[188])^(a[192] & b[189])^(a[191] & b[190])^(a[190] & b[191])^(a[189] & b[192])^(a[188] & b[193])^(a[187] & b[194])^(a[186] & b[195])^(a[185] & b[196])^(a[184] & b[197])^(a[183] & b[198])^(a[182] & b[199])^(a[181] & b[200])^(a[180] & b[201])^(a[179] & b[202])^(a[178] & b[203])^(a[177] & b[204])^(a[176] & b[205])^(a[175] & b[206])^(a[174] & b[207])^(a[173] & b[208])^(a[172] & b[209])^(a[171] & b[210])^(a[170] & b[211])^(a[169] & b[212])^(a[168] & b[213])^(a[167] & b[214])^(a[166] & b[215])^(a[165] & b[216])^(a[164] & b[217])^(a[163] & b[218])^(a[162] & b[219])^(a[161] & b[220])^(a[160] & b[221])^(a[159] & b[222])^(a[158] & b[223])^(a[157] & b[224])^(a[156] & b[225])^(a[155] & b[226])^(a[154] & b[227])^(a[153] & b[228])^(a[152] & b[229])^(a[151] & b[230])^(a[150] & b[231])^(a[149] & b[232]);
assign y[382] = (a[232] & b[150])^(a[231] & b[151])^(a[230] & b[152])^(a[229] & b[153])^(a[228] & b[154])^(a[227] & b[155])^(a[226] & b[156])^(a[225] & b[157])^(a[224] & b[158])^(a[223] & b[159])^(a[222] & b[160])^(a[221] & b[161])^(a[220] & b[162])^(a[219] & b[163])^(a[218] & b[164])^(a[217] & b[165])^(a[216] & b[166])^(a[215] & b[167])^(a[214] & b[168])^(a[213] & b[169])^(a[212] & b[170])^(a[211] & b[171])^(a[210] & b[172])^(a[209] & b[173])^(a[208] & b[174])^(a[207] & b[175])^(a[206] & b[176])^(a[205] & b[177])^(a[204] & b[178])^(a[203] & b[179])^(a[202] & b[180])^(a[201] & b[181])^(a[200] & b[182])^(a[199] & b[183])^(a[198] & b[184])^(a[197] & b[185])^(a[196] & b[186])^(a[195] & b[187])^(a[194] & b[188])^(a[193] & b[189])^(a[192] & b[190])^(a[191] & b[191])^(a[190] & b[192])^(a[189] & b[193])^(a[188] & b[194])^(a[187] & b[195])^(a[186] & b[196])^(a[185] & b[197])^(a[184] & b[198])^(a[183] & b[199])^(a[182] & b[200])^(a[181] & b[201])^(a[180] & b[202])^(a[179] & b[203])^(a[178] & b[204])^(a[177] & b[205])^(a[176] & b[206])^(a[175] & b[207])^(a[174] & b[208])^(a[173] & b[209])^(a[172] & b[210])^(a[171] & b[211])^(a[170] & b[212])^(a[169] & b[213])^(a[168] & b[214])^(a[167] & b[215])^(a[166] & b[216])^(a[165] & b[217])^(a[164] & b[218])^(a[163] & b[219])^(a[162] & b[220])^(a[161] & b[221])^(a[160] & b[222])^(a[159] & b[223])^(a[158] & b[224])^(a[157] & b[225])^(a[156] & b[226])^(a[155] & b[227])^(a[154] & b[228])^(a[153] & b[229])^(a[152] & b[230])^(a[151] & b[231])^(a[150] & b[232]);
assign y[383] = (a[232] & b[151])^(a[231] & b[152])^(a[230] & b[153])^(a[229] & b[154])^(a[228] & b[155])^(a[227] & b[156])^(a[226] & b[157])^(a[225] & b[158])^(a[224] & b[159])^(a[223] & b[160])^(a[222] & b[161])^(a[221] & b[162])^(a[220] & b[163])^(a[219] & b[164])^(a[218] & b[165])^(a[217] & b[166])^(a[216] & b[167])^(a[215] & b[168])^(a[214] & b[169])^(a[213] & b[170])^(a[212] & b[171])^(a[211] & b[172])^(a[210] & b[173])^(a[209] & b[174])^(a[208] & b[175])^(a[207] & b[176])^(a[206] & b[177])^(a[205] & b[178])^(a[204] & b[179])^(a[203] & b[180])^(a[202] & b[181])^(a[201] & b[182])^(a[200] & b[183])^(a[199] & b[184])^(a[198] & b[185])^(a[197] & b[186])^(a[196] & b[187])^(a[195] & b[188])^(a[194] & b[189])^(a[193] & b[190])^(a[192] & b[191])^(a[191] & b[192])^(a[190] & b[193])^(a[189] & b[194])^(a[188] & b[195])^(a[187] & b[196])^(a[186] & b[197])^(a[185] & b[198])^(a[184] & b[199])^(a[183] & b[200])^(a[182] & b[201])^(a[181] & b[202])^(a[180] & b[203])^(a[179] & b[204])^(a[178] & b[205])^(a[177] & b[206])^(a[176] & b[207])^(a[175] & b[208])^(a[174] & b[209])^(a[173] & b[210])^(a[172] & b[211])^(a[171] & b[212])^(a[170] & b[213])^(a[169] & b[214])^(a[168] & b[215])^(a[167] & b[216])^(a[166] & b[217])^(a[165] & b[218])^(a[164] & b[219])^(a[163] & b[220])^(a[162] & b[221])^(a[161] & b[222])^(a[160] & b[223])^(a[159] & b[224])^(a[158] & b[225])^(a[157] & b[226])^(a[156] & b[227])^(a[155] & b[228])^(a[154] & b[229])^(a[153] & b[230])^(a[152] & b[231])^(a[151] & b[232]);
assign y[384] = (a[232] & b[152])^(a[231] & b[153])^(a[230] & b[154])^(a[229] & b[155])^(a[228] & b[156])^(a[227] & b[157])^(a[226] & b[158])^(a[225] & b[159])^(a[224] & b[160])^(a[223] & b[161])^(a[222] & b[162])^(a[221] & b[163])^(a[220] & b[164])^(a[219] & b[165])^(a[218] & b[166])^(a[217] & b[167])^(a[216] & b[168])^(a[215] & b[169])^(a[214] & b[170])^(a[213] & b[171])^(a[212] & b[172])^(a[211] & b[173])^(a[210] & b[174])^(a[209] & b[175])^(a[208] & b[176])^(a[207] & b[177])^(a[206] & b[178])^(a[205] & b[179])^(a[204] & b[180])^(a[203] & b[181])^(a[202] & b[182])^(a[201] & b[183])^(a[200] & b[184])^(a[199] & b[185])^(a[198] & b[186])^(a[197] & b[187])^(a[196] & b[188])^(a[195] & b[189])^(a[194] & b[190])^(a[193] & b[191])^(a[192] & b[192])^(a[191] & b[193])^(a[190] & b[194])^(a[189] & b[195])^(a[188] & b[196])^(a[187] & b[197])^(a[186] & b[198])^(a[185] & b[199])^(a[184] & b[200])^(a[183] & b[201])^(a[182] & b[202])^(a[181] & b[203])^(a[180] & b[204])^(a[179] & b[205])^(a[178] & b[206])^(a[177] & b[207])^(a[176] & b[208])^(a[175] & b[209])^(a[174] & b[210])^(a[173] & b[211])^(a[172] & b[212])^(a[171] & b[213])^(a[170] & b[214])^(a[169] & b[215])^(a[168] & b[216])^(a[167] & b[217])^(a[166] & b[218])^(a[165] & b[219])^(a[164] & b[220])^(a[163] & b[221])^(a[162] & b[222])^(a[161] & b[223])^(a[160] & b[224])^(a[159] & b[225])^(a[158] & b[226])^(a[157] & b[227])^(a[156] & b[228])^(a[155] & b[229])^(a[154] & b[230])^(a[153] & b[231])^(a[152] & b[232]);
assign y[385] = (a[232] & b[153])^(a[231] & b[154])^(a[230] & b[155])^(a[229] & b[156])^(a[228] & b[157])^(a[227] & b[158])^(a[226] & b[159])^(a[225] & b[160])^(a[224] & b[161])^(a[223] & b[162])^(a[222] & b[163])^(a[221] & b[164])^(a[220] & b[165])^(a[219] & b[166])^(a[218] & b[167])^(a[217] & b[168])^(a[216] & b[169])^(a[215] & b[170])^(a[214] & b[171])^(a[213] & b[172])^(a[212] & b[173])^(a[211] & b[174])^(a[210] & b[175])^(a[209] & b[176])^(a[208] & b[177])^(a[207] & b[178])^(a[206] & b[179])^(a[205] & b[180])^(a[204] & b[181])^(a[203] & b[182])^(a[202] & b[183])^(a[201] & b[184])^(a[200] & b[185])^(a[199] & b[186])^(a[198] & b[187])^(a[197] & b[188])^(a[196] & b[189])^(a[195] & b[190])^(a[194] & b[191])^(a[193] & b[192])^(a[192] & b[193])^(a[191] & b[194])^(a[190] & b[195])^(a[189] & b[196])^(a[188] & b[197])^(a[187] & b[198])^(a[186] & b[199])^(a[185] & b[200])^(a[184] & b[201])^(a[183] & b[202])^(a[182] & b[203])^(a[181] & b[204])^(a[180] & b[205])^(a[179] & b[206])^(a[178] & b[207])^(a[177] & b[208])^(a[176] & b[209])^(a[175] & b[210])^(a[174] & b[211])^(a[173] & b[212])^(a[172] & b[213])^(a[171] & b[214])^(a[170] & b[215])^(a[169] & b[216])^(a[168] & b[217])^(a[167] & b[218])^(a[166] & b[219])^(a[165] & b[220])^(a[164] & b[221])^(a[163] & b[222])^(a[162] & b[223])^(a[161] & b[224])^(a[160] & b[225])^(a[159] & b[226])^(a[158] & b[227])^(a[157] & b[228])^(a[156] & b[229])^(a[155] & b[230])^(a[154] & b[231])^(a[153] & b[232]);
assign y[386] = (a[232] & b[154])^(a[231] & b[155])^(a[230] & b[156])^(a[229] & b[157])^(a[228] & b[158])^(a[227] & b[159])^(a[226] & b[160])^(a[225] & b[161])^(a[224] & b[162])^(a[223] & b[163])^(a[222] & b[164])^(a[221] & b[165])^(a[220] & b[166])^(a[219] & b[167])^(a[218] & b[168])^(a[217] & b[169])^(a[216] & b[170])^(a[215] & b[171])^(a[214] & b[172])^(a[213] & b[173])^(a[212] & b[174])^(a[211] & b[175])^(a[210] & b[176])^(a[209] & b[177])^(a[208] & b[178])^(a[207] & b[179])^(a[206] & b[180])^(a[205] & b[181])^(a[204] & b[182])^(a[203] & b[183])^(a[202] & b[184])^(a[201] & b[185])^(a[200] & b[186])^(a[199] & b[187])^(a[198] & b[188])^(a[197] & b[189])^(a[196] & b[190])^(a[195] & b[191])^(a[194] & b[192])^(a[193] & b[193])^(a[192] & b[194])^(a[191] & b[195])^(a[190] & b[196])^(a[189] & b[197])^(a[188] & b[198])^(a[187] & b[199])^(a[186] & b[200])^(a[185] & b[201])^(a[184] & b[202])^(a[183] & b[203])^(a[182] & b[204])^(a[181] & b[205])^(a[180] & b[206])^(a[179] & b[207])^(a[178] & b[208])^(a[177] & b[209])^(a[176] & b[210])^(a[175] & b[211])^(a[174] & b[212])^(a[173] & b[213])^(a[172] & b[214])^(a[171] & b[215])^(a[170] & b[216])^(a[169] & b[217])^(a[168] & b[218])^(a[167] & b[219])^(a[166] & b[220])^(a[165] & b[221])^(a[164] & b[222])^(a[163] & b[223])^(a[162] & b[224])^(a[161] & b[225])^(a[160] & b[226])^(a[159] & b[227])^(a[158] & b[228])^(a[157] & b[229])^(a[156] & b[230])^(a[155] & b[231])^(a[154] & b[232]);
assign y[387] = (a[232] & b[155])^(a[231] & b[156])^(a[230] & b[157])^(a[229] & b[158])^(a[228] & b[159])^(a[227] & b[160])^(a[226] & b[161])^(a[225] & b[162])^(a[224] & b[163])^(a[223] & b[164])^(a[222] & b[165])^(a[221] & b[166])^(a[220] & b[167])^(a[219] & b[168])^(a[218] & b[169])^(a[217] & b[170])^(a[216] & b[171])^(a[215] & b[172])^(a[214] & b[173])^(a[213] & b[174])^(a[212] & b[175])^(a[211] & b[176])^(a[210] & b[177])^(a[209] & b[178])^(a[208] & b[179])^(a[207] & b[180])^(a[206] & b[181])^(a[205] & b[182])^(a[204] & b[183])^(a[203] & b[184])^(a[202] & b[185])^(a[201] & b[186])^(a[200] & b[187])^(a[199] & b[188])^(a[198] & b[189])^(a[197] & b[190])^(a[196] & b[191])^(a[195] & b[192])^(a[194] & b[193])^(a[193] & b[194])^(a[192] & b[195])^(a[191] & b[196])^(a[190] & b[197])^(a[189] & b[198])^(a[188] & b[199])^(a[187] & b[200])^(a[186] & b[201])^(a[185] & b[202])^(a[184] & b[203])^(a[183] & b[204])^(a[182] & b[205])^(a[181] & b[206])^(a[180] & b[207])^(a[179] & b[208])^(a[178] & b[209])^(a[177] & b[210])^(a[176] & b[211])^(a[175] & b[212])^(a[174] & b[213])^(a[173] & b[214])^(a[172] & b[215])^(a[171] & b[216])^(a[170] & b[217])^(a[169] & b[218])^(a[168] & b[219])^(a[167] & b[220])^(a[166] & b[221])^(a[165] & b[222])^(a[164] & b[223])^(a[163] & b[224])^(a[162] & b[225])^(a[161] & b[226])^(a[160] & b[227])^(a[159] & b[228])^(a[158] & b[229])^(a[157] & b[230])^(a[156] & b[231])^(a[155] & b[232]);
assign y[388] = (a[232] & b[156])^(a[231] & b[157])^(a[230] & b[158])^(a[229] & b[159])^(a[228] & b[160])^(a[227] & b[161])^(a[226] & b[162])^(a[225] & b[163])^(a[224] & b[164])^(a[223] & b[165])^(a[222] & b[166])^(a[221] & b[167])^(a[220] & b[168])^(a[219] & b[169])^(a[218] & b[170])^(a[217] & b[171])^(a[216] & b[172])^(a[215] & b[173])^(a[214] & b[174])^(a[213] & b[175])^(a[212] & b[176])^(a[211] & b[177])^(a[210] & b[178])^(a[209] & b[179])^(a[208] & b[180])^(a[207] & b[181])^(a[206] & b[182])^(a[205] & b[183])^(a[204] & b[184])^(a[203] & b[185])^(a[202] & b[186])^(a[201] & b[187])^(a[200] & b[188])^(a[199] & b[189])^(a[198] & b[190])^(a[197] & b[191])^(a[196] & b[192])^(a[195] & b[193])^(a[194] & b[194])^(a[193] & b[195])^(a[192] & b[196])^(a[191] & b[197])^(a[190] & b[198])^(a[189] & b[199])^(a[188] & b[200])^(a[187] & b[201])^(a[186] & b[202])^(a[185] & b[203])^(a[184] & b[204])^(a[183] & b[205])^(a[182] & b[206])^(a[181] & b[207])^(a[180] & b[208])^(a[179] & b[209])^(a[178] & b[210])^(a[177] & b[211])^(a[176] & b[212])^(a[175] & b[213])^(a[174] & b[214])^(a[173] & b[215])^(a[172] & b[216])^(a[171] & b[217])^(a[170] & b[218])^(a[169] & b[219])^(a[168] & b[220])^(a[167] & b[221])^(a[166] & b[222])^(a[165] & b[223])^(a[164] & b[224])^(a[163] & b[225])^(a[162] & b[226])^(a[161] & b[227])^(a[160] & b[228])^(a[159] & b[229])^(a[158] & b[230])^(a[157] & b[231])^(a[156] & b[232]);
assign y[389] = (a[232] & b[157])^(a[231] & b[158])^(a[230] & b[159])^(a[229] & b[160])^(a[228] & b[161])^(a[227] & b[162])^(a[226] & b[163])^(a[225] & b[164])^(a[224] & b[165])^(a[223] & b[166])^(a[222] & b[167])^(a[221] & b[168])^(a[220] & b[169])^(a[219] & b[170])^(a[218] & b[171])^(a[217] & b[172])^(a[216] & b[173])^(a[215] & b[174])^(a[214] & b[175])^(a[213] & b[176])^(a[212] & b[177])^(a[211] & b[178])^(a[210] & b[179])^(a[209] & b[180])^(a[208] & b[181])^(a[207] & b[182])^(a[206] & b[183])^(a[205] & b[184])^(a[204] & b[185])^(a[203] & b[186])^(a[202] & b[187])^(a[201] & b[188])^(a[200] & b[189])^(a[199] & b[190])^(a[198] & b[191])^(a[197] & b[192])^(a[196] & b[193])^(a[195] & b[194])^(a[194] & b[195])^(a[193] & b[196])^(a[192] & b[197])^(a[191] & b[198])^(a[190] & b[199])^(a[189] & b[200])^(a[188] & b[201])^(a[187] & b[202])^(a[186] & b[203])^(a[185] & b[204])^(a[184] & b[205])^(a[183] & b[206])^(a[182] & b[207])^(a[181] & b[208])^(a[180] & b[209])^(a[179] & b[210])^(a[178] & b[211])^(a[177] & b[212])^(a[176] & b[213])^(a[175] & b[214])^(a[174] & b[215])^(a[173] & b[216])^(a[172] & b[217])^(a[171] & b[218])^(a[170] & b[219])^(a[169] & b[220])^(a[168] & b[221])^(a[167] & b[222])^(a[166] & b[223])^(a[165] & b[224])^(a[164] & b[225])^(a[163] & b[226])^(a[162] & b[227])^(a[161] & b[228])^(a[160] & b[229])^(a[159] & b[230])^(a[158] & b[231])^(a[157] & b[232]);
assign y[390] = (a[232] & b[158])^(a[231] & b[159])^(a[230] & b[160])^(a[229] & b[161])^(a[228] & b[162])^(a[227] & b[163])^(a[226] & b[164])^(a[225] & b[165])^(a[224] & b[166])^(a[223] & b[167])^(a[222] & b[168])^(a[221] & b[169])^(a[220] & b[170])^(a[219] & b[171])^(a[218] & b[172])^(a[217] & b[173])^(a[216] & b[174])^(a[215] & b[175])^(a[214] & b[176])^(a[213] & b[177])^(a[212] & b[178])^(a[211] & b[179])^(a[210] & b[180])^(a[209] & b[181])^(a[208] & b[182])^(a[207] & b[183])^(a[206] & b[184])^(a[205] & b[185])^(a[204] & b[186])^(a[203] & b[187])^(a[202] & b[188])^(a[201] & b[189])^(a[200] & b[190])^(a[199] & b[191])^(a[198] & b[192])^(a[197] & b[193])^(a[196] & b[194])^(a[195] & b[195])^(a[194] & b[196])^(a[193] & b[197])^(a[192] & b[198])^(a[191] & b[199])^(a[190] & b[200])^(a[189] & b[201])^(a[188] & b[202])^(a[187] & b[203])^(a[186] & b[204])^(a[185] & b[205])^(a[184] & b[206])^(a[183] & b[207])^(a[182] & b[208])^(a[181] & b[209])^(a[180] & b[210])^(a[179] & b[211])^(a[178] & b[212])^(a[177] & b[213])^(a[176] & b[214])^(a[175] & b[215])^(a[174] & b[216])^(a[173] & b[217])^(a[172] & b[218])^(a[171] & b[219])^(a[170] & b[220])^(a[169] & b[221])^(a[168] & b[222])^(a[167] & b[223])^(a[166] & b[224])^(a[165] & b[225])^(a[164] & b[226])^(a[163] & b[227])^(a[162] & b[228])^(a[161] & b[229])^(a[160] & b[230])^(a[159] & b[231])^(a[158] & b[232]);
assign y[391] = (a[232] & b[159])^(a[231] & b[160])^(a[230] & b[161])^(a[229] & b[162])^(a[228] & b[163])^(a[227] & b[164])^(a[226] & b[165])^(a[225] & b[166])^(a[224] & b[167])^(a[223] & b[168])^(a[222] & b[169])^(a[221] & b[170])^(a[220] & b[171])^(a[219] & b[172])^(a[218] & b[173])^(a[217] & b[174])^(a[216] & b[175])^(a[215] & b[176])^(a[214] & b[177])^(a[213] & b[178])^(a[212] & b[179])^(a[211] & b[180])^(a[210] & b[181])^(a[209] & b[182])^(a[208] & b[183])^(a[207] & b[184])^(a[206] & b[185])^(a[205] & b[186])^(a[204] & b[187])^(a[203] & b[188])^(a[202] & b[189])^(a[201] & b[190])^(a[200] & b[191])^(a[199] & b[192])^(a[198] & b[193])^(a[197] & b[194])^(a[196] & b[195])^(a[195] & b[196])^(a[194] & b[197])^(a[193] & b[198])^(a[192] & b[199])^(a[191] & b[200])^(a[190] & b[201])^(a[189] & b[202])^(a[188] & b[203])^(a[187] & b[204])^(a[186] & b[205])^(a[185] & b[206])^(a[184] & b[207])^(a[183] & b[208])^(a[182] & b[209])^(a[181] & b[210])^(a[180] & b[211])^(a[179] & b[212])^(a[178] & b[213])^(a[177] & b[214])^(a[176] & b[215])^(a[175] & b[216])^(a[174] & b[217])^(a[173] & b[218])^(a[172] & b[219])^(a[171] & b[220])^(a[170] & b[221])^(a[169] & b[222])^(a[168] & b[223])^(a[167] & b[224])^(a[166] & b[225])^(a[165] & b[226])^(a[164] & b[227])^(a[163] & b[228])^(a[162] & b[229])^(a[161] & b[230])^(a[160] & b[231])^(a[159] & b[232]);
assign y[392] = (a[232] & b[160])^(a[231] & b[161])^(a[230] & b[162])^(a[229] & b[163])^(a[228] & b[164])^(a[227] & b[165])^(a[226] & b[166])^(a[225] & b[167])^(a[224] & b[168])^(a[223] & b[169])^(a[222] & b[170])^(a[221] & b[171])^(a[220] & b[172])^(a[219] & b[173])^(a[218] & b[174])^(a[217] & b[175])^(a[216] & b[176])^(a[215] & b[177])^(a[214] & b[178])^(a[213] & b[179])^(a[212] & b[180])^(a[211] & b[181])^(a[210] & b[182])^(a[209] & b[183])^(a[208] & b[184])^(a[207] & b[185])^(a[206] & b[186])^(a[205] & b[187])^(a[204] & b[188])^(a[203] & b[189])^(a[202] & b[190])^(a[201] & b[191])^(a[200] & b[192])^(a[199] & b[193])^(a[198] & b[194])^(a[197] & b[195])^(a[196] & b[196])^(a[195] & b[197])^(a[194] & b[198])^(a[193] & b[199])^(a[192] & b[200])^(a[191] & b[201])^(a[190] & b[202])^(a[189] & b[203])^(a[188] & b[204])^(a[187] & b[205])^(a[186] & b[206])^(a[185] & b[207])^(a[184] & b[208])^(a[183] & b[209])^(a[182] & b[210])^(a[181] & b[211])^(a[180] & b[212])^(a[179] & b[213])^(a[178] & b[214])^(a[177] & b[215])^(a[176] & b[216])^(a[175] & b[217])^(a[174] & b[218])^(a[173] & b[219])^(a[172] & b[220])^(a[171] & b[221])^(a[170] & b[222])^(a[169] & b[223])^(a[168] & b[224])^(a[167] & b[225])^(a[166] & b[226])^(a[165] & b[227])^(a[164] & b[228])^(a[163] & b[229])^(a[162] & b[230])^(a[161] & b[231])^(a[160] & b[232]);
assign y[393] = (a[232] & b[161])^(a[231] & b[162])^(a[230] & b[163])^(a[229] & b[164])^(a[228] & b[165])^(a[227] & b[166])^(a[226] & b[167])^(a[225] & b[168])^(a[224] & b[169])^(a[223] & b[170])^(a[222] & b[171])^(a[221] & b[172])^(a[220] & b[173])^(a[219] & b[174])^(a[218] & b[175])^(a[217] & b[176])^(a[216] & b[177])^(a[215] & b[178])^(a[214] & b[179])^(a[213] & b[180])^(a[212] & b[181])^(a[211] & b[182])^(a[210] & b[183])^(a[209] & b[184])^(a[208] & b[185])^(a[207] & b[186])^(a[206] & b[187])^(a[205] & b[188])^(a[204] & b[189])^(a[203] & b[190])^(a[202] & b[191])^(a[201] & b[192])^(a[200] & b[193])^(a[199] & b[194])^(a[198] & b[195])^(a[197] & b[196])^(a[196] & b[197])^(a[195] & b[198])^(a[194] & b[199])^(a[193] & b[200])^(a[192] & b[201])^(a[191] & b[202])^(a[190] & b[203])^(a[189] & b[204])^(a[188] & b[205])^(a[187] & b[206])^(a[186] & b[207])^(a[185] & b[208])^(a[184] & b[209])^(a[183] & b[210])^(a[182] & b[211])^(a[181] & b[212])^(a[180] & b[213])^(a[179] & b[214])^(a[178] & b[215])^(a[177] & b[216])^(a[176] & b[217])^(a[175] & b[218])^(a[174] & b[219])^(a[173] & b[220])^(a[172] & b[221])^(a[171] & b[222])^(a[170] & b[223])^(a[169] & b[224])^(a[168] & b[225])^(a[167] & b[226])^(a[166] & b[227])^(a[165] & b[228])^(a[164] & b[229])^(a[163] & b[230])^(a[162] & b[231])^(a[161] & b[232]);
assign y[394] = (a[232] & b[162])^(a[231] & b[163])^(a[230] & b[164])^(a[229] & b[165])^(a[228] & b[166])^(a[227] & b[167])^(a[226] & b[168])^(a[225] & b[169])^(a[224] & b[170])^(a[223] & b[171])^(a[222] & b[172])^(a[221] & b[173])^(a[220] & b[174])^(a[219] & b[175])^(a[218] & b[176])^(a[217] & b[177])^(a[216] & b[178])^(a[215] & b[179])^(a[214] & b[180])^(a[213] & b[181])^(a[212] & b[182])^(a[211] & b[183])^(a[210] & b[184])^(a[209] & b[185])^(a[208] & b[186])^(a[207] & b[187])^(a[206] & b[188])^(a[205] & b[189])^(a[204] & b[190])^(a[203] & b[191])^(a[202] & b[192])^(a[201] & b[193])^(a[200] & b[194])^(a[199] & b[195])^(a[198] & b[196])^(a[197] & b[197])^(a[196] & b[198])^(a[195] & b[199])^(a[194] & b[200])^(a[193] & b[201])^(a[192] & b[202])^(a[191] & b[203])^(a[190] & b[204])^(a[189] & b[205])^(a[188] & b[206])^(a[187] & b[207])^(a[186] & b[208])^(a[185] & b[209])^(a[184] & b[210])^(a[183] & b[211])^(a[182] & b[212])^(a[181] & b[213])^(a[180] & b[214])^(a[179] & b[215])^(a[178] & b[216])^(a[177] & b[217])^(a[176] & b[218])^(a[175] & b[219])^(a[174] & b[220])^(a[173] & b[221])^(a[172] & b[222])^(a[171] & b[223])^(a[170] & b[224])^(a[169] & b[225])^(a[168] & b[226])^(a[167] & b[227])^(a[166] & b[228])^(a[165] & b[229])^(a[164] & b[230])^(a[163] & b[231])^(a[162] & b[232]);
assign y[395] = (a[232] & b[163])^(a[231] & b[164])^(a[230] & b[165])^(a[229] & b[166])^(a[228] & b[167])^(a[227] & b[168])^(a[226] & b[169])^(a[225] & b[170])^(a[224] & b[171])^(a[223] & b[172])^(a[222] & b[173])^(a[221] & b[174])^(a[220] & b[175])^(a[219] & b[176])^(a[218] & b[177])^(a[217] & b[178])^(a[216] & b[179])^(a[215] & b[180])^(a[214] & b[181])^(a[213] & b[182])^(a[212] & b[183])^(a[211] & b[184])^(a[210] & b[185])^(a[209] & b[186])^(a[208] & b[187])^(a[207] & b[188])^(a[206] & b[189])^(a[205] & b[190])^(a[204] & b[191])^(a[203] & b[192])^(a[202] & b[193])^(a[201] & b[194])^(a[200] & b[195])^(a[199] & b[196])^(a[198] & b[197])^(a[197] & b[198])^(a[196] & b[199])^(a[195] & b[200])^(a[194] & b[201])^(a[193] & b[202])^(a[192] & b[203])^(a[191] & b[204])^(a[190] & b[205])^(a[189] & b[206])^(a[188] & b[207])^(a[187] & b[208])^(a[186] & b[209])^(a[185] & b[210])^(a[184] & b[211])^(a[183] & b[212])^(a[182] & b[213])^(a[181] & b[214])^(a[180] & b[215])^(a[179] & b[216])^(a[178] & b[217])^(a[177] & b[218])^(a[176] & b[219])^(a[175] & b[220])^(a[174] & b[221])^(a[173] & b[222])^(a[172] & b[223])^(a[171] & b[224])^(a[170] & b[225])^(a[169] & b[226])^(a[168] & b[227])^(a[167] & b[228])^(a[166] & b[229])^(a[165] & b[230])^(a[164] & b[231])^(a[163] & b[232]);
assign y[396] = (a[232] & b[164])^(a[231] & b[165])^(a[230] & b[166])^(a[229] & b[167])^(a[228] & b[168])^(a[227] & b[169])^(a[226] & b[170])^(a[225] & b[171])^(a[224] & b[172])^(a[223] & b[173])^(a[222] & b[174])^(a[221] & b[175])^(a[220] & b[176])^(a[219] & b[177])^(a[218] & b[178])^(a[217] & b[179])^(a[216] & b[180])^(a[215] & b[181])^(a[214] & b[182])^(a[213] & b[183])^(a[212] & b[184])^(a[211] & b[185])^(a[210] & b[186])^(a[209] & b[187])^(a[208] & b[188])^(a[207] & b[189])^(a[206] & b[190])^(a[205] & b[191])^(a[204] & b[192])^(a[203] & b[193])^(a[202] & b[194])^(a[201] & b[195])^(a[200] & b[196])^(a[199] & b[197])^(a[198] & b[198])^(a[197] & b[199])^(a[196] & b[200])^(a[195] & b[201])^(a[194] & b[202])^(a[193] & b[203])^(a[192] & b[204])^(a[191] & b[205])^(a[190] & b[206])^(a[189] & b[207])^(a[188] & b[208])^(a[187] & b[209])^(a[186] & b[210])^(a[185] & b[211])^(a[184] & b[212])^(a[183] & b[213])^(a[182] & b[214])^(a[181] & b[215])^(a[180] & b[216])^(a[179] & b[217])^(a[178] & b[218])^(a[177] & b[219])^(a[176] & b[220])^(a[175] & b[221])^(a[174] & b[222])^(a[173] & b[223])^(a[172] & b[224])^(a[171] & b[225])^(a[170] & b[226])^(a[169] & b[227])^(a[168] & b[228])^(a[167] & b[229])^(a[166] & b[230])^(a[165] & b[231])^(a[164] & b[232]);
assign y[397] = (a[232] & b[165])^(a[231] & b[166])^(a[230] & b[167])^(a[229] & b[168])^(a[228] & b[169])^(a[227] & b[170])^(a[226] & b[171])^(a[225] & b[172])^(a[224] & b[173])^(a[223] & b[174])^(a[222] & b[175])^(a[221] & b[176])^(a[220] & b[177])^(a[219] & b[178])^(a[218] & b[179])^(a[217] & b[180])^(a[216] & b[181])^(a[215] & b[182])^(a[214] & b[183])^(a[213] & b[184])^(a[212] & b[185])^(a[211] & b[186])^(a[210] & b[187])^(a[209] & b[188])^(a[208] & b[189])^(a[207] & b[190])^(a[206] & b[191])^(a[205] & b[192])^(a[204] & b[193])^(a[203] & b[194])^(a[202] & b[195])^(a[201] & b[196])^(a[200] & b[197])^(a[199] & b[198])^(a[198] & b[199])^(a[197] & b[200])^(a[196] & b[201])^(a[195] & b[202])^(a[194] & b[203])^(a[193] & b[204])^(a[192] & b[205])^(a[191] & b[206])^(a[190] & b[207])^(a[189] & b[208])^(a[188] & b[209])^(a[187] & b[210])^(a[186] & b[211])^(a[185] & b[212])^(a[184] & b[213])^(a[183] & b[214])^(a[182] & b[215])^(a[181] & b[216])^(a[180] & b[217])^(a[179] & b[218])^(a[178] & b[219])^(a[177] & b[220])^(a[176] & b[221])^(a[175] & b[222])^(a[174] & b[223])^(a[173] & b[224])^(a[172] & b[225])^(a[171] & b[226])^(a[170] & b[227])^(a[169] & b[228])^(a[168] & b[229])^(a[167] & b[230])^(a[166] & b[231])^(a[165] & b[232]);
assign y[398] = (a[232] & b[166])^(a[231] & b[167])^(a[230] & b[168])^(a[229] & b[169])^(a[228] & b[170])^(a[227] & b[171])^(a[226] & b[172])^(a[225] & b[173])^(a[224] & b[174])^(a[223] & b[175])^(a[222] & b[176])^(a[221] & b[177])^(a[220] & b[178])^(a[219] & b[179])^(a[218] & b[180])^(a[217] & b[181])^(a[216] & b[182])^(a[215] & b[183])^(a[214] & b[184])^(a[213] & b[185])^(a[212] & b[186])^(a[211] & b[187])^(a[210] & b[188])^(a[209] & b[189])^(a[208] & b[190])^(a[207] & b[191])^(a[206] & b[192])^(a[205] & b[193])^(a[204] & b[194])^(a[203] & b[195])^(a[202] & b[196])^(a[201] & b[197])^(a[200] & b[198])^(a[199] & b[199])^(a[198] & b[200])^(a[197] & b[201])^(a[196] & b[202])^(a[195] & b[203])^(a[194] & b[204])^(a[193] & b[205])^(a[192] & b[206])^(a[191] & b[207])^(a[190] & b[208])^(a[189] & b[209])^(a[188] & b[210])^(a[187] & b[211])^(a[186] & b[212])^(a[185] & b[213])^(a[184] & b[214])^(a[183] & b[215])^(a[182] & b[216])^(a[181] & b[217])^(a[180] & b[218])^(a[179] & b[219])^(a[178] & b[220])^(a[177] & b[221])^(a[176] & b[222])^(a[175] & b[223])^(a[174] & b[224])^(a[173] & b[225])^(a[172] & b[226])^(a[171] & b[227])^(a[170] & b[228])^(a[169] & b[229])^(a[168] & b[230])^(a[167] & b[231])^(a[166] & b[232]);
assign y[399] = (a[232] & b[167])^(a[231] & b[168])^(a[230] & b[169])^(a[229] & b[170])^(a[228] & b[171])^(a[227] & b[172])^(a[226] & b[173])^(a[225] & b[174])^(a[224] & b[175])^(a[223] & b[176])^(a[222] & b[177])^(a[221] & b[178])^(a[220] & b[179])^(a[219] & b[180])^(a[218] & b[181])^(a[217] & b[182])^(a[216] & b[183])^(a[215] & b[184])^(a[214] & b[185])^(a[213] & b[186])^(a[212] & b[187])^(a[211] & b[188])^(a[210] & b[189])^(a[209] & b[190])^(a[208] & b[191])^(a[207] & b[192])^(a[206] & b[193])^(a[205] & b[194])^(a[204] & b[195])^(a[203] & b[196])^(a[202] & b[197])^(a[201] & b[198])^(a[200] & b[199])^(a[199] & b[200])^(a[198] & b[201])^(a[197] & b[202])^(a[196] & b[203])^(a[195] & b[204])^(a[194] & b[205])^(a[193] & b[206])^(a[192] & b[207])^(a[191] & b[208])^(a[190] & b[209])^(a[189] & b[210])^(a[188] & b[211])^(a[187] & b[212])^(a[186] & b[213])^(a[185] & b[214])^(a[184] & b[215])^(a[183] & b[216])^(a[182] & b[217])^(a[181] & b[218])^(a[180] & b[219])^(a[179] & b[220])^(a[178] & b[221])^(a[177] & b[222])^(a[176] & b[223])^(a[175] & b[224])^(a[174] & b[225])^(a[173] & b[226])^(a[172] & b[227])^(a[171] & b[228])^(a[170] & b[229])^(a[169] & b[230])^(a[168] & b[231])^(a[167] & b[232]);
assign y[400] = (a[232] & b[168])^(a[231] & b[169])^(a[230] & b[170])^(a[229] & b[171])^(a[228] & b[172])^(a[227] & b[173])^(a[226] & b[174])^(a[225] & b[175])^(a[224] & b[176])^(a[223] & b[177])^(a[222] & b[178])^(a[221] & b[179])^(a[220] & b[180])^(a[219] & b[181])^(a[218] & b[182])^(a[217] & b[183])^(a[216] & b[184])^(a[215] & b[185])^(a[214] & b[186])^(a[213] & b[187])^(a[212] & b[188])^(a[211] & b[189])^(a[210] & b[190])^(a[209] & b[191])^(a[208] & b[192])^(a[207] & b[193])^(a[206] & b[194])^(a[205] & b[195])^(a[204] & b[196])^(a[203] & b[197])^(a[202] & b[198])^(a[201] & b[199])^(a[200] & b[200])^(a[199] & b[201])^(a[198] & b[202])^(a[197] & b[203])^(a[196] & b[204])^(a[195] & b[205])^(a[194] & b[206])^(a[193] & b[207])^(a[192] & b[208])^(a[191] & b[209])^(a[190] & b[210])^(a[189] & b[211])^(a[188] & b[212])^(a[187] & b[213])^(a[186] & b[214])^(a[185] & b[215])^(a[184] & b[216])^(a[183] & b[217])^(a[182] & b[218])^(a[181] & b[219])^(a[180] & b[220])^(a[179] & b[221])^(a[178] & b[222])^(a[177] & b[223])^(a[176] & b[224])^(a[175] & b[225])^(a[174] & b[226])^(a[173] & b[227])^(a[172] & b[228])^(a[171] & b[229])^(a[170] & b[230])^(a[169] & b[231])^(a[168] & b[232]);
assign y[401] = (a[232] & b[169])^(a[231] & b[170])^(a[230] & b[171])^(a[229] & b[172])^(a[228] & b[173])^(a[227] & b[174])^(a[226] & b[175])^(a[225] & b[176])^(a[224] & b[177])^(a[223] & b[178])^(a[222] & b[179])^(a[221] & b[180])^(a[220] & b[181])^(a[219] & b[182])^(a[218] & b[183])^(a[217] & b[184])^(a[216] & b[185])^(a[215] & b[186])^(a[214] & b[187])^(a[213] & b[188])^(a[212] & b[189])^(a[211] & b[190])^(a[210] & b[191])^(a[209] & b[192])^(a[208] & b[193])^(a[207] & b[194])^(a[206] & b[195])^(a[205] & b[196])^(a[204] & b[197])^(a[203] & b[198])^(a[202] & b[199])^(a[201] & b[200])^(a[200] & b[201])^(a[199] & b[202])^(a[198] & b[203])^(a[197] & b[204])^(a[196] & b[205])^(a[195] & b[206])^(a[194] & b[207])^(a[193] & b[208])^(a[192] & b[209])^(a[191] & b[210])^(a[190] & b[211])^(a[189] & b[212])^(a[188] & b[213])^(a[187] & b[214])^(a[186] & b[215])^(a[185] & b[216])^(a[184] & b[217])^(a[183] & b[218])^(a[182] & b[219])^(a[181] & b[220])^(a[180] & b[221])^(a[179] & b[222])^(a[178] & b[223])^(a[177] & b[224])^(a[176] & b[225])^(a[175] & b[226])^(a[174] & b[227])^(a[173] & b[228])^(a[172] & b[229])^(a[171] & b[230])^(a[170] & b[231])^(a[169] & b[232]);
assign y[402] = (a[232] & b[170])^(a[231] & b[171])^(a[230] & b[172])^(a[229] & b[173])^(a[228] & b[174])^(a[227] & b[175])^(a[226] & b[176])^(a[225] & b[177])^(a[224] & b[178])^(a[223] & b[179])^(a[222] & b[180])^(a[221] & b[181])^(a[220] & b[182])^(a[219] & b[183])^(a[218] & b[184])^(a[217] & b[185])^(a[216] & b[186])^(a[215] & b[187])^(a[214] & b[188])^(a[213] & b[189])^(a[212] & b[190])^(a[211] & b[191])^(a[210] & b[192])^(a[209] & b[193])^(a[208] & b[194])^(a[207] & b[195])^(a[206] & b[196])^(a[205] & b[197])^(a[204] & b[198])^(a[203] & b[199])^(a[202] & b[200])^(a[201] & b[201])^(a[200] & b[202])^(a[199] & b[203])^(a[198] & b[204])^(a[197] & b[205])^(a[196] & b[206])^(a[195] & b[207])^(a[194] & b[208])^(a[193] & b[209])^(a[192] & b[210])^(a[191] & b[211])^(a[190] & b[212])^(a[189] & b[213])^(a[188] & b[214])^(a[187] & b[215])^(a[186] & b[216])^(a[185] & b[217])^(a[184] & b[218])^(a[183] & b[219])^(a[182] & b[220])^(a[181] & b[221])^(a[180] & b[222])^(a[179] & b[223])^(a[178] & b[224])^(a[177] & b[225])^(a[176] & b[226])^(a[175] & b[227])^(a[174] & b[228])^(a[173] & b[229])^(a[172] & b[230])^(a[171] & b[231])^(a[170] & b[232]);
assign y[403] = (a[232] & b[171])^(a[231] & b[172])^(a[230] & b[173])^(a[229] & b[174])^(a[228] & b[175])^(a[227] & b[176])^(a[226] & b[177])^(a[225] & b[178])^(a[224] & b[179])^(a[223] & b[180])^(a[222] & b[181])^(a[221] & b[182])^(a[220] & b[183])^(a[219] & b[184])^(a[218] & b[185])^(a[217] & b[186])^(a[216] & b[187])^(a[215] & b[188])^(a[214] & b[189])^(a[213] & b[190])^(a[212] & b[191])^(a[211] & b[192])^(a[210] & b[193])^(a[209] & b[194])^(a[208] & b[195])^(a[207] & b[196])^(a[206] & b[197])^(a[205] & b[198])^(a[204] & b[199])^(a[203] & b[200])^(a[202] & b[201])^(a[201] & b[202])^(a[200] & b[203])^(a[199] & b[204])^(a[198] & b[205])^(a[197] & b[206])^(a[196] & b[207])^(a[195] & b[208])^(a[194] & b[209])^(a[193] & b[210])^(a[192] & b[211])^(a[191] & b[212])^(a[190] & b[213])^(a[189] & b[214])^(a[188] & b[215])^(a[187] & b[216])^(a[186] & b[217])^(a[185] & b[218])^(a[184] & b[219])^(a[183] & b[220])^(a[182] & b[221])^(a[181] & b[222])^(a[180] & b[223])^(a[179] & b[224])^(a[178] & b[225])^(a[177] & b[226])^(a[176] & b[227])^(a[175] & b[228])^(a[174] & b[229])^(a[173] & b[230])^(a[172] & b[231])^(a[171] & b[232]);
assign y[404] = (a[232] & b[172])^(a[231] & b[173])^(a[230] & b[174])^(a[229] & b[175])^(a[228] & b[176])^(a[227] & b[177])^(a[226] & b[178])^(a[225] & b[179])^(a[224] & b[180])^(a[223] & b[181])^(a[222] & b[182])^(a[221] & b[183])^(a[220] & b[184])^(a[219] & b[185])^(a[218] & b[186])^(a[217] & b[187])^(a[216] & b[188])^(a[215] & b[189])^(a[214] & b[190])^(a[213] & b[191])^(a[212] & b[192])^(a[211] & b[193])^(a[210] & b[194])^(a[209] & b[195])^(a[208] & b[196])^(a[207] & b[197])^(a[206] & b[198])^(a[205] & b[199])^(a[204] & b[200])^(a[203] & b[201])^(a[202] & b[202])^(a[201] & b[203])^(a[200] & b[204])^(a[199] & b[205])^(a[198] & b[206])^(a[197] & b[207])^(a[196] & b[208])^(a[195] & b[209])^(a[194] & b[210])^(a[193] & b[211])^(a[192] & b[212])^(a[191] & b[213])^(a[190] & b[214])^(a[189] & b[215])^(a[188] & b[216])^(a[187] & b[217])^(a[186] & b[218])^(a[185] & b[219])^(a[184] & b[220])^(a[183] & b[221])^(a[182] & b[222])^(a[181] & b[223])^(a[180] & b[224])^(a[179] & b[225])^(a[178] & b[226])^(a[177] & b[227])^(a[176] & b[228])^(a[175] & b[229])^(a[174] & b[230])^(a[173] & b[231])^(a[172] & b[232]);
assign y[405] = (a[232] & b[173])^(a[231] & b[174])^(a[230] & b[175])^(a[229] & b[176])^(a[228] & b[177])^(a[227] & b[178])^(a[226] & b[179])^(a[225] & b[180])^(a[224] & b[181])^(a[223] & b[182])^(a[222] & b[183])^(a[221] & b[184])^(a[220] & b[185])^(a[219] & b[186])^(a[218] & b[187])^(a[217] & b[188])^(a[216] & b[189])^(a[215] & b[190])^(a[214] & b[191])^(a[213] & b[192])^(a[212] & b[193])^(a[211] & b[194])^(a[210] & b[195])^(a[209] & b[196])^(a[208] & b[197])^(a[207] & b[198])^(a[206] & b[199])^(a[205] & b[200])^(a[204] & b[201])^(a[203] & b[202])^(a[202] & b[203])^(a[201] & b[204])^(a[200] & b[205])^(a[199] & b[206])^(a[198] & b[207])^(a[197] & b[208])^(a[196] & b[209])^(a[195] & b[210])^(a[194] & b[211])^(a[193] & b[212])^(a[192] & b[213])^(a[191] & b[214])^(a[190] & b[215])^(a[189] & b[216])^(a[188] & b[217])^(a[187] & b[218])^(a[186] & b[219])^(a[185] & b[220])^(a[184] & b[221])^(a[183] & b[222])^(a[182] & b[223])^(a[181] & b[224])^(a[180] & b[225])^(a[179] & b[226])^(a[178] & b[227])^(a[177] & b[228])^(a[176] & b[229])^(a[175] & b[230])^(a[174] & b[231])^(a[173] & b[232]);
assign y[406] = (a[232] & b[174])^(a[231] & b[175])^(a[230] & b[176])^(a[229] & b[177])^(a[228] & b[178])^(a[227] & b[179])^(a[226] & b[180])^(a[225] & b[181])^(a[224] & b[182])^(a[223] & b[183])^(a[222] & b[184])^(a[221] & b[185])^(a[220] & b[186])^(a[219] & b[187])^(a[218] & b[188])^(a[217] & b[189])^(a[216] & b[190])^(a[215] & b[191])^(a[214] & b[192])^(a[213] & b[193])^(a[212] & b[194])^(a[211] & b[195])^(a[210] & b[196])^(a[209] & b[197])^(a[208] & b[198])^(a[207] & b[199])^(a[206] & b[200])^(a[205] & b[201])^(a[204] & b[202])^(a[203] & b[203])^(a[202] & b[204])^(a[201] & b[205])^(a[200] & b[206])^(a[199] & b[207])^(a[198] & b[208])^(a[197] & b[209])^(a[196] & b[210])^(a[195] & b[211])^(a[194] & b[212])^(a[193] & b[213])^(a[192] & b[214])^(a[191] & b[215])^(a[190] & b[216])^(a[189] & b[217])^(a[188] & b[218])^(a[187] & b[219])^(a[186] & b[220])^(a[185] & b[221])^(a[184] & b[222])^(a[183] & b[223])^(a[182] & b[224])^(a[181] & b[225])^(a[180] & b[226])^(a[179] & b[227])^(a[178] & b[228])^(a[177] & b[229])^(a[176] & b[230])^(a[175] & b[231])^(a[174] & b[232]);
assign y[407] = (a[232] & b[175])^(a[231] & b[176])^(a[230] & b[177])^(a[229] & b[178])^(a[228] & b[179])^(a[227] & b[180])^(a[226] & b[181])^(a[225] & b[182])^(a[224] & b[183])^(a[223] & b[184])^(a[222] & b[185])^(a[221] & b[186])^(a[220] & b[187])^(a[219] & b[188])^(a[218] & b[189])^(a[217] & b[190])^(a[216] & b[191])^(a[215] & b[192])^(a[214] & b[193])^(a[213] & b[194])^(a[212] & b[195])^(a[211] & b[196])^(a[210] & b[197])^(a[209] & b[198])^(a[208] & b[199])^(a[207] & b[200])^(a[206] & b[201])^(a[205] & b[202])^(a[204] & b[203])^(a[203] & b[204])^(a[202] & b[205])^(a[201] & b[206])^(a[200] & b[207])^(a[199] & b[208])^(a[198] & b[209])^(a[197] & b[210])^(a[196] & b[211])^(a[195] & b[212])^(a[194] & b[213])^(a[193] & b[214])^(a[192] & b[215])^(a[191] & b[216])^(a[190] & b[217])^(a[189] & b[218])^(a[188] & b[219])^(a[187] & b[220])^(a[186] & b[221])^(a[185] & b[222])^(a[184] & b[223])^(a[183] & b[224])^(a[182] & b[225])^(a[181] & b[226])^(a[180] & b[227])^(a[179] & b[228])^(a[178] & b[229])^(a[177] & b[230])^(a[176] & b[231])^(a[175] & b[232]);
assign y[408] = (a[232] & b[176])^(a[231] & b[177])^(a[230] & b[178])^(a[229] & b[179])^(a[228] & b[180])^(a[227] & b[181])^(a[226] & b[182])^(a[225] & b[183])^(a[224] & b[184])^(a[223] & b[185])^(a[222] & b[186])^(a[221] & b[187])^(a[220] & b[188])^(a[219] & b[189])^(a[218] & b[190])^(a[217] & b[191])^(a[216] & b[192])^(a[215] & b[193])^(a[214] & b[194])^(a[213] & b[195])^(a[212] & b[196])^(a[211] & b[197])^(a[210] & b[198])^(a[209] & b[199])^(a[208] & b[200])^(a[207] & b[201])^(a[206] & b[202])^(a[205] & b[203])^(a[204] & b[204])^(a[203] & b[205])^(a[202] & b[206])^(a[201] & b[207])^(a[200] & b[208])^(a[199] & b[209])^(a[198] & b[210])^(a[197] & b[211])^(a[196] & b[212])^(a[195] & b[213])^(a[194] & b[214])^(a[193] & b[215])^(a[192] & b[216])^(a[191] & b[217])^(a[190] & b[218])^(a[189] & b[219])^(a[188] & b[220])^(a[187] & b[221])^(a[186] & b[222])^(a[185] & b[223])^(a[184] & b[224])^(a[183] & b[225])^(a[182] & b[226])^(a[181] & b[227])^(a[180] & b[228])^(a[179] & b[229])^(a[178] & b[230])^(a[177] & b[231])^(a[176] & b[232]);
assign y[409] = (a[232] & b[177])^(a[231] & b[178])^(a[230] & b[179])^(a[229] & b[180])^(a[228] & b[181])^(a[227] & b[182])^(a[226] & b[183])^(a[225] & b[184])^(a[224] & b[185])^(a[223] & b[186])^(a[222] & b[187])^(a[221] & b[188])^(a[220] & b[189])^(a[219] & b[190])^(a[218] & b[191])^(a[217] & b[192])^(a[216] & b[193])^(a[215] & b[194])^(a[214] & b[195])^(a[213] & b[196])^(a[212] & b[197])^(a[211] & b[198])^(a[210] & b[199])^(a[209] & b[200])^(a[208] & b[201])^(a[207] & b[202])^(a[206] & b[203])^(a[205] & b[204])^(a[204] & b[205])^(a[203] & b[206])^(a[202] & b[207])^(a[201] & b[208])^(a[200] & b[209])^(a[199] & b[210])^(a[198] & b[211])^(a[197] & b[212])^(a[196] & b[213])^(a[195] & b[214])^(a[194] & b[215])^(a[193] & b[216])^(a[192] & b[217])^(a[191] & b[218])^(a[190] & b[219])^(a[189] & b[220])^(a[188] & b[221])^(a[187] & b[222])^(a[186] & b[223])^(a[185] & b[224])^(a[184] & b[225])^(a[183] & b[226])^(a[182] & b[227])^(a[181] & b[228])^(a[180] & b[229])^(a[179] & b[230])^(a[178] & b[231])^(a[177] & b[232]);
assign y[410] = (a[232] & b[178])^(a[231] & b[179])^(a[230] & b[180])^(a[229] & b[181])^(a[228] & b[182])^(a[227] & b[183])^(a[226] & b[184])^(a[225] & b[185])^(a[224] & b[186])^(a[223] & b[187])^(a[222] & b[188])^(a[221] & b[189])^(a[220] & b[190])^(a[219] & b[191])^(a[218] & b[192])^(a[217] & b[193])^(a[216] & b[194])^(a[215] & b[195])^(a[214] & b[196])^(a[213] & b[197])^(a[212] & b[198])^(a[211] & b[199])^(a[210] & b[200])^(a[209] & b[201])^(a[208] & b[202])^(a[207] & b[203])^(a[206] & b[204])^(a[205] & b[205])^(a[204] & b[206])^(a[203] & b[207])^(a[202] & b[208])^(a[201] & b[209])^(a[200] & b[210])^(a[199] & b[211])^(a[198] & b[212])^(a[197] & b[213])^(a[196] & b[214])^(a[195] & b[215])^(a[194] & b[216])^(a[193] & b[217])^(a[192] & b[218])^(a[191] & b[219])^(a[190] & b[220])^(a[189] & b[221])^(a[188] & b[222])^(a[187] & b[223])^(a[186] & b[224])^(a[185] & b[225])^(a[184] & b[226])^(a[183] & b[227])^(a[182] & b[228])^(a[181] & b[229])^(a[180] & b[230])^(a[179] & b[231])^(a[178] & b[232]);
assign y[411] = (a[232] & b[179])^(a[231] & b[180])^(a[230] & b[181])^(a[229] & b[182])^(a[228] & b[183])^(a[227] & b[184])^(a[226] & b[185])^(a[225] & b[186])^(a[224] & b[187])^(a[223] & b[188])^(a[222] & b[189])^(a[221] & b[190])^(a[220] & b[191])^(a[219] & b[192])^(a[218] & b[193])^(a[217] & b[194])^(a[216] & b[195])^(a[215] & b[196])^(a[214] & b[197])^(a[213] & b[198])^(a[212] & b[199])^(a[211] & b[200])^(a[210] & b[201])^(a[209] & b[202])^(a[208] & b[203])^(a[207] & b[204])^(a[206] & b[205])^(a[205] & b[206])^(a[204] & b[207])^(a[203] & b[208])^(a[202] & b[209])^(a[201] & b[210])^(a[200] & b[211])^(a[199] & b[212])^(a[198] & b[213])^(a[197] & b[214])^(a[196] & b[215])^(a[195] & b[216])^(a[194] & b[217])^(a[193] & b[218])^(a[192] & b[219])^(a[191] & b[220])^(a[190] & b[221])^(a[189] & b[222])^(a[188] & b[223])^(a[187] & b[224])^(a[186] & b[225])^(a[185] & b[226])^(a[184] & b[227])^(a[183] & b[228])^(a[182] & b[229])^(a[181] & b[230])^(a[180] & b[231])^(a[179] & b[232]);
assign y[412] = (a[232] & b[180])^(a[231] & b[181])^(a[230] & b[182])^(a[229] & b[183])^(a[228] & b[184])^(a[227] & b[185])^(a[226] & b[186])^(a[225] & b[187])^(a[224] & b[188])^(a[223] & b[189])^(a[222] & b[190])^(a[221] & b[191])^(a[220] & b[192])^(a[219] & b[193])^(a[218] & b[194])^(a[217] & b[195])^(a[216] & b[196])^(a[215] & b[197])^(a[214] & b[198])^(a[213] & b[199])^(a[212] & b[200])^(a[211] & b[201])^(a[210] & b[202])^(a[209] & b[203])^(a[208] & b[204])^(a[207] & b[205])^(a[206] & b[206])^(a[205] & b[207])^(a[204] & b[208])^(a[203] & b[209])^(a[202] & b[210])^(a[201] & b[211])^(a[200] & b[212])^(a[199] & b[213])^(a[198] & b[214])^(a[197] & b[215])^(a[196] & b[216])^(a[195] & b[217])^(a[194] & b[218])^(a[193] & b[219])^(a[192] & b[220])^(a[191] & b[221])^(a[190] & b[222])^(a[189] & b[223])^(a[188] & b[224])^(a[187] & b[225])^(a[186] & b[226])^(a[185] & b[227])^(a[184] & b[228])^(a[183] & b[229])^(a[182] & b[230])^(a[181] & b[231])^(a[180] & b[232]);
assign y[413] = (a[232] & b[181])^(a[231] & b[182])^(a[230] & b[183])^(a[229] & b[184])^(a[228] & b[185])^(a[227] & b[186])^(a[226] & b[187])^(a[225] & b[188])^(a[224] & b[189])^(a[223] & b[190])^(a[222] & b[191])^(a[221] & b[192])^(a[220] & b[193])^(a[219] & b[194])^(a[218] & b[195])^(a[217] & b[196])^(a[216] & b[197])^(a[215] & b[198])^(a[214] & b[199])^(a[213] & b[200])^(a[212] & b[201])^(a[211] & b[202])^(a[210] & b[203])^(a[209] & b[204])^(a[208] & b[205])^(a[207] & b[206])^(a[206] & b[207])^(a[205] & b[208])^(a[204] & b[209])^(a[203] & b[210])^(a[202] & b[211])^(a[201] & b[212])^(a[200] & b[213])^(a[199] & b[214])^(a[198] & b[215])^(a[197] & b[216])^(a[196] & b[217])^(a[195] & b[218])^(a[194] & b[219])^(a[193] & b[220])^(a[192] & b[221])^(a[191] & b[222])^(a[190] & b[223])^(a[189] & b[224])^(a[188] & b[225])^(a[187] & b[226])^(a[186] & b[227])^(a[185] & b[228])^(a[184] & b[229])^(a[183] & b[230])^(a[182] & b[231])^(a[181] & b[232]);
assign y[414] = (a[232] & b[182])^(a[231] & b[183])^(a[230] & b[184])^(a[229] & b[185])^(a[228] & b[186])^(a[227] & b[187])^(a[226] & b[188])^(a[225] & b[189])^(a[224] & b[190])^(a[223] & b[191])^(a[222] & b[192])^(a[221] & b[193])^(a[220] & b[194])^(a[219] & b[195])^(a[218] & b[196])^(a[217] & b[197])^(a[216] & b[198])^(a[215] & b[199])^(a[214] & b[200])^(a[213] & b[201])^(a[212] & b[202])^(a[211] & b[203])^(a[210] & b[204])^(a[209] & b[205])^(a[208] & b[206])^(a[207] & b[207])^(a[206] & b[208])^(a[205] & b[209])^(a[204] & b[210])^(a[203] & b[211])^(a[202] & b[212])^(a[201] & b[213])^(a[200] & b[214])^(a[199] & b[215])^(a[198] & b[216])^(a[197] & b[217])^(a[196] & b[218])^(a[195] & b[219])^(a[194] & b[220])^(a[193] & b[221])^(a[192] & b[222])^(a[191] & b[223])^(a[190] & b[224])^(a[189] & b[225])^(a[188] & b[226])^(a[187] & b[227])^(a[186] & b[228])^(a[185] & b[229])^(a[184] & b[230])^(a[183] & b[231])^(a[182] & b[232]);
assign y[415] = (a[232] & b[183])^(a[231] & b[184])^(a[230] & b[185])^(a[229] & b[186])^(a[228] & b[187])^(a[227] & b[188])^(a[226] & b[189])^(a[225] & b[190])^(a[224] & b[191])^(a[223] & b[192])^(a[222] & b[193])^(a[221] & b[194])^(a[220] & b[195])^(a[219] & b[196])^(a[218] & b[197])^(a[217] & b[198])^(a[216] & b[199])^(a[215] & b[200])^(a[214] & b[201])^(a[213] & b[202])^(a[212] & b[203])^(a[211] & b[204])^(a[210] & b[205])^(a[209] & b[206])^(a[208] & b[207])^(a[207] & b[208])^(a[206] & b[209])^(a[205] & b[210])^(a[204] & b[211])^(a[203] & b[212])^(a[202] & b[213])^(a[201] & b[214])^(a[200] & b[215])^(a[199] & b[216])^(a[198] & b[217])^(a[197] & b[218])^(a[196] & b[219])^(a[195] & b[220])^(a[194] & b[221])^(a[193] & b[222])^(a[192] & b[223])^(a[191] & b[224])^(a[190] & b[225])^(a[189] & b[226])^(a[188] & b[227])^(a[187] & b[228])^(a[186] & b[229])^(a[185] & b[230])^(a[184] & b[231])^(a[183] & b[232]);
assign y[416] = (a[232] & b[184])^(a[231] & b[185])^(a[230] & b[186])^(a[229] & b[187])^(a[228] & b[188])^(a[227] & b[189])^(a[226] & b[190])^(a[225] & b[191])^(a[224] & b[192])^(a[223] & b[193])^(a[222] & b[194])^(a[221] & b[195])^(a[220] & b[196])^(a[219] & b[197])^(a[218] & b[198])^(a[217] & b[199])^(a[216] & b[200])^(a[215] & b[201])^(a[214] & b[202])^(a[213] & b[203])^(a[212] & b[204])^(a[211] & b[205])^(a[210] & b[206])^(a[209] & b[207])^(a[208] & b[208])^(a[207] & b[209])^(a[206] & b[210])^(a[205] & b[211])^(a[204] & b[212])^(a[203] & b[213])^(a[202] & b[214])^(a[201] & b[215])^(a[200] & b[216])^(a[199] & b[217])^(a[198] & b[218])^(a[197] & b[219])^(a[196] & b[220])^(a[195] & b[221])^(a[194] & b[222])^(a[193] & b[223])^(a[192] & b[224])^(a[191] & b[225])^(a[190] & b[226])^(a[189] & b[227])^(a[188] & b[228])^(a[187] & b[229])^(a[186] & b[230])^(a[185] & b[231])^(a[184] & b[232]);
assign y[417] = (a[232] & b[185])^(a[231] & b[186])^(a[230] & b[187])^(a[229] & b[188])^(a[228] & b[189])^(a[227] & b[190])^(a[226] & b[191])^(a[225] & b[192])^(a[224] & b[193])^(a[223] & b[194])^(a[222] & b[195])^(a[221] & b[196])^(a[220] & b[197])^(a[219] & b[198])^(a[218] & b[199])^(a[217] & b[200])^(a[216] & b[201])^(a[215] & b[202])^(a[214] & b[203])^(a[213] & b[204])^(a[212] & b[205])^(a[211] & b[206])^(a[210] & b[207])^(a[209] & b[208])^(a[208] & b[209])^(a[207] & b[210])^(a[206] & b[211])^(a[205] & b[212])^(a[204] & b[213])^(a[203] & b[214])^(a[202] & b[215])^(a[201] & b[216])^(a[200] & b[217])^(a[199] & b[218])^(a[198] & b[219])^(a[197] & b[220])^(a[196] & b[221])^(a[195] & b[222])^(a[194] & b[223])^(a[193] & b[224])^(a[192] & b[225])^(a[191] & b[226])^(a[190] & b[227])^(a[189] & b[228])^(a[188] & b[229])^(a[187] & b[230])^(a[186] & b[231])^(a[185] & b[232]);
assign y[418] = (a[232] & b[186])^(a[231] & b[187])^(a[230] & b[188])^(a[229] & b[189])^(a[228] & b[190])^(a[227] & b[191])^(a[226] & b[192])^(a[225] & b[193])^(a[224] & b[194])^(a[223] & b[195])^(a[222] & b[196])^(a[221] & b[197])^(a[220] & b[198])^(a[219] & b[199])^(a[218] & b[200])^(a[217] & b[201])^(a[216] & b[202])^(a[215] & b[203])^(a[214] & b[204])^(a[213] & b[205])^(a[212] & b[206])^(a[211] & b[207])^(a[210] & b[208])^(a[209] & b[209])^(a[208] & b[210])^(a[207] & b[211])^(a[206] & b[212])^(a[205] & b[213])^(a[204] & b[214])^(a[203] & b[215])^(a[202] & b[216])^(a[201] & b[217])^(a[200] & b[218])^(a[199] & b[219])^(a[198] & b[220])^(a[197] & b[221])^(a[196] & b[222])^(a[195] & b[223])^(a[194] & b[224])^(a[193] & b[225])^(a[192] & b[226])^(a[191] & b[227])^(a[190] & b[228])^(a[189] & b[229])^(a[188] & b[230])^(a[187] & b[231])^(a[186] & b[232]);
assign y[419] = (a[232] & b[187])^(a[231] & b[188])^(a[230] & b[189])^(a[229] & b[190])^(a[228] & b[191])^(a[227] & b[192])^(a[226] & b[193])^(a[225] & b[194])^(a[224] & b[195])^(a[223] & b[196])^(a[222] & b[197])^(a[221] & b[198])^(a[220] & b[199])^(a[219] & b[200])^(a[218] & b[201])^(a[217] & b[202])^(a[216] & b[203])^(a[215] & b[204])^(a[214] & b[205])^(a[213] & b[206])^(a[212] & b[207])^(a[211] & b[208])^(a[210] & b[209])^(a[209] & b[210])^(a[208] & b[211])^(a[207] & b[212])^(a[206] & b[213])^(a[205] & b[214])^(a[204] & b[215])^(a[203] & b[216])^(a[202] & b[217])^(a[201] & b[218])^(a[200] & b[219])^(a[199] & b[220])^(a[198] & b[221])^(a[197] & b[222])^(a[196] & b[223])^(a[195] & b[224])^(a[194] & b[225])^(a[193] & b[226])^(a[192] & b[227])^(a[191] & b[228])^(a[190] & b[229])^(a[189] & b[230])^(a[188] & b[231])^(a[187] & b[232]);
assign y[420] = (a[232] & b[188])^(a[231] & b[189])^(a[230] & b[190])^(a[229] & b[191])^(a[228] & b[192])^(a[227] & b[193])^(a[226] & b[194])^(a[225] & b[195])^(a[224] & b[196])^(a[223] & b[197])^(a[222] & b[198])^(a[221] & b[199])^(a[220] & b[200])^(a[219] & b[201])^(a[218] & b[202])^(a[217] & b[203])^(a[216] & b[204])^(a[215] & b[205])^(a[214] & b[206])^(a[213] & b[207])^(a[212] & b[208])^(a[211] & b[209])^(a[210] & b[210])^(a[209] & b[211])^(a[208] & b[212])^(a[207] & b[213])^(a[206] & b[214])^(a[205] & b[215])^(a[204] & b[216])^(a[203] & b[217])^(a[202] & b[218])^(a[201] & b[219])^(a[200] & b[220])^(a[199] & b[221])^(a[198] & b[222])^(a[197] & b[223])^(a[196] & b[224])^(a[195] & b[225])^(a[194] & b[226])^(a[193] & b[227])^(a[192] & b[228])^(a[191] & b[229])^(a[190] & b[230])^(a[189] & b[231])^(a[188] & b[232]);
assign y[421] = (a[232] & b[189])^(a[231] & b[190])^(a[230] & b[191])^(a[229] & b[192])^(a[228] & b[193])^(a[227] & b[194])^(a[226] & b[195])^(a[225] & b[196])^(a[224] & b[197])^(a[223] & b[198])^(a[222] & b[199])^(a[221] & b[200])^(a[220] & b[201])^(a[219] & b[202])^(a[218] & b[203])^(a[217] & b[204])^(a[216] & b[205])^(a[215] & b[206])^(a[214] & b[207])^(a[213] & b[208])^(a[212] & b[209])^(a[211] & b[210])^(a[210] & b[211])^(a[209] & b[212])^(a[208] & b[213])^(a[207] & b[214])^(a[206] & b[215])^(a[205] & b[216])^(a[204] & b[217])^(a[203] & b[218])^(a[202] & b[219])^(a[201] & b[220])^(a[200] & b[221])^(a[199] & b[222])^(a[198] & b[223])^(a[197] & b[224])^(a[196] & b[225])^(a[195] & b[226])^(a[194] & b[227])^(a[193] & b[228])^(a[192] & b[229])^(a[191] & b[230])^(a[190] & b[231])^(a[189] & b[232]);
assign y[422] = (a[232] & b[190])^(a[231] & b[191])^(a[230] & b[192])^(a[229] & b[193])^(a[228] & b[194])^(a[227] & b[195])^(a[226] & b[196])^(a[225] & b[197])^(a[224] & b[198])^(a[223] & b[199])^(a[222] & b[200])^(a[221] & b[201])^(a[220] & b[202])^(a[219] & b[203])^(a[218] & b[204])^(a[217] & b[205])^(a[216] & b[206])^(a[215] & b[207])^(a[214] & b[208])^(a[213] & b[209])^(a[212] & b[210])^(a[211] & b[211])^(a[210] & b[212])^(a[209] & b[213])^(a[208] & b[214])^(a[207] & b[215])^(a[206] & b[216])^(a[205] & b[217])^(a[204] & b[218])^(a[203] & b[219])^(a[202] & b[220])^(a[201] & b[221])^(a[200] & b[222])^(a[199] & b[223])^(a[198] & b[224])^(a[197] & b[225])^(a[196] & b[226])^(a[195] & b[227])^(a[194] & b[228])^(a[193] & b[229])^(a[192] & b[230])^(a[191] & b[231])^(a[190] & b[232]);
assign y[423] = (a[232] & b[191])^(a[231] & b[192])^(a[230] & b[193])^(a[229] & b[194])^(a[228] & b[195])^(a[227] & b[196])^(a[226] & b[197])^(a[225] & b[198])^(a[224] & b[199])^(a[223] & b[200])^(a[222] & b[201])^(a[221] & b[202])^(a[220] & b[203])^(a[219] & b[204])^(a[218] & b[205])^(a[217] & b[206])^(a[216] & b[207])^(a[215] & b[208])^(a[214] & b[209])^(a[213] & b[210])^(a[212] & b[211])^(a[211] & b[212])^(a[210] & b[213])^(a[209] & b[214])^(a[208] & b[215])^(a[207] & b[216])^(a[206] & b[217])^(a[205] & b[218])^(a[204] & b[219])^(a[203] & b[220])^(a[202] & b[221])^(a[201] & b[222])^(a[200] & b[223])^(a[199] & b[224])^(a[198] & b[225])^(a[197] & b[226])^(a[196] & b[227])^(a[195] & b[228])^(a[194] & b[229])^(a[193] & b[230])^(a[192] & b[231])^(a[191] & b[232]);
assign y[424] = (a[232] & b[192])^(a[231] & b[193])^(a[230] & b[194])^(a[229] & b[195])^(a[228] & b[196])^(a[227] & b[197])^(a[226] & b[198])^(a[225] & b[199])^(a[224] & b[200])^(a[223] & b[201])^(a[222] & b[202])^(a[221] & b[203])^(a[220] & b[204])^(a[219] & b[205])^(a[218] & b[206])^(a[217] & b[207])^(a[216] & b[208])^(a[215] & b[209])^(a[214] & b[210])^(a[213] & b[211])^(a[212] & b[212])^(a[211] & b[213])^(a[210] & b[214])^(a[209] & b[215])^(a[208] & b[216])^(a[207] & b[217])^(a[206] & b[218])^(a[205] & b[219])^(a[204] & b[220])^(a[203] & b[221])^(a[202] & b[222])^(a[201] & b[223])^(a[200] & b[224])^(a[199] & b[225])^(a[198] & b[226])^(a[197] & b[227])^(a[196] & b[228])^(a[195] & b[229])^(a[194] & b[230])^(a[193] & b[231])^(a[192] & b[232]);
assign y[425] = (a[232] & b[193])^(a[231] & b[194])^(a[230] & b[195])^(a[229] & b[196])^(a[228] & b[197])^(a[227] & b[198])^(a[226] & b[199])^(a[225] & b[200])^(a[224] & b[201])^(a[223] & b[202])^(a[222] & b[203])^(a[221] & b[204])^(a[220] & b[205])^(a[219] & b[206])^(a[218] & b[207])^(a[217] & b[208])^(a[216] & b[209])^(a[215] & b[210])^(a[214] & b[211])^(a[213] & b[212])^(a[212] & b[213])^(a[211] & b[214])^(a[210] & b[215])^(a[209] & b[216])^(a[208] & b[217])^(a[207] & b[218])^(a[206] & b[219])^(a[205] & b[220])^(a[204] & b[221])^(a[203] & b[222])^(a[202] & b[223])^(a[201] & b[224])^(a[200] & b[225])^(a[199] & b[226])^(a[198] & b[227])^(a[197] & b[228])^(a[196] & b[229])^(a[195] & b[230])^(a[194] & b[231])^(a[193] & b[232]);
assign y[426] = (a[232] & b[194])^(a[231] & b[195])^(a[230] & b[196])^(a[229] & b[197])^(a[228] & b[198])^(a[227] & b[199])^(a[226] & b[200])^(a[225] & b[201])^(a[224] & b[202])^(a[223] & b[203])^(a[222] & b[204])^(a[221] & b[205])^(a[220] & b[206])^(a[219] & b[207])^(a[218] & b[208])^(a[217] & b[209])^(a[216] & b[210])^(a[215] & b[211])^(a[214] & b[212])^(a[213] & b[213])^(a[212] & b[214])^(a[211] & b[215])^(a[210] & b[216])^(a[209] & b[217])^(a[208] & b[218])^(a[207] & b[219])^(a[206] & b[220])^(a[205] & b[221])^(a[204] & b[222])^(a[203] & b[223])^(a[202] & b[224])^(a[201] & b[225])^(a[200] & b[226])^(a[199] & b[227])^(a[198] & b[228])^(a[197] & b[229])^(a[196] & b[230])^(a[195] & b[231])^(a[194] & b[232]);
assign y[427] = (a[232] & b[195])^(a[231] & b[196])^(a[230] & b[197])^(a[229] & b[198])^(a[228] & b[199])^(a[227] & b[200])^(a[226] & b[201])^(a[225] & b[202])^(a[224] & b[203])^(a[223] & b[204])^(a[222] & b[205])^(a[221] & b[206])^(a[220] & b[207])^(a[219] & b[208])^(a[218] & b[209])^(a[217] & b[210])^(a[216] & b[211])^(a[215] & b[212])^(a[214] & b[213])^(a[213] & b[214])^(a[212] & b[215])^(a[211] & b[216])^(a[210] & b[217])^(a[209] & b[218])^(a[208] & b[219])^(a[207] & b[220])^(a[206] & b[221])^(a[205] & b[222])^(a[204] & b[223])^(a[203] & b[224])^(a[202] & b[225])^(a[201] & b[226])^(a[200] & b[227])^(a[199] & b[228])^(a[198] & b[229])^(a[197] & b[230])^(a[196] & b[231])^(a[195] & b[232]);
assign y[428] = (a[232] & b[196])^(a[231] & b[197])^(a[230] & b[198])^(a[229] & b[199])^(a[228] & b[200])^(a[227] & b[201])^(a[226] & b[202])^(a[225] & b[203])^(a[224] & b[204])^(a[223] & b[205])^(a[222] & b[206])^(a[221] & b[207])^(a[220] & b[208])^(a[219] & b[209])^(a[218] & b[210])^(a[217] & b[211])^(a[216] & b[212])^(a[215] & b[213])^(a[214] & b[214])^(a[213] & b[215])^(a[212] & b[216])^(a[211] & b[217])^(a[210] & b[218])^(a[209] & b[219])^(a[208] & b[220])^(a[207] & b[221])^(a[206] & b[222])^(a[205] & b[223])^(a[204] & b[224])^(a[203] & b[225])^(a[202] & b[226])^(a[201] & b[227])^(a[200] & b[228])^(a[199] & b[229])^(a[198] & b[230])^(a[197] & b[231])^(a[196] & b[232]);
assign y[429] = (a[232] & b[197])^(a[231] & b[198])^(a[230] & b[199])^(a[229] & b[200])^(a[228] & b[201])^(a[227] & b[202])^(a[226] & b[203])^(a[225] & b[204])^(a[224] & b[205])^(a[223] & b[206])^(a[222] & b[207])^(a[221] & b[208])^(a[220] & b[209])^(a[219] & b[210])^(a[218] & b[211])^(a[217] & b[212])^(a[216] & b[213])^(a[215] & b[214])^(a[214] & b[215])^(a[213] & b[216])^(a[212] & b[217])^(a[211] & b[218])^(a[210] & b[219])^(a[209] & b[220])^(a[208] & b[221])^(a[207] & b[222])^(a[206] & b[223])^(a[205] & b[224])^(a[204] & b[225])^(a[203] & b[226])^(a[202] & b[227])^(a[201] & b[228])^(a[200] & b[229])^(a[199] & b[230])^(a[198] & b[231])^(a[197] & b[232]);
assign y[430] = (a[232] & b[198])^(a[231] & b[199])^(a[230] & b[200])^(a[229] & b[201])^(a[228] & b[202])^(a[227] & b[203])^(a[226] & b[204])^(a[225] & b[205])^(a[224] & b[206])^(a[223] & b[207])^(a[222] & b[208])^(a[221] & b[209])^(a[220] & b[210])^(a[219] & b[211])^(a[218] & b[212])^(a[217] & b[213])^(a[216] & b[214])^(a[215] & b[215])^(a[214] & b[216])^(a[213] & b[217])^(a[212] & b[218])^(a[211] & b[219])^(a[210] & b[220])^(a[209] & b[221])^(a[208] & b[222])^(a[207] & b[223])^(a[206] & b[224])^(a[205] & b[225])^(a[204] & b[226])^(a[203] & b[227])^(a[202] & b[228])^(a[201] & b[229])^(a[200] & b[230])^(a[199] & b[231])^(a[198] & b[232]);
assign y[431] = (a[232] & b[199])^(a[231] & b[200])^(a[230] & b[201])^(a[229] & b[202])^(a[228] & b[203])^(a[227] & b[204])^(a[226] & b[205])^(a[225] & b[206])^(a[224] & b[207])^(a[223] & b[208])^(a[222] & b[209])^(a[221] & b[210])^(a[220] & b[211])^(a[219] & b[212])^(a[218] & b[213])^(a[217] & b[214])^(a[216] & b[215])^(a[215] & b[216])^(a[214] & b[217])^(a[213] & b[218])^(a[212] & b[219])^(a[211] & b[220])^(a[210] & b[221])^(a[209] & b[222])^(a[208] & b[223])^(a[207] & b[224])^(a[206] & b[225])^(a[205] & b[226])^(a[204] & b[227])^(a[203] & b[228])^(a[202] & b[229])^(a[201] & b[230])^(a[200] & b[231])^(a[199] & b[232]);
assign y[432] = (a[232] & b[200])^(a[231] & b[201])^(a[230] & b[202])^(a[229] & b[203])^(a[228] & b[204])^(a[227] & b[205])^(a[226] & b[206])^(a[225] & b[207])^(a[224] & b[208])^(a[223] & b[209])^(a[222] & b[210])^(a[221] & b[211])^(a[220] & b[212])^(a[219] & b[213])^(a[218] & b[214])^(a[217] & b[215])^(a[216] & b[216])^(a[215] & b[217])^(a[214] & b[218])^(a[213] & b[219])^(a[212] & b[220])^(a[211] & b[221])^(a[210] & b[222])^(a[209] & b[223])^(a[208] & b[224])^(a[207] & b[225])^(a[206] & b[226])^(a[205] & b[227])^(a[204] & b[228])^(a[203] & b[229])^(a[202] & b[230])^(a[201] & b[231])^(a[200] & b[232]);
assign y[433] = (a[232] & b[201])^(a[231] & b[202])^(a[230] & b[203])^(a[229] & b[204])^(a[228] & b[205])^(a[227] & b[206])^(a[226] & b[207])^(a[225] & b[208])^(a[224] & b[209])^(a[223] & b[210])^(a[222] & b[211])^(a[221] & b[212])^(a[220] & b[213])^(a[219] & b[214])^(a[218] & b[215])^(a[217] & b[216])^(a[216] & b[217])^(a[215] & b[218])^(a[214] & b[219])^(a[213] & b[220])^(a[212] & b[221])^(a[211] & b[222])^(a[210] & b[223])^(a[209] & b[224])^(a[208] & b[225])^(a[207] & b[226])^(a[206] & b[227])^(a[205] & b[228])^(a[204] & b[229])^(a[203] & b[230])^(a[202] & b[231])^(a[201] & b[232]);
assign y[434] = (a[232] & b[202])^(a[231] & b[203])^(a[230] & b[204])^(a[229] & b[205])^(a[228] & b[206])^(a[227] & b[207])^(a[226] & b[208])^(a[225] & b[209])^(a[224] & b[210])^(a[223] & b[211])^(a[222] & b[212])^(a[221] & b[213])^(a[220] & b[214])^(a[219] & b[215])^(a[218] & b[216])^(a[217] & b[217])^(a[216] & b[218])^(a[215] & b[219])^(a[214] & b[220])^(a[213] & b[221])^(a[212] & b[222])^(a[211] & b[223])^(a[210] & b[224])^(a[209] & b[225])^(a[208] & b[226])^(a[207] & b[227])^(a[206] & b[228])^(a[205] & b[229])^(a[204] & b[230])^(a[203] & b[231])^(a[202] & b[232]);
assign y[435] = (a[232] & b[203])^(a[231] & b[204])^(a[230] & b[205])^(a[229] & b[206])^(a[228] & b[207])^(a[227] & b[208])^(a[226] & b[209])^(a[225] & b[210])^(a[224] & b[211])^(a[223] & b[212])^(a[222] & b[213])^(a[221] & b[214])^(a[220] & b[215])^(a[219] & b[216])^(a[218] & b[217])^(a[217] & b[218])^(a[216] & b[219])^(a[215] & b[220])^(a[214] & b[221])^(a[213] & b[222])^(a[212] & b[223])^(a[211] & b[224])^(a[210] & b[225])^(a[209] & b[226])^(a[208] & b[227])^(a[207] & b[228])^(a[206] & b[229])^(a[205] & b[230])^(a[204] & b[231])^(a[203] & b[232]);
assign y[436] = (a[232] & b[204])^(a[231] & b[205])^(a[230] & b[206])^(a[229] & b[207])^(a[228] & b[208])^(a[227] & b[209])^(a[226] & b[210])^(a[225] & b[211])^(a[224] & b[212])^(a[223] & b[213])^(a[222] & b[214])^(a[221] & b[215])^(a[220] & b[216])^(a[219] & b[217])^(a[218] & b[218])^(a[217] & b[219])^(a[216] & b[220])^(a[215] & b[221])^(a[214] & b[222])^(a[213] & b[223])^(a[212] & b[224])^(a[211] & b[225])^(a[210] & b[226])^(a[209] & b[227])^(a[208] & b[228])^(a[207] & b[229])^(a[206] & b[230])^(a[205] & b[231])^(a[204] & b[232]);
assign y[437] = (a[232] & b[205])^(a[231] & b[206])^(a[230] & b[207])^(a[229] & b[208])^(a[228] & b[209])^(a[227] & b[210])^(a[226] & b[211])^(a[225] & b[212])^(a[224] & b[213])^(a[223] & b[214])^(a[222] & b[215])^(a[221] & b[216])^(a[220] & b[217])^(a[219] & b[218])^(a[218] & b[219])^(a[217] & b[220])^(a[216] & b[221])^(a[215] & b[222])^(a[214] & b[223])^(a[213] & b[224])^(a[212] & b[225])^(a[211] & b[226])^(a[210] & b[227])^(a[209] & b[228])^(a[208] & b[229])^(a[207] & b[230])^(a[206] & b[231])^(a[205] & b[232]);
assign y[438] = (a[232] & b[206])^(a[231] & b[207])^(a[230] & b[208])^(a[229] & b[209])^(a[228] & b[210])^(a[227] & b[211])^(a[226] & b[212])^(a[225] & b[213])^(a[224] & b[214])^(a[223] & b[215])^(a[222] & b[216])^(a[221] & b[217])^(a[220] & b[218])^(a[219] & b[219])^(a[218] & b[220])^(a[217] & b[221])^(a[216] & b[222])^(a[215] & b[223])^(a[214] & b[224])^(a[213] & b[225])^(a[212] & b[226])^(a[211] & b[227])^(a[210] & b[228])^(a[209] & b[229])^(a[208] & b[230])^(a[207] & b[231])^(a[206] & b[232]);
assign y[439] = (a[232] & b[207])^(a[231] & b[208])^(a[230] & b[209])^(a[229] & b[210])^(a[228] & b[211])^(a[227] & b[212])^(a[226] & b[213])^(a[225] & b[214])^(a[224] & b[215])^(a[223] & b[216])^(a[222] & b[217])^(a[221] & b[218])^(a[220] & b[219])^(a[219] & b[220])^(a[218] & b[221])^(a[217] & b[222])^(a[216] & b[223])^(a[215] & b[224])^(a[214] & b[225])^(a[213] & b[226])^(a[212] & b[227])^(a[211] & b[228])^(a[210] & b[229])^(a[209] & b[230])^(a[208] & b[231])^(a[207] & b[232]);
assign y[440] = (a[232] & b[208])^(a[231] & b[209])^(a[230] & b[210])^(a[229] & b[211])^(a[228] & b[212])^(a[227] & b[213])^(a[226] & b[214])^(a[225] & b[215])^(a[224] & b[216])^(a[223] & b[217])^(a[222] & b[218])^(a[221] & b[219])^(a[220] & b[220])^(a[219] & b[221])^(a[218] & b[222])^(a[217] & b[223])^(a[216] & b[224])^(a[215] & b[225])^(a[214] & b[226])^(a[213] & b[227])^(a[212] & b[228])^(a[211] & b[229])^(a[210] & b[230])^(a[209] & b[231])^(a[208] & b[232]);
assign y[441] = (a[232] & b[209])^(a[231] & b[210])^(a[230] & b[211])^(a[229] & b[212])^(a[228] & b[213])^(a[227] & b[214])^(a[226] & b[215])^(a[225] & b[216])^(a[224] & b[217])^(a[223] & b[218])^(a[222] & b[219])^(a[221] & b[220])^(a[220] & b[221])^(a[219] & b[222])^(a[218] & b[223])^(a[217] & b[224])^(a[216] & b[225])^(a[215] & b[226])^(a[214] & b[227])^(a[213] & b[228])^(a[212] & b[229])^(a[211] & b[230])^(a[210] & b[231])^(a[209] & b[232]);
assign y[442] = (a[232] & b[210])^(a[231] & b[211])^(a[230] & b[212])^(a[229] & b[213])^(a[228] & b[214])^(a[227] & b[215])^(a[226] & b[216])^(a[225] & b[217])^(a[224] & b[218])^(a[223] & b[219])^(a[222] & b[220])^(a[221] & b[221])^(a[220] & b[222])^(a[219] & b[223])^(a[218] & b[224])^(a[217] & b[225])^(a[216] & b[226])^(a[215] & b[227])^(a[214] & b[228])^(a[213] & b[229])^(a[212] & b[230])^(a[211] & b[231])^(a[210] & b[232]);
assign y[443] = (a[232] & b[211])^(a[231] & b[212])^(a[230] & b[213])^(a[229] & b[214])^(a[228] & b[215])^(a[227] & b[216])^(a[226] & b[217])^(a[225] & b[218])^(a[224] & b[219])^(a[223] & b[220])^(a[222] & b[221])^(a[221] & b[222])^(a[220] & b[223])^(a[219] & b[224])^(a[218] & b[225])^(a[217] & b[226])^(a[216] & b[227])^(a[215] & b[228])^(a[214] & b[229])^(a[213] & b[230])^(a[212] & b[231])^(a[211] & b[232]);
assign y[444] = (a[232] & b[212])^(a[231] & b[213])^(a[230] & b[214])^(a[229] & b[215])^(a[228] & b[216])^(a[227] & b[217])^(a[226] & b[218])^(a[225] & b[219])^(a[224] & b[220])^(a[223] & b[221])^(a[222] & b[222])^(a[221] & b[223])^(a[220] & b[224])^(a[219] & b[225])^(a[218] & b[226])^(a[217] & b[227])^(a[216] & b[228])^(a[215] & b[229])^(a[214] & b[230])^(a[213] & b[231])^(a[212] & b[232]);
assign y[445] = (a[232] & b[213])^(a[231] & b[214])^(a[230] & b[215])^(a[229] & b[216])^(a[228] & b[217])^(a[227] & b[218])^(a[226] & b[219])^(a[225] & b[220])^(a[224] & b[221])^(a[223] & b[222])^(a[222] & b[223])^(a[221] & b[224])^(a[220] & b[225])^(a[219] & b[226])^(a[218] & b[227])^(a[217] & b[228])^(a[216] & b[229])^(a[215] & b[230])^(a[214] & b[231])^(a[213] & b[232]);
assign y[446] = (a[232] & b[214])^(a[231] & b[215])^(a[230] & b[216])^(a[229] & b[217])^(a[228] & b[218])^(a[227] & b[219])^(a[226] & b[220])^(a[225] & b[221])^(a[224] & b[222])^(a[223] & b[223])^(a[222] & b[224])^(a[221] & b[225])^(a[220] & b[226])^(a[219] & b[227])^(a[218] & b[228])^(a[217] & b[229])^(a[216] & b[230])^(a[215] & b[231])^(a[214] & b[232]);
assign y[447] = (a[232] & b[215])^(a[231] & b[216])^(a[230] & b[217])^(a[229] & b[218])^(a[228] & b[219])^(a[227] & b[220])^(a[226] & b[221])^(a[225] & b[222])^(a[224] & b[223])^(a[223] & b[224])^(a[222] & b[225])^(a[221] & b[226])^(a[220] & b[227])^(a[219] & b[228])^(a[218] & b[229])^(a[217] & b[230])^(a[216] & b[231])^(a[215] & b[232]);
assign y[448] = (a[232] & b[216])^(a[231] & b[217])^(a[230] & b[218])^(a[229] & b[219])^(a[228] & b[220])^(a[227] & b[221])^(a[226] & b[222])^(a[225] & b[223])^(a[224] & b[224])^(a[223] & b[225])^(a[222] & b[226])^(a[221] & b[227])^(a[220] & b[228])^(a[219] & b[229])^(a[218] & b[230])^(a[217] & b[231])^(a[216] & b[232]);
assign y[449] = (a[232] & b[217])^(a[231] & b[218])^(a[230] & b[219])^(a[229] & b[220])^(a[228] & b[221])^(a[227] & b[222])^(a[226] & b[223])^(a[225] & b[224])^(a[224] & b[225])^(a[223] & b[226])^(a[222] & b[227])^(a[221] & b[228])^(a[220] & b[229])^(a[219] & b[230])^(a[218] & b[231])^(a[217] & b[232]);
assign y[450] = (a[232] & b[218])^(a[231] & b[219])^(a[230] & b[220])^(a[229] & b[221])^(a[228] & b[222])^(a[227] & b[223])^(a[226] & b[224])^(a[225] & b[225])^(a[224] & b[226])^(a[223] & b[227])^(a[222] & b[228])^(a[221] & b[229])^(a[220] & b[230])^(a[219] & b[231])^(a[218] & b[232]);
assign y[451] = (a[232] & b[219])^(a[231] & b[220])^(a[230] & b[221])^(a[229] & b[222])^(a[228] & b[223])^(a[227] & b[224])^(a[226] & b[225])^(a[225] & b[226])^(a[224] & b[227])^(a[223] & b[228])^(a[222] & b[229])^(a[221] & b[230])^(a[220] & b[231])^(a[219] & b[232]);
assign y[452] = (a[232] & b[220])^(a[231] & b[221])^(a[230] & b[222])^(a[229] & b[223])^(a[228] & b[224])^(a[227] & b[225])^(a[226] & b[226])^(a[225] & b[227])^(a[224] & b[228])^(a[223] & b[229])^(a[222] & b[230])^(a[221] & b[231])^(a[220] & b[232]);
assign y[453] = (a[232] & b[221])^(a[231] & b[222])^(a[230] & b[223])^(a[229] & b[224])^(a[228] & b[225])^(a[227] & b[226])^(a[226] & b[227])^(a[225] & b[228])^(a[224] & b[229])^(a[223] & b[230])^(a[222] & b[231])^(a[221] & b[232]);
assign y[454] = (a[232] & b[222])^(a[231] & b[223])^(a[230] & b[224])^(a[229] & b[225])^(a[228] & b[226])^(a[227] & b[227])^(a[226] & b[228])^(a[225] & b[229])^(a[224] & b[230])^(a[223] & b[231])^(a[222] & b[232]);
assign y[455] = (a[232] & b[223])^(a[231] & b[224])^(a[230] & b[225])^(a[229] & b[226])^(a[228] & b[227])^(a[227] & b[228])^(a[226] & b[229])^(a[225] & b[230])^(a[224] & b[231])^(a[223] & b[232]);
assign y[456] = (a[232] & b[224])^(a[231] & b[225])^(a[230] & b[226])^(a[229] & b[227])^(a[228] & b[228])^(a[227] & b[229])^(a[226] & b[230])^(a[225] & b[231])^(a[224] & b[232]);
assign y[457] = (a[232] & b[225])^(a[231] & b[226])^(a[230] & b[227])^(a[229] & b[228])^(a[228] & b[229])^(a[227] & b[230])^(a[226] & b[231])^(a[225] & b[232]);
assign y[458] = (a[232] & b[226])^(a[231] & b[227])^(a[230] & b[228])^(a[229] & b[229])^(a[228] & b[230])^(a[227] & b[231])^(a[226] & b[232]);
assign y[459] = (a[232] & b[227])^(a[231] & b[228])^(a[230] & b[229])^(a[229] & b[230])^(a[228] & b[231])^(a[227] & b[232]);
assign y[460] = (a[232] & b[228])^(a[231] & b[229])^(a[230] & b[230])^(a[229] & b[231])^(a[228] & b[232]);
assign y[461] = (a[232] & b[229])^(a[231] & b[230])^(a[230] & b[231])^(a[229] & b[232]);
assign y[462] = (a[232] & b[230])^(a[231] & b[231])^(a[230] & b[232]);
assign y[463] = (a[232] & b[231])^(a[231] & b[232]);
assign y[464] = (a[232] & b[232]);



endmodule
