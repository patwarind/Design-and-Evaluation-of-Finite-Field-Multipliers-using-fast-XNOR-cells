`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Nitin D. Patwari
// 
// Create Date: 20.01.2022 22:25:39
// Design Name: 
// Module Name: CA_409bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CA_409bit(
    a,
    b,
    y
    );

input [408:0] a;
input [408:0] b;

output [816:0] y;




assign y[0] = (a[0] & b[0]);
assign y[1] = (a[1] & b[0])^(a[0] & b[1]);
assign y[2] = (a[2] & b[0])^(a[1] & b[1])^(a[0] & b[2]);
assign y[3] = (a[3] & b[0])^(a[2] & b[1])^(a[1] & b[2])^(a[0] & b[3]);
assign y[4] = (a[4] & b[0])^(a[3] & b[1])^(a[2] & b[2])^(a[1] & b[3])^(a[0] & b[4]);
assign y[5] = (a[5] & b[0])^(a[4] & b[1])^(a[3] & b[2])^(a[2] & b[3])^(a[1] & b[4])^(a[0] & b[5]);
assign y[6] = (a[6] & b[0])^(a[5] & b[1])^(a[4] & b[2])^(a[3] & b[3])^(a[2] & b[4])^(a[1] & b[5])^(a[0] & b[6]);
assign y[7] = (a[7] & b[0])^(a[6] & b[1])^(a[5] & b[2])^(a[4] & b[3])^(a[3] & b[4])^(a[2] & b[5])^(a[1] & b[6])^(a[0] & b[7]);
assign y[8] = (a[8] & b[0])^(a[7] & b[1])^(a[6] & b[2])^(a[5] & b[3])^(a[4] & b[4])^(a[3] & b[5])^(a[2] & b[6])^(a[1] & b[7])^(a[0] & b[8]);
assign y[9] = (a[9] & b[0])^(a[8] & b[1])^(a[7] & b[2])^(a[6] & b[3])^(a[5] & b[4])^(a[4] & b[5])^(a[3] & b[6])^(a[2] & b[7])^(a[1] & b[8])^(a[0] & b[9]);
assign y[10] = (a[10] & b[0])^(a[9] & b[1])^(a[8] & b[2])^(a[7] & b[3])^(a[6] & b[4])^(a[5] & b[5])^(a[4] & b[6])^(a[3] & b[7])^(a[2] & b[8])^(a[1] & b[9])^(a[0] & b[10]);
assign y[11] = (a[11] & b[0])^(a[10] & b[1])^(a[9] & b[2])^(a[8] & b[3])^(a[7] & b[4])^(a[6] & b[5])^(a[5] & b[6])^(a[4] & b[7])^(a[3] & b[8])^(a[2] & b[9])^(a[1] & b[10])^(a[0] & b[11]);
assign y[12] = (a[12] & b[0])^(a[11] & b[1])^(a[10] & b[2])^(a[9] & b[3])^(a[8] & b[4])^(a[7] & b[5])^(a[6] & b[6])^(a[5] & b[7])^(a[4] & b[8])^(a[3] & b[9])^(a[2] & b[10])^(a[1] & b[11])^(a[0] & b[12]);
assign y[13] = (a[13] & b[0])^(a[12] & b[1])^(a[11] & b[2])^(a[10] & b[3])^(a[9] & b[4])^(a[8] & b[5])^(a[7] & b[6])^(a[6] & b[7])^(a[5] & b[8])^(a[4] & b[9])^(a[3] & b[10])^(a[2] & b[11])^(a[1] & b[12])^(a[0] & b[13]);
assign y[14] = (a[14] & b[0])^(a[13] & b[1])^(a[12] & b[2])^(a[11] & b[3])^(a[10] & b[4])^(a[9] & b[5])^(a[8] & b[6])^(a[7] & b[7])^(a[6] & b[8])^(a[5] & b[9])^(a[4] & b[10])^(a[3] & b[11])^(a[2] & b[12])^(a[1] & b[13])^(a[0] & b[14]);
assign y[15] = (a[15] & b[0])^(a[14] & b[1])^(a[13] & b[2])^(a[12] & b[3])^(a[11] & b[4])^(a[10] & b[5])^(a[9] & b[6])^(a[8] & b[7])^(a[7] & b[8])^(a[6] & b[9])^(a[5] & b[10])^(a[4] & b[11])^(a[3] & b[12])^(a[2] & b[13])^(a[1] & b[14])^(a[0] & b[15]);
assign y[16] = (a[16] & b[0])^(a[15] & b[1])^(a[14] & b[2])^(a[13] & b[3])^(a[12] & b[4])^(a[11] & b[5])^(a[10] & b[6])^(a[9] & b[7])^(a[8] & b[8])^(a[7] & b[9])^(a[6] & b[10])^(a[5] & b[11])^(a[4] & b[12])^(a[3] & b[13])^(a[2] & b[14])^(a[1] & b[15])^(a[0] & b[16]);
assign y[17] = (a[17] & b[0])^(a[16] & b[1])^(a[15] & b[2])^(a[14] & b[3])^(a[13] & b[4])^(a[12] & b[5])^(a[11] & b[6])^(a[10] & b[7])^(a[9] & b[8])^(a[8] & b[9])^(a[7] & b[10])^(a[6] & b[11])^(a[5] & b[12])^(a[4] & b[13])^(a[3] & b[14])^(a[2] & b[15])^(a[1] & b[16])^(a[0] & b[17]);
assign y[18] = (a[18] & b[0])^(a[17] & b[1])^(a[16] & b[2])^(a[15] & b[3])^(a[14] & b[4])^(a[13] & b[5])^(a[12] & b[6])^(a[11] & b[7])^(a[10] & b[8])^(a[9] & b[9])^(a[8] & b[10])^(a[7] & b[11])^(a[6] & b[12])^(a[5] & b[13])^(a[4] & b[14])^(a[3] & b[15])^(a[2] & b[16])^(a[1] & b[17])^(a[0] & b[18]);
assign y[19] = (a[19] & b[0])^(a[18] & b[1])^(a[17] & b[2])^(a[16] & b[3])^(a[15] & b[4])^(a[14] & b[5])^(a[13] & b[6])^(a[12] & b[7])^(a[11] & b[8])^(a[10] & b[9])^(a[9] & b[10])^(a[8] & b[11])^(a[7] & b[12])^(a[6] & b[13])^(a[5] & b[14])^(a[4] & b[15])^(a[3] & b[16])^(a[2] & b[17])^(a[1] & b[18])^(a[0] & b[19]);
assign y[20] = (a[20] & b[0])^(a[19] & b[1])^(a[18] & b[2])^(a[17] & b[3])^(a[16] & b[4])^(a[15] & b[5])^(a[14] & b[6])^(a[13] & b[7])^(a[12] & b[8])^(a[11] & b[9])^(a[10] & b[10])^(a[9] & b[11])^(a[8] & b[12])^(a[7] & b[13])^(a[6] & b[14])^(a[5] & b[15])^(a[4] & b[16])^(a[3] & b[17])^(a[2] & b[18])^(a[1] & b[19])^(a[0] & b[20]);
assign y[21] = (a[21] & b[0])^(a[20] & b[1])^(a[19] & b[2])^(a[18] & b[3])^(a[17] & b[4])^(a[16] & b[5])^(a[15] & b[6])^(a[14] & b[7])^(a[13] & b[8])^(a[12] & b[9])^(a[11] & b[10])^(a[10] & b[11])^(a[9] & b[12])^(a[8] & b[13])^(a[7] & b[14])^(a[6] & b[15])^(a[5] & b[16])^(a[4] & b[17])^(a[3] & b[18])^(a[2] & b[19])^(a[1] & b[20])^(a[0] & b[21]);
assign y[22] = (a[22] & b[0])^(a[21] & b[1])^(a[20] & b[2])^(a[19] & b[3])^(a[18] & b[4])^(a[17] & b[5])^(a[16] & b[6])^(a[15] & b[7])^(a[14] & b[8])^(a[13] & b[9])^(a[12] & b[10])^(a[11] & b[11])^(a[10] & b[12])^(a[9] & b[13])^(a[8] & b[14])^(a[7] & b[15])^(a[6] & b[16])^(a[5] & b[17])^(a[4] & b[18])^(a[3] & b[19])^(a[2] & b[20])^(a[1] & b[21])^(a[0] & b[22]);
assign y[23] = (a[23] & b[0])^(a[22] & b[1])^(a[21] & b[2])^(a[20] & b[3])^(a[19] & b[4])^(a[18] & b[5])^(a[17] & b[6])^(a[16] & b[7])^(a[15] & b[8])^(a[14] & b[9])^(a[13] & b[10])^(a[12] & b[11])^(a[11] & b[12])^(a[10] & b[13])^(a[9] & b[14])^(a[8] & b[15])^(a[7] & b[16])^(a[6] & b[17])^(a[5] & b[18])^(a[4] & b[19])^(a[3] & b[20])^(a[2] & b[21])^(a[1] & b[22])^(a[0] & b[23]);
assign y[24] = (a[24] & b[0])^(a[23] & b[1])^(a[22] & b[2])^(a[21] & b[3])^(a[20] & b[4])^(a[19] & b[5])^(a[18] & b[6])^(a[17] & b[7])^(a[16] & b[8])^(a[15] & b[9])^(a[14] & b[10])^(a[13] & b[11])^(a[12] & b[12])^(a[11] & b[13])^(a[10] & b[14])^(a[9] & b[15])^(a[8] & b[16])^(a[7] & b[17])^(a[6] & b[18])^(a[5] & b[19])^(a[4] & b[20])^(a[3] & b[21])^(a[2] & b[22])^(a[1] & b[23])^(a[0] & b[24]);
assign y[25] = (a[25] & b[0])^(a[24] & b[1])^(a[23] & b[2])^(a[22] & b[3])^(a[21] & b[4])^(a[20] & b[5])^(a[19] & b[6])^(a[18] & b[7])^(a[17] & b[8])^(a[16] & b[9])^(a[15] & b[10])^(a[14] & b[11])^(a[13] & b[12])^(a[12] & b[13])^(a[11] & b[14])^(a[10] & b[15])^(a[9] & b[16])^(a[8] & b[17])^(a[7] & b[18])^(a[6] & b[19])^(a[5] & b[20])^(a[4] & b[21])^(a[3] & b[22])^(a[2] & b[23])^(a[1] & b[24])^(a[0] & b[25]);
assign y[26] = (a[26] & b[0])^(a[25] & b[1])^(a[24] & b[2])^(a[23] & b[3])^(a[22] & b[4])^(a[21] & b[5])^(a[20] & b[6])^(a[19] & b[7])^(a[18] & b[8])^(a[17] & b[9])^(a[16] & b[10])^(a[15] & b[11])^(a[14] & b[12])^(a[13] & b[13])^(a[12] & b[14])^(a[11] & b[15])^(a[10] & b[16])^(a[9] & b[17])^(a[8] & b[18])^(a[7] & b[19])^(a[6] & b[20])^(a[5] & b[21])^(a[4] & b[22])^(a[3] & b[23])^(a[2] & b[24])^(a[1] & b[25])^(a[0] & b[26]);
assign y[27] = (a[27] & b[0])^(a[26] & b[1])^(a[25] & b[2])^(a[24] & b[3])^(a[23] & b[4])^(a[22] & b[5])^(a[21] & b[6])^(a[20] & b[7])^(a[19] & b[8])^(a[18] & b[9])^(a[17] & b[10])^(a[16] & b[11])^(a[15] & b[12])^(a[14] & b[13])^(a[13] & b[14])^(a[12] & b[15])^(a[11] & b[16])^(a[10] & b[17])^(a[9] & b[18])^(a[8] & b[19])^(a[7] & b[20])^(a[6] & b[21])^(a[5] & b[22])^(a[4] & b[23])^(a[3] & b[24])^(a[2] & b[25])^(a[1] & b[26])^(a[0] & b[27]);
assign y[28] = (a[28] & b[0])^(a[27] & b[1])^(a[26] & b[2])^(a[25] & b[3])^(a[24] & b[4])^(a[23] & b[5])^(a[22] & b[6])^(a[21] & b[7])^(a[20] & b[8])^(a[19] & b[9])^(a[18] & b[10])^(a[17] & b[11])^(a[16] & b[12])^(a[15] & b[13])^(a[14] & b[14])^(a[13] & b[15])^(a[12] & b[16])^(a[11] & b[17])^(a[10] & b[18])^(a[9] & b[19])^(a[8] & b[20])^(a[7] & b[21])^(a[6] & b[22])^(a[5] & b[23])^(a[4] & b[24])^(a[3] & b[25])^(a[2] & b[26])^(a[1] & b[27])^(a[0] & b[28]);
assign y[29] = (a[29] & b[0])^(a[28] & b[1])^(a[27] & b[2])^(a[26] & b[3])^(a[25] & b[4])^(a[24] & b[5])^(a[23] & b[6])^(a[22] & b[7])^(a[21] & b[8])^(a[20] & b[9])^(a[19] & b[10])^(a[18] & b[11])^(a[17] & b[12])^(a[16] & b[13])^(a[15] & b[14])^(a[14] & b[15])^(a[13] & b[16])^(a[12] & b[17])^(a[11] & b[18])^(a[10] & b[19])^(a[9] & b[20])^(a[8] & b[21])^(a[7] & b[22])^(a[6] & b[23])^(a[5] & b[24])^(a[4] & b[25])^(a[3] & b[26])^(a[2] & b[27])^(a[1] & b[28])^(a[0] & b[29]);
assign y[30] = (a[30] & b[0])^(a[29] & b[1])^(a[28] & b[2])^(a[27] & b[3])^(a[26] & b[4])^(a[25] & b[5])^(a[24] & b[6])^(a[23] & b[7])^(a[22] & b[8])^(a[21] & b[9])^(a[20] & b[10])^(a[19] & b[11])^(a[18] & b[12])^(a[17] & b[13])^(a[16] & b[14])^(a[15] & b[15])^(a[14] & b[16])^(a[13] & b[17])^(a[12] & b[18])^(a[11] & b[19])^(a[10] & b[20])^(a[9] & b[21])^(a[8] & b[22])^(a[7] & b[23])^(a[6] & b[24])^(a[5] & b[25])^(a[4] & b[26])^(a[3] & b[27])^(a[2] & b[28])^(a[1] & b[29])^(a[0] & b[30]);
assign y[31] = (a[31] & b[0])^(a[30] & b[1])^(a[29] & b[2])^(a[28] & b[3])^(a[27] & b[4])^(a[26] & b[5])^(a[25] & b[6])^(a[24] & b[7])^(a[23] & b[8])^(a[22] & b[9])^(a[21] & b[10])^(a[20] & b[11])^(a[19] & b[12])^(a[18] & b[13])^(a[17] & b[14])^(a[16] & b[15])^(a[15] & b[16])^(a[14] & b[17])^(a[13] & b[18])^(a[12] & b[19])^(a[11] & b[20])^(a[10] & b[21])^(a[9] & b[22])^(a[8] & b[23])^(a[7] & b[24])^(a[6] & b[25])^(a[5] & b[26])^(a[4] & b[27])^(a[3] & b[28])^(a[2] & b[29])^(a[1] & b[30])^(a[0] & b[31]);
assign y[32] = (a[32] & b[0])^(a[31] & b[1])^(a[30] & b[2])^(a[29] & b[3])^(a[28] & b[4])^(a[27] & b[5])^(a[26] & b[6])^(a[25] & b[7])^(a[24] & b[8])^(a[23] & b[9])^(a[22] & b[10])^(a[21] & b[11])^(a[20] & b[12])^(a[19] & b[13])^(a[18] & b[14])^(a[17] & b[15])^(a[16] & b[16])^(a[15] & b[17])^(a[14] & b[18])^(a[13] & b[19])^(a[12] & b[20])^(a[11] & b[21])^(a[10] & b[22])^(a[9] & b[23])^(a[8] & b[24])^(a[7] & b[25])^(a[6] & b[26])^(a[5] & b[27])^(a[4] & b[28])^(a[3] & b[29])^(a[2] & b[30])^(a[1] & b[31])^(a[0] & b[32]);
assign y[33] = (a[33] & b[0])^(a[32] & b[1])^(a[31] & b[2])^(a[30] & b[3])^(a[29] & b[4])^(a[28] & b[5])^(a[27] & b[6])^(a[26] & b[7])^(a[25] & b[8])^(a[24] & b[9])^(a[23] & b[10])^(a[22] & b[11])^(a[21] & b[12])^(a[20] & b[13])^(a[19] & b[14])^(a[18] & b[15])^(a[17] & b[16])^(a[16] & b[17])^(a[15] & b[18])^(a[14] & b[19])^(a[13] & b[20])^(a[12] & b[21])^(a[11] & b[22])^(a[10] & b[23])^(a[9] & b[24])^(a[8] & b[25])^(a[7] & b[26])^(a[6] & b[27])^(a[5] & b[28])^(a[4] & b[29])^(a[3] & b[30])^(a[2] & b[31])^(a[1] & b[32])^(a[0] & b[33]);
assign y[34] = (a[34] & b[0])^(a[33] & b[1])^(a[32] & b[2])^(a[31] & b[3])^(a[30] & b[4])^(a[29] & b[5])^(a[28] & b[6])^(a[27] & b[7])^(a[26] & b[8])^(a[25] & b[9])^(a[24] & b[10])^(a[23] & b[11])^(a[22] & b[12])^(a[21] & b[13])^(a[20] & b[14])^(a[19] & b[15])^(a[18] & b[16])^(a[17] & b[17])^(a[16] & b[18])^(a[15] & b[19])^(a[14] & b[20])^(a[13] & b[21])^(a[12] & b[22])^(a[11] & b[23])^(a[10] & b[24])^(a[9] & b[25])^(a[8] & b[26])^(a[7] & b[27])^(a[6] & b[28])^(a[5] & b[29])^(a[4] & b[30])^(a[3] & b[31])^(a[2] & b[32])^(a[1] & b[33])^(a[0] & b[34]);
assign y[35] = (a[35] & b[0])^(a[34] & b[1])^(a[33] & b[2])^(a[32] & b[3])^(a[31] & b[4])^(a[30] & b[5])^(a[29] & b[6])^(a[28] & b[7])^(a[27] & b[8])^(a[26] & b[9])^(a[25] & b[10])^(a[24] & b[11])^(a[23] & b[12])^(a[22] & b[13])^(a[21] & b[14])^(a[20] & b[15])^(a[19] & b[16])^(a[18] & b[17])^(a[17] & b[18])^(a[16] & b[19])^(a[15] & b[20])^(a[14] & b[21])^(a[13] & b[22])^(a[12] & b[23])^(a[11] & b[24])^(a[10] & b[25])^(a[9] & b[26])^(a[8] & b[27])^(a[7] & b[28])^(a[6] & b[29])^(a[5] & b[30])^(a[4] & b[31])^(a[3] & b[32])^(a[2] & b[33])^(a[1] & b[34])^(a[0] & b[35]);
assign y[36] = (a[36] & b[0])^(a[35] & b[1])^(a[34] & b[2])^(a[33] & b[3])^(a[32] & b[4])^(a[31] & b[5])^(a[30] & b[6])^(a[29] & b[7])^(a[28] & b[8])^(a[27] & b[9])^(a[26] & b[10])^(a[25] & b[11])^(a[24] & b[12])^(a[23] & b[13])^(a[22] & b[14])^(a[21] & b[15])^(a[20] & b[16])^(a[19] & b[17])^(a[18] & b[18])^(a[17] & b[19])^(a[16] & b[20])^(a[15] & b[21])^(a[14] & b[22])^(a[13] & b[23])^(a[12] & b[24])^(a[11] & b[25])^(a[10] & b[26])^(a[9] & b[27])^(a[8] & b[28])^(a[7] & b[29])^(a[6] & b[30])^(a[5] & b[31])^(a[4] & b[32])^(a[3] & b[33])^(a[2] & b[34])^(a[1] & b[35])^(a[0] & b[36]);
assign y[37] = (a[37] & b[0])^(a[36] & b[1])^(a[35] & b[2])^(a[34] & b[3])^(a[33] & b[4])^(a[32] & b[5])^(a[31] & b[6])^(a[30] & b[7])^(a[29] & b[8])^(a[28] & b[9])^(a[27] & b[10])^(a[26] & b[11])^(a[25] & b[12])^(a[24] & b[13])^(a[23] & b[14])^(a[22] & b[15])^(a[21] & b[16])^(a[20] & b[17])^(a[19] & b[18])^(a[18] & b[19])^(a[17] & b[20])^(a[16] & b[21])^(a[15] & b[22])^(a[14] & b[23])^(a[13] & b[24])^(a[12] & b[25])^(a[11] & b[26])^(a[10] & b[27])^(a[9] & b[28])^(a[8] & b[29])^(a[7] & b[30])^(a[6] & b[31])^(a[5] & b[32])^(a[4] & b[33])^(a[3] & b[34])^(a[2] & b[35])^(a[1] & b[36])^(a[0] & b[37]);
assign y[38] = (a[38] & b[0])^(a[37] & b[1])^(a[36] & b[2])^(a[35] & b[3])^(a[34] & b[4])^(a[33] & b[5])^(a[32] & b[6])^(a[31] & b[7])^(a[30] & b[8])^(a[29] & b[9])^(a[28] & b[10])^(a[27] & b[11])^(a[26] & b[12])^(a[25] & b[13])^(a[24] & b[14])^(a[23] & b[15])^(a[22] & b[16])^(a[21] & b[17])^(a[20] & b[18])^(a[19] & b[19])^(a[18] & b[20])^(a[17] & b[21])^(a[16] & b[22])^(a[15] & b[23])^(a[14] & b[24])^(a[13] & b[25])^(a[12] & b[26])^(a[11] & b[27])^(a[10] & b[28])^(a[9] & b[29])^(a[8] & b[30])^(a[7] & b[31])^(a[6] & b[32])^(a[5] & b[33])^(a[4] & b[34])^(a[3] & b[35])^(a[2] & b[36])^(a[1] & b[37])^(a[0] & b[38]);
assign y[39] = (a[39] & b[0])^(a[38] & b[1])^(a[37] & b[2])^(a[36] & b[3])^(a[35] & b[4])^(a[34] & b[5])^(a[33] & b[6])^(a[32] & b[7])^(a[31] & b[8])^(a[30] & b[9])^(a[29] & b[10])^(a[28] & b[11])^(a[27] & b[12])^(a[26] & b[13])^(a[25] & b[14])^(a[24] & b[15])^(a[23] & b[16])^(a[22] & b[17])^(a[21] & b[18])^(a[20] & b[19])^(a[19] & b[20])^(a[18] & b[21])^(a[17] & b[22])^(a[16] & b[23])^(a[15] & b[24])^(a[14] & b[25])^(a[13] & b[26])^(a[12] & b[27])^(a[11] & b[28])^(a[10] & b[29])^(a[9] & b[30])^(a[8] & b[31])^(a[7] & b[32])^(a[6] & b[33])^(a[5] & b[34])^(a[4] & b[35])^(a[3] & b[36])^(a[2] & b[37])^(a[1] & b[38])^(a[0] & b[39]);
assign y[40] = (a[40] & b[0])^(a[39] & b[1])^(a[38] & b[2])^(a[37] & b[3])^(a[36] & b[4])^(a[35] & b[5])^(a[34] & b[6])^(a[33] & b[7])^(a[32] & b[8])^(a[31] & b[9])^(a[30] & b[10])^(a[29] & b[11])^(a[28] & b[12])^(a[27] & b[13])^(a[26] & b[14])^(a[25] & b[15])^(a[24] & b[16])^(a[23] & b[17])^(a[22] & b[18])^(a[21] & b[19])^(a[20] & b[20])^(a[19] & b[21])^(a[18] & b[22])^(a[17] & b[23])^(a[16] & b[24])^(a[15] & b[25])^(a[14] & b[26])^(a[13] & b[27])^(a[12] & b[28])^(a[11] & b[29])^(a[10] & b[30])^(a[9] & b[31])^(a[8] & b[32])^(a[7] & b[33])^(a[6] & b[34])^(a[5] & b[35])^(a[4] & b[36])^(a[3] & b[37])^(a[2] & b[38])^(a[1] & b[39])^(a[0] & b[40]);
assign y[41] = (a[41] & b[0])^(a[40] & b[1])^(a[39] & b[2])^(a[38] & b[3])^(a[37] & b[4])^(a[36] & b[5])^(a[35] & b[6])^(a[34] & b[7])^(a[33] & b[8])^(a[32] & b[9])^(a[31] & b[10])^(a[30] & b[11])^(a[29] & b[12])^(a[28] & b[13])^(a[27] & b[14])^(a[26] & b[15])^(a[25] & b[16])^(a[24] & b[17])^(a[23] & b[18])^(a[22] & b[19])^(a[21] & b[20])^(a[20] & b[21])^(a[19] & b[22])^(a[18] & b[23])^(a[17] & b[24])^(a[16] & b[25])^(a[15] & b[26])^(a[14] & b[27])^(a[13] & b[28])^(a[12] & b[29])^(a[11] & b[30])^(a[10] & b[31])^(a[9] & b[32])^(a[8] & b[33])^(a[7] & b[34])^(a[6] & b[35])^(a[5] & b[36])^(a[4] & b[37])^(a[3] & b[38])^(a[2] & b[39])^(a[1] & b[40])^(a[0] & b[41]);
assign y[42] = (a[42] & b[0])^(a[41] & b[1])^(a[40] & b[2])^(a[39] & b[3])^(a[38] & b[4])^(a[37] & b[5])^(a[36] & b[6])^(a[35] & b[7])^(a[34] & b[8])^(a[33] & b[9])^(a[32] & b[10])^(a[31] & b[11])^(a[30] & b[12])^(a[29] & b[13])^(a[28] & b[14])^(a[27] & b[15])^(a[26] & b[16])^(a[25] & b[17])^(a[24] & b[18])^(a[23] & b[19])^(a[22] & b[20])^(a[21] & b[21])^(a[20] & b[22])^(a[19] & b[23])^(a[18] & b[24])^(a[17] & b[25])^(a[16] & b[26])^(a[15] & b[27])^(a[14] & b[28])^(a[13] & b[29])^(a[12] & b[30])^(a[11] & b[31])^(a[10] & b[32])^(a[9] & b[33])^(a[8] & b[34])^(a[7] & b[35])^(a[6] & b[36])^(a[5] & b[37])^(a[4] & b[38])^(a[3] & b[39])^(a[2] & b[40])^(a[1] & b[41])^(a[0] & b[42]);
assign y[43] = (a[43] & b[0])^(a[42] & b[1])^(a[41] & b[2])^(a[40] & b[3])^(a[39] & b[4])^(a[38] & b[5])^(a[37] & b[6])^(a[36] & b[7])^(a[35] & b[8])^(a[34] & b[9])^(a[33] & b[10])^(a[32] & b[11])^(a[31] & b[12])^(a[30] & b[13])^(a[29] & b[14])^(a[28] & b[15])^(a[27] & b[16])^(a[26] & b[17])^(a[25] & b[18])^(a[24] & b[19])^(a[23] & b[20])^(a[22] & b[21])^(a[21] & b[22])^(a[20] & b[23])^(a[19] & b[24])^(a[18] & b[25])^(a[17] & b[26])^(a[16] & b[27])^(a[15] & b[28])^(a[14] & b[29])^(a[13] & b[30])^(a[12] & b[31])^(a[11] & b[32])^(a[10] & b[33])^(a[9] & b[34])^(a[8] & b[35])^(a[7] & b[36])^(a[6] & b[37])^(a[5] & b[38])^(a[4] & b[39])^(a[3] & b[40])^(a[2] & b[41])^(a[1] & b[42])^(a[0] & b[43]);
assign y[44] = (a[44] & b[0])^(a[43] & b[1])^(a[42] & b[2])^(a[41] & b[3])^(a[40] & b[4])^(a[39] & b[5])^(a[38] & b[6])^(a[37] & b[7])^(a[36] & b[8])^(a[35] & b[9])^(a[34] & b[10])^(a[33] & b[11])^(a[32] & b[12])^(a[31] & b[13])^(a[30] & b[14])^(a[29] & b[15])^(a[28] & b[16])^(a[27] & b[17])^(a[26] & b[18])^(a[25] & b[19])^(a[24] & b[20])^(a[23] & b[21])^(a[22] & b[22])^(a[21] & b[23])^(a[20] & b[24])^(a[19] & b[25])^(a[18] & b[26])^(a[17] & b[27])^(a[16] & b[28])^(a[15] & b[29])^(a[14] & b[30])^(a[13] & b[31])^(a[12] & b[32])^(a[11] & b[33])^(a[10] & b[34])^(a[9] & b[35])^(a[8] & b[36])^(a[7] & b[37])^(a[6] & b[38])^(a[5] & b[39])^(a[4] & b[40])^(a[3] & b[41])^(a[2] & b[42])^(a[1] & b[43])^(a[0] & b[44]);
assign y[45] = (a[45] & b[0])^(a[44] & b[1])^(a[43] & b[2])^(a[42] & b[3])^(a[41] & b[4])^(a[40] & b[5])^(a[39] & b[6])^(a[38] & b[7])^(a[37] & b[8])^(a[36] & b[9])^(a[35] & b[10])^(a[34] & b[11])^(a[33] & b[12])^(a[32] & b[13])^(a[31] & b[14])^(a[30] & b[15])^(a[29] & b[16])^(a[28] & b[17])^(a[27] & b[18])^(a[26] & b[19])^(a[25] & b[20])^(a[24] & b[21])^(a[23] & b[22])^(a[22] & b[23])^(a[21] & b[24])^(a[20] & b[25])^(a[19] & b[26])^(a[18] & b[27])^(a[17] & b[28])^(a[16] & b[29])^(a[15] & b[30])^(a[14] & b[31])^(a[13] & b[32])^(a[12] & b[33])^(a[11] & b[34])^(a[10] & b[35])^(a[9] & b[36])^(a[8] & b[37])^(a[7] & b[38])^(a[6] & b[39])^(a[5] & b[40])^(a[4] & b[41])^(a[3] & b[42])^(a[2] & b[43])^(a[1] & b[44])^(a[0] & b[45]);
assign y[46] = (a[46] & b[0])^(a[45] & b[1])^(a[44] & b[2])^(a[43] & b[3])^(a[42] & b[4])^(a[41] & b[5])^(a[40] & b[6])^(a[39] & b[7])^(a[38] & b[8])^(a[37] & b[9])^(a[36] & b[10])^(a[35] & b[11])^(a[34] & b[12])^(a[33] & b[13])^(a[32] & b[14])^(a[31] & b[15])^(a[30] & b[16])^(a[29] & b[17])^(a[28] & b[18])^(a[27] & b[19])^(a[26] & b[20])^(a[25] & b[21])^(a[24] & b[22])^(a[23] & b[23])^(a[22] & b[24])^(a[21] & b[25])^(a[20] & b[26])^(a[19] & b[27])^(a[18] & b[28])^(a[17] & b[29])^(a[16] & b[30])^(a[15] & b[31])^(a[14] & b[32])^(a[13] & b[33])^(a[12] & b[34])^(a[11] & b[35])^(a[10] & b[36])^(a[9] & b[37])^(a[8] & b[38])^(a[7] & b[39])^(a[6] & b[40])^(a[5] & b[41])^(a[4] & b[42])^(a[3] & b[43])^(a[2] & b[44])^(a[1] & b[45])^(a[0] & b[46]);
assign y[47] = (a[47] & b[0])^(a[46] & b[1])^(a[45] & b[2])^(a[44] & b[3])^(a[43] & b[4])^(a[42] & b[5])^(a[41] & b[6])^(a[40] & b[7])^(a[39] & b[8])^(a[38] & b[9])^(a[37] & b[10])^(a[36] & b[11])^(a[35] & b[12])^(a[34] & b[13])^(a[33] & b[14])^(a[32] & b[15])^(a[31] & b[16])^(a[30] & b[17])^(a[29] & b[18])^(a[28] & b[19])^(a[27] & b[20])^(a[26] & b[21])^(a[25] & b[22])^(a[24] & b[23])^(a[23] & b[24])^(a[22] & b[25])^(a[21] & b[26])^(a[20] & b[27])^(a[19] & b[28])^(a[18] & b[29])^(a[17] & b[30])^(a[16] & b[31])^(a[15] & b[32])^(a[14] & b[33])^(a[13] & b[34])^(a[12] & b[35])^(a[11] & b[36])^(a[10] & b[37])^(a[9] & b[38])^(a[8] & b[39])^(a[7] & b[40])^(a[6] & b[41])^(a[5] & b[42])^(a[4] & b[43])^(a[3] & b[44])^(a[2] & b[45])^(a[1] & b[46])^(a[0] & b[47]);
assign y[48] = (a[48] & b[0])^(a[47] & b[1])^(a[46] & b[2])^(a[45] & b[3])^(a[44] & b[4])^(a[43] & b[5])^(a[42] & b[6])^(a[41] & b[7])^(a[40] & b[8])^(a[39] & b[9])^(a[38] & b[10])^(a[37] & b[11])^(a[36] & b[12])^(a[35] & b[13])^(a[34] & b[14])^(a[33] & b[15])^(a[32] & b[16])^(a[31] & b[17])^(a[30] & b[18])^(a[29] & b[19])^(a[28] & b[20])^(a[27] & b[21])^(a[26] & b[22])^(a[25] & b[23])^(a[24] & b[24])^(a[23] & b[25])^(a[22] & b[26])^(a[21] & b[27])^(a[20] & b[28])^(a[19] & b[29])^(a[18] & b[30])^(a[17] & b[31])^(a[16] & b[32])^(a[15] & b[33])^(a[14] & b[34])^(a[13] & b[35])^(a[12] & b[36])^(a[11] & b[37])^(a[10] & b[38])^(a[9] & b[39])^(a[8] & b[40])^(a[7] & b[41])^(a[6] & b[42])^(a[5] & b[43])^(a[4] & b[44])^(a[3] & b[45])^(a[2] & b[46])^(a[1] & b[47])^(a[0] & b[48]);
assign y[49] = (a[49] & b[0])^(a[48] & b[1])^(a[47] & b[2])^(a[46] & b[3])^(a[45] & b[4])^(a[44] & b[5])^(a[43] & b[6])^(a[42] & b[7])^(a[41] & b[8])^(a[40] & b[9])^(a[39] & b[10])^(a[38] & b[11])^(a[37] & b[12])^(a[36] & b[13])^(a[35] & b[14])^(a[34] & b[15])^(a[33] & b[16])^(a[32] & b[17])^(a[31] & b[18])^(a[30] & b[19])^(a[29] & b[20])^(a[28] & b[21])^(a[27] & b[22])^(a[26] & b[23])^(a[25] & b[24])^(a[24] & b[25])^(a[23] & b[26])^(a[22] & b[27])^(a[21] & b[28])^(a[20] & b[29])^(a[19] & b[30])^(a[18] & b[31])^(a[17] & b[32])^(a[16] & b[33])^(a[15] & b[34])^(a[14] & b[35])^(a[13] & b[36])^(a[12] & b[37])^(a[11] & b[38])^(a[10] & b[39])^(a[9] & b[40])^(a[8] & b[41])^(a[7] & b[42])^(a[6] & b[43])^(a[5] & b[44])^(a[4] & b[45])^(a[3] & b[46])^(a[2] & b[47])^(a[1] & b[48])^(a[0] & b[49]);
assign y[50] = (a[50] & b[0])^(a[49] & b[1])^(a[48] & b[2])^(a[47] & b[3])^(a[46] & b[4])^(a[45] & b[5])^(a[44] & b[6])^(a[43] & b[7])^(a[42] & b[8])^(a[41] & b[9])^(a[40] & b[10])^(a[39] & b[11])^(a[38] & b[12])^(a[37] & b[13])^(a[36] & b[14])^(a[35] & b[15])^(a[34] & b[16])^(a[33] & b[17])^(a[32] & b[18])^(a[31] & b[19])^(a[30] & b[20])^(a[29] & b[21])^(a[28] & b[22])^(a[27] & b[23])^(a[26] & b[24])^(a[25] & b[25])^(a[24] & b[26])^(a[23] & b[27])^(a[22] & b[28])^(a[21] & b[29])^(a[20] & b[30])^(a[19] & b[31])^(a[18] & b[32])^(a[17] & b[33])^(a[16] & b[34])^(a[15] & b[35])^(a[14] & b[36])^(a[13] & b[37])^(a[12] & b[38])^(a[11] & b[39])^(a[10] & b[40])^(a[9] & b[41])^(a[8] & b[42])^(a[7] & b[43])^(a[6] & b[44])^(a[5] & b[45])^(a[4] & b[46])^(a[3] & b[47])^(a[2] & b[48])^(a[1] & b[49])^(a[0] & b[50]);
assign y[51] = (a[51] & b[0])^(a[50] & b[1])^(a[49] & b[2])^(a[48] & b[3])^(a[47] & b[4])^(a[46] & b[5])^(a[45] & b[6])^(a[44] & b[7])^(a[43] & b[8])^(a[42] & b[9])^(a[41] & b[10])^(a[40] & b[11])^(a[39] & b[12])^(a[38] & b[13])^(a[37] & b[14])^(a[36] & b[15])^(a[35] & b[16])^(a[34] & b[17])^(a[33] & b[18])^(a[32] & b[19])^(a[31] & b[20])^(a[30] & b[21])^(a[29] & b[22])^(a[28] & b[23])^(a[27] & b[24])^(a[26] & b[25])^(a[25] & b[26])^(a[24] & b[27])^(a[23] & b[28])^(a[22] & b[29])^(a[21] & b[30])^(a[20] & b[31])^(a[19] & b[32])^(a[18] & b[33])^(a[17] & b[34])^(a[16] & b[35])^(a[15] & b[36])^(a[14] & b[37])^(a[13] & b[38])^(a[12] & b[39])^(a[11] & b[40])^(a[10] & b[41])^(a[9] & b[42])^(a[8] & b[43])^(a[7] & b[44])^(a[6] & b[45])^(a[5] & b[46])^(a[4] & b[47])^(a[3] & b[48])^(a[2] & b[49])^(a[1] & b[50])^(a[0] & b[51]);
assign y[52] = (a[52] & b[0])^(a[51] & b[1])^(a[50] & b[2])^(a[49] & b[3])^(a[48] & b[4])^(a[47] & b[5])^(a[46] & b[6])^(a[45] & b[7])^(a[44] & b[8])^(a[43] & b[9])^(a[42] & b[10])^(a[41] & b[11])^(a[40] & b[12])^(a[39] & b[13])^(a[38] & b[14])^(a[37] & b[15])^(a[36] & b[16])^(a[35] & b[17])^(a[34] & b[18])^(a[33] & b[19])^(a[32] & b[20])^(a[31] & b[21])^(a[30] & b[22])^(a[29] & b[23])^(a[28] & b[24])^(a[27] & b[25])^(a[26] & b[26])^(a[25] & b[27])^(a[24] & b[28])^(a[23] & b[29])^(a[22] & b[30])^(a[21] & b[31])^(a[20] & b[32])^(a[19] & b[33])^(a[18] & b[34])^(a[17] & b[35])^(a[16] & b[36])^(a[15] & b[37])^(a[14] & b[38])^(a[13] & b[39])^(a[12] & b[40])^(a[11] & b[41])^(a[10] & b[42])^(a[9] & b[43])^(a[8] & b[44])^(a[7] & b[45])^(a[6] & b[46])^(a[5] & b[47])^(a[4] & b[48])^(a[3] & b[49])^(a[2] & b[50])^(a[1] & b[51])^(a[0] & b[52]);
assign y[53] = (a[53] & b[0])^(a[52] & b[1])^(a[51] & b[2])^(a[50] & b[3])^(a[49] & b[4])^(a[48] & b[5])^(a[47] & b[6])^(a[46] & b[7])^(a[45] & b[8])^(a[44] & b[9])^(a[43] & b[10])^(a[42] & b[11])^(a[41] & b[12])^(a[40] & b[13])^(a[39] & b[14])^(a[38] & b[15])^(a[37] & b[16])^(a[36] & b[17])^(a[35] & b[18])^(a[34] & b[19])^(a[33] & b[20])^(a[32] & b[21])^(a[31] & b[22])^(a[30] & b[23])^(a[29] & b[24])^(a[28] & b[25])^(a[27] & b[26])^(a[26] & b[27])^(a[25] & b[28])^(a[24] & b[29])^(a[23] & b[30])^(a[22] & b[31])^(a[21] & b[32])^(a[20] & b[33])^(a[19] & b[34])^(a[18] & b[35])^(a[17] & b[36])^(a[16] & b[37])^(a[15] & b[38])^(a[14] & b[39])^(a[13] & b[40])^(a[12] & b[41])^(a[11] & b[42])^(a[10] & b[43])^(a[9] & b[44])^(a[8] & b[45])^(a[7] & b[46])^(a[6] & b[47])^(a[5] & b[48])^(a[4] & b[49])^(a[3] & b[50])^(a[2] & b[51])^(a[1] & b[52])^(a[0] & b[53]);
assign y[54] = (a[54] & b[0])^(a[53] & b[1])^(a[52] & b[2])^(a[51] & b[3])^(a[50] & b[4])^(a[49] & b[5])^(a[48] & b[6])^(a[47] & b[7])^(a[46] & b[8])^(a[45] & b[9])^(a[44] & b[10])^(a[43] & b[11])^(a[42] & b[12])^(a[41] & b[13])^(a[40] & b[14])^(a[39] & b[15])^(a[38] & b[16])^(a[37] & b[17])^(a[36] & b[18])^(a[35] & b[19])^(a[34] & b[20])^(a[33] & b[21])^(a[32] & b[22])^(a[31] & b[23])^(a[30] & b[24])^(a[29] & b[25])^(a[28] & b[26])^(a[27] & b[27])^(a[26] & b[28])^(a[25] & b[29])^(a[24] & b[30])^(a[23] & b[31])^(a[22] & b[32])^(a[21] & b[33])^(a[20] & b[34])^(a[19] & b[35])^(a[18] & b[36])^(a[17] & b[37])^(a[16] & b[38])^(a[15] & b[39])^(a[14] & b[40])^(a[13] & b[41])^(a[12] & b[42])^(a[11] & b[43])^(a[10] & b[44])^(a[9] & b[45])^(a[8] & b[46])^(a[7] & b[47])^(a[6] & b[48])^(a[5] & b[49])^(a[4] & b[50])^(a[3] & b[51])^(a[2] & b[52])^(a[1] & b[53])^(a[0] & b[54]);
assign y[55] = (a[55] & b[0])^(a[54] & b[1])^(a[53] & b[2])^(a[52] & b[3])^(a[51] & b[4])^(a[50] & b[5])^(a[49] & b[6])^(a[48] & b[7])^(a[47] & b[8])^(a[46] & b[9])^(a[45] & b[10])^(a[44] & b[11])^(a[43] & b[12])^(a[42] & b[13])^(a[41] & b[14])^(a[40] & b[15])^(a[39] & b[16])^(a[38] & b[17])^(a[37] & b[18])^(a[36] & b[19])^(a[35] & b[20])^(a[34] & b[21])^(a[33] & b[22])^(a[32] & b[23])^(a[31] & b[24])^(a[30] & b[25])^(a[29] & b[26])^(a[28] & b[27])^(a[27] & b[28])^(a[26] & b[29])^(a[25] & b[30])^(a[24] & b[31])^(a[23] & b[32])^(a[22] & b[33])^(a[21] & b[34])^(a[20] & b[35])^(a[19] & b[36])^(a[18] & b[37])^(a[17] & b[38])^(a[16] & b[39])^(a[15] & b[40])^(a[14] & b[41])^(a[13] & b[42])^(a[12] & b[43])^(a[11] & b[44])^(a[10] & b[45])^(a[9] & b[46])^(a[8] & b[47])^(a[7] & b[48])^(a[6] & b[49])^(a[5] & b[50])^(a[4] & b[51])^(a[3] & b[52])^(a[2] & b[53])^(a[1] & b[54])^(a[0] & b[55]);
assign y[56] = (a[56] & b[0])^(a[55] & b[1])^(a[54] & b[2])^(a[53] & b[3])^(a[52] & b[4])^(a[51] & b[5])^(a[50] & b[6])^(a[49] & b[7])^(a[48] & b[8])^(a[47] & b[9])^(a[46] & b[10])^(a[45] & b[11])^(a[44] & b[12])^(a[43] & b[13])^(a[42] & b[14])^(a[41] & b[15])^(a[40] & b[16])^(a[39] & b[17])^(a[38] & b[18])^(a[37] & b[19])^(a[36] & b[20])^(a[35] & b[21])^(a[34] & b[22])^(a[33] & b[23])^(a[32] & b[24])^(a[31] & b[25])^(a[30] & b[26])^(a[29] & b[27])^(a[28] & b[28])^(a[27] & b[29])^(a[26] & b[30])^(a[25] & b[31])^(a[24] & b[32])^(a[23] & b[33])^(a[22] & b[34])^(a[21] & b[35])^(a[20] & b[36])^(a[19] & b[37])^(a[18] & b[38])^(a[17] & b[39])^(a[16] & b[40])^(a[15] & b[41])^(a[14] & b[42])^(a[13] & b[43])^(a[12] & b[44])^(a[11] & b[45])^(a[10] & b[46])^(a[9] & b[47])^(a[8] & b[48])^(a[7] & b[49])^(a[6] & b[50])^(a[5] & b[51])^(a[4] & b[52])^(a[3] & b[53])^(a[2] & b[54])^(a[1] & b[55])^(a[0] & b[56]);
assign y[57] = (a[57] & b[0])^(a[56] & b[1])^(a[55] & b[2])^(a[54] & b[3])^(a[53] & b[4])^(a[52] & b[5])^(a[51] & b[6])^(a[50] & b[7])^(a[49] & b[8])^(a[48] & b[9])^(a[47] & b[10])^(a[46] & b[11])^(a[45] & b[12])^(a[44] & b[13])^(a[43] & b[14])^(a[42] & b[15])^(a[41] & b[16])^(a[40] & b[17])^(a[39] & b[18])^(a[38] & b[19])^(a[37] & b[20])^(a[36] & b[21])^(a[35] & b[22])^(a[34] & b[23])^(a[33] & b[24])^(a[32] & b[25])^(a[31] & b[26])^(a[30] & b[27])^(a[29] & b[28])^(a[28] & b[29])^(a[27] & b[30])^(a[26] & b[31])^(a[25] & b[32])^(a[24] & b[33])^(a[23] & b[34])^(a[22] & b[35])^(a[21] & b[36])^(a[20] & b[37])^(a[19] & b[38])^(a[18] & b[39])^(a[17] & b[40])^(a[16] & b[41])^(a[15] & b[42])^(a[14] & b[43])^(a[13] & b[44])^(a[12] & b[45])^(a[11] & b[46])^(a[10] & b[47])^(a[9] & b[48])^(a[8] & b[49])^(a[7] & b[50])^(a[6] & b[51])^(a[5] & b[52])^(a[4] & b[53])^(a[3] & b[54])^(a[2] & b[55])^(a[1] & b[56])^(a[0] & b[57]);
assign y[58] = (a[58] & b[0])^(a[57] & b[1])^(a[56] & b[2])^(a[55] & b[3])^(a[54] & b[4])^(a[53] & b[5])^(a[52] & b[6])^(a[51] & b[7])^(a[50] & b[8])^(a[49] & b[9])^(a[48] & b[10])^(a[47] & b[11])^(a[46] & b[12])^(a[45] & b[13])^(a[44] & b[14])^(a[43] & b[15])^(a[42] & b[16])^(a[41] & b[17])^(a[40] & b[18])^(a[39] & b[19])^(a[38] & b[20])^(a[37] & b[21])^(a[36] & b[22])^(a[35] & b[23])^(a[34] & b[24])^(a[33] & b[25])^(a[32] & b[26])^(a[31] & b[27])^(a[30] & b[28])^(a[29] & b[29])^(a[28] & b[30])^(a[27] & b[31])^(a[26] & b[32])^(a[25] & b[33])^(a[24] & b[34])^(a[23] & b[35])^(a[22] & b[36])^(a[21] & b[37])^(a[20] & b[38])^(a[19] & b[39])^(a[18] & b[40])^(a[17] & b[41])^(a[16] & b[42])^(a[15] & b[43])^(a[14] & b[44])^(a[13] & b[45])^(a[12] & b[46])^(a[11] & b[47])^(a[10] & b[48])^(a[9] & b[49])^(a[8] & b[50])^(a[7] & b[51])^(a[6] & b[52])^(a[5] & b[53])^(a[4] & b[54])^(a[3] & b[55])^(a[2] & b[56])^(a[1] & b[57])^(a[0] & b[58]);
assign y[59] = (a[59] & b[0])^(a[58] & b[1])^(a[57] & b[2])^(a[56] & b[3])^(a[55] & b[4])^(a[54] & b[5])^(a[53] & b[6])^(a[52] & b[7])^(a[51] & b[8])^(a[50] & b[9])^(a[49] & b[10])^(a[48] & b[11])^(a[47] & b[12])^(a[46] & b[13])^(a[45] & b[14])^(a[44] & b[15])^(a[43] & b[16])^(a[42] & b[17])^(a[41] & b[18])^(a[40] & b[19])^(a[39] & b[20])^(a[38] & b[21])^(a[37] & b[22])^(a[36] & b[23])^(a[35] & b[24])^(a[34] & b[25])^(a[33] & b[26])^(a[32] & b[27])^(a[31] & b[28])^(a[30] & b[29])^(a[29] & b[30])^(a[28] & b[31])^(a[27] & b[32])^(a[26] & b[33])^(a[25] & b[34])^(a[24] & b[35])^(a[23] & b[36])^(a[22] & b[37])^(a[21] & b[38])^(a[20] & b[39])^(a[19] & b[40])^(a[18] & b[41])^(a[17] & b[42])^(a[16] & b[43])^(a[15] & b[44])^(a[14] & b[45])^(a[13] & b[46])^(a[12] & b[47])^(a[11] & b[48])^(a[10] & b[49])^(a[9] & b[50])^(a[8] & b[51])^(a[7] & b[52])^(a[6] & b[53])^(a[5] & b[54])^(a[4] & b[55])^(a[3] & b[56])^(a[2] & b[57])^(a[1] & b[58])^(a[0] & b[59]);
assign y[60] = (a[60] & b[0])^(a[59] & b[1])^(a[58] & b[2])^(a[57] & b[3])^(a[56] & b[4])^(a[55] & b[5])^(a[54] & b[6])^(a[53] & b[7])^(a[52] & b[8])^(a[51] & b[9])^(a[50] & b[10])^(a[49] & b[11])^(a[48] & b[12])^(a[47] & b[13])^(a[46] & b[14])^(a[45] & b[15])^(a[44] & b[16])^(a[43] & b[17])^(a[42] & b[18])^(a[41] & b[19])^(a[40] & b[20])^(a[39] & b[21])^(a[38] & b[22])^(a[37] & b[23])^(a[36] & b[24])^(a[35] & b[25])^(a[34] & b[26])^(a[33] & b[27])^(a[32] & b[28])^(a[31] & b[29])^(a[30] & b[30])^(a[29] & b[31])^(a[28] & b[32])^(a[27] & b[33])^(a[26] & b[34])^(a[25] & b[35])^(a[24] & b[36])^(a[23] & b[37])^(a[22] & b[38])^(a[21] & b[39])^(a[20] & b[40])^(a[19] & b[41])^(a[18] & b[42])^(a[17] & b[43])^(a[16] & b[44])^(a[15] & b[45])^(a[14] & b[46])^(a[13] & b[47])^(a[12] & b[48])^(a[11] & b[49])^(a[10] & b[50])^(a[9] & b[51])^(a[8] & b[52])^(a[7] & b[53])^(a[6] & b[54])^(a[5] & b[55])^(a[4] & b[56])^(a[3] & b[57])^(a[2] & b[58])^(a[1] & b[59])^(a[0] & b[60]);
assign y[61] = (a[61] & b[0])^(a[60] & b[1])^(a[59] & b[2])^(a[58] & b[3])^(a[57] & b[4])^(a[56] & b[5])^(a[55] & b[6])^(a[54] & b[7])^(a[53] & b[8])^(a[52] & b[9])^(a[51] & b[10])^(a[50] & b[11])^(a[49] & b[12])^(a[48] & b[13])^(a[47] & b[14])^(a[46] & b[15])^(a[45] & b[16])^(a[44] & b[17])^(a[43] & b[18])^(a[42] & b[19])^(a[41] & b[20])^(a[40] & b[21])^(a[39] & b[22])^(a[38] & b[23])^(a[37] & b[24])^(a[36] & b[25])^(a[35] & b[26])^(a[34] & b[27])^(a[33] & b[28])^(a[32] & b[29])^(a[31] & b[30])^(a[30] & b[31])^(a[29] & b[32])^(a[28] & b[33])^(a[27] & b[34])^(a[26] & b[35])^(a[25] & b[36])^(a[24] & b[37])^(a[23] & b[38])^(a[22] & b[39])^(a[21] & b[40])^(a[20] & b[41])^(a[19] & b[42])^(a[18] & b[43])^(a[17] & b[44])^(a[16] & b[45])^(a[15] & b[46])^(a[14] & b[47])^(a[13] & b[48])^(a[12] & b[49])^(a[11] & b[50])^(a[10] & b[51])^(a[9] & b[52])^(a[8] & b[53])^(a[7] & b[54])^(a[6] & b[55])^(a[5] & b[56])^(a[4] & b[57])^(a[3] & b[58])^(a[2] & b[59])^(a[1] & b[60])^(a[0] & b[61]);
assign y[62] = (a[62] & b[0])^(a[61] & b[1])^(a[60] & b[2])^(a[59] & b[3])^(a[58] & b[4])^(a[57] & b[5])^(a[56] & b[6])^(a[55] & b[7])^(a[54] & b[8])^(a[53] & b[9])^(a[52] & b[10])^(a[51] & b[11])^(a[50] & b[12])^(a[49] & b[13])^(a[48] & b[14])^(a[47] & b[15])^(a[46] & b[16])^(a[45] & b[17])^(a[44] & b[18])^(a[43] & b[19])^(a[42] & b[20])^(a[41] & b[21])^(a[40] & b[22])^(a[39] & b[23])^(a[38] & b[24])^(a[37] & b[25])^(a[36] & b[26])^(a[35] & b[27])^(a[34] & b[28])^(a[33] & b[29])^(a[32] & b[30])^(a[31] & b[31])^(a[30] & b[32])^(a[29] & b[33])^(a[28] & b[34])^(a[27] & b[35])^(a[26] & b[36])^(a[25] & b[37])^(a[24] & b[38])^(a[23] & b[39])^(a[22] & b[40])^(a[21] & b[41])^(a[20] & b[42])^(a[19] & b[43])^(a[18] & b[44])^(a[17] & b[45])^(a[16] & b[46])^(a[15] & b[47])^(a[14] & b[48])^(a[13] & b[49])^(a[12] & b[50])^(a[11] & b[51])^(a[10] & b[52])^(a[9] & b[53])^(a[8] & b[54])^(a[7] & b[55])^(a[6] & b[56])^(a[5] & b[57])^(a[4] & b[58])^(a[3] & b[59])^(a[2] & b[60])^(a[1] & b[61])^(a[0] & b[62]);
assign y[63] = (a[63] & b[0])^(a[62] & b[1])^(a[61] & b[2])^(a[60] & b[3])^(a[59] & b[4])^(a[58] & b[5])^(a[57] & b[6])^(a[56] & b[7])^(a[55] & b[8])^(a[54] & b[9])^(a[53] & b[10])^(a[52] & b[11])^(a[51] & b[12])^(a[50] & b[13])^(a[49] & b[14])^(a[48] & b[15])^(a[47] & b[16])^(a[46] & b[17])^(a[45] & b[18])^(a[44] & b[19])^(a[43] & b[20])^(a[42] & b[21])^(a[41] & b[22])^(a[40] & b[23])^(a[39] & b[24])^(a[38] & b[25])^(a[37] & b[26])^(a[36] & b[27])^(a[35] & b[28])^(a[34] & b[29])^(a[33] & b[30])^(a[32] & b[31])^(a[31] & b[32])^(a[30] & b[33])^(a[29] & b[34])^(a[28] & b[35])^(a[27] & b[36])^(a[26] & b[37])^(a[25] & b[38])^(a[24] & b[39])^(a[23] & b[40])^(a[22] & b[41])^(a[21] & b[42])^(a[20] & b[43])^(a[19] & b[44])^(a[18] & b[45])^(a[17] & b[46])^(a[16] & b[47])^(a[15] & b[48])^(a[14] & b[49])^(a[13] & b[50])^(a[12] & b[51])^(a[11] & b[52])^(a[10] & b[53])^(a[9] & b[54])^(a[8] & b[55])^(a[7] & b[56])^(a[6] & b[57])^(a[5] & b[58])^(a[4] & b[59])^(a[3] & b[60])^(a[2] & b[61])^(a[1] & b[62])^(a[0] & b[63]);
assign y[64] = (a[64] & b[0])^(a[63] & b[1])^(a[62] & b[2])^(a[61] & b[3])^(a[60] & b[4])^(a[59] & b[5])^(a[58] & b[6])^(a[57] & b[7])^(a[56] & b[8])^(a[55] & b[9])^(a[54] & b[10])^(a[53] & b[11])^(a[52] & b[12])^(a[51] & b[13])^(a[50] & b[14])^(a[49] & b[15])^(a[48] & b[16])^(a[47] & b[17])^(a[46] & b[18])^(a[45] & b[19])^(a[44] & b[20])^(a[43] & b[21])^(a[42] & b[22])^(a[41] & b[23])^(a[40] & b[24])^(a[39] & b[25])^(a[38] & b[26])^(a[37] & b[27])^(a[36] & b[28])^(a[35] & b[29])^(a[34] & b[30])^(a[33] & b[31])^(a[32] & b[32])^(a[31] & b[33])^(a[30] & b[34])^(a[29] & b[35])^(a[28] & b[36])^(a[27] & b[37])^(a[26] & b[38])^(a[25] & b[39])^(a[24] & b[40])^(a[23] & b[41])^(a[22] & b[42])^(a[21] & b[43])^(a[20] & b[44])^(a[19] & b[45])^(a[18] & b[46])^(a[17] & b[47])^(a[16] & b[48])^(a[15] & b[49])^(a[14] & b[50])^(a[13] & b[51])^(a[12] & b[52])^(a[11] & b[53])^(a[10] & b[54])^(a[9] & b[55])^(a[8] & b[56])^(a[7] & b[57])^(a[6] & b[58])^(a[5] & b[59])^(a[4] & b[60])^(a[3] & b[61])^(a[2] & b[62])^(a[1] & b[63])^(a[0] & b[64]);
assign y[65] = (a[65] & b[0])^(a[64] & b[1])^(a[63] & b[2])^(a[62] & b[3])^(a[61] & b[4])^(a[60] & b[5])^(a[59] & b[6])^(a[58] & b[7])^(a[57] & b[8])^(a[56] & b[9])^(a[55] & b[10])^(a[54] & b[11])^(a[53] & b[12])^(a[52] & b[13])^(a[51] & b[14])^(a[50] & b[15])^(a[49] & b[16])^(a[48] & b[17])^(a[47] & b[18])^(a[46] & b[19])^(a[45] & b[20])^(a[44] & b[21])^(a[43] & b[22])^(a[42] & b[23])^(a[41] & b[24])^(a[40] & b[25])^(a[39] & b[26])^(a[38] & b[27])^(a[37] & b[28])^(a[36] & b[29])^(a[35] & b[30])^(a[34] & b[31])^(a[33] & b[32])^(a[32] & b[33])^(a[31] & b[34])^(a[30] & b[35])^(a[29] & b[36])^(a[28] & b[37])^(a[27] & b[38])^(a[26] & b[39])^(a[25] & b[40])^(a[24] & b[41])^(a[23] & b[42])^(a[22] & b[43])^(a[21] & b[44])^(a[20] & b[45])^(a[19] & b[46])^(a[18] & b[47])^(a[17] & b[48])^(a[16] & b[49])^(a[15] & b[50])^(a[14] & b[51])^(a[13] & b[52])^(a[12] & b[53])^(a[11] & b[54])^(a[10] & b[55])^(a[9] & b[56])^(a[8] & b[57])^(a[7] & b[58])^(a[6] & b[59])^(a[5] & b[60])^(a[4] & b[61])^(a[3] & b[62])^(a[2] & b[63])^(a[1] & b[64])^(a[0] & b[65]);
assign y[66] = (a[66] & b[0])^(a[65] & b[1])^(a[64] & b[2])^(a[63] & b[3])^(a[62] & b[4])^(a[61] & b[5])^(a[60] & b[6])^(a[59] & b[7])^(a[58] & b[8])^(a[57] & b[9])^(a[56] & b[10])^(a[55] & b[11])^(a[54] & b[12])^(a[53] & b[13])^(a[52] & b[14])^(a[51] & b[15])^(a[50] & b[16])^(a[49] & b[17])^(a[48] & b[18])^(a[47] & b[19])^(a[46] & b[20])^(a[45] & b[21])^(a[44] & b[22])^(a[43] & b[23])^(a[42] & b[24])^(a[41] & b[25])^(a[40] & b[26])^(a[39] & b[27])^(a[38] & b[28])^(a[37] & b[29])^(a[36] & b[30])^(a[35] & b[31])^(a[34] & b[32])^(a[33] & b[33])^(a[32] & b[34])^(a[31] & b[35])^(a[30] & b[36])^(a[29] & b[37])^(a[28] & b[38])^(a[27] & b[39])^(a[26] & b[40])^(a[25] & b[41])^(a[24] & b[42])^(a[23] & b[43])^(a[22] & b[44])^(a[21] & b[45])^(a[20] & b[46])^(a[19] & b[47])^(a[18] & b[48])^(a[17] & b[49])^(a[16] & b[50])^(a[15] & b[51])^(a[14] & b[52])^(a[13] & b[53])^(a[12] & b[54])^(a[11] & b[55])^(a[10] & b[56])^(a[9] & b[57])^(a[8] & b[58])^(a[7] & b[59])^(a[6] & b[60])^(a[5] & b[61])^(a[4] & b[62])^(a[3] & b[63])^(a[2] & b[64])^(a[1] & b[65])^(a[0] & b[66]);
assign y[67] = (a[67] & b[0])^(a[66] & b[1])^(a[65] & b[2])^(a[64] & b[3])^(a[63] & b[4])^(a[62] & b[5])^(a[61] & b[6])^(a[60] & b[7])^(a[59] & b[8])^(a[58] & b[9])^(a[57] & b[10])^(a[56] & b[11])^(a[55] & b[12])^(a[54] & b[13])^(a[53] & b[14])^(a[52] & b[15])^(a[51] & b[16])^(a[50] & b[17])^(a[49] & b[18])^(a[48] & b[19])^(a[47] & b[20])^(a[46] & b[21])^(a[45] & b[22])^(a[44] & b[23])^(a[43] & b[24])^(a[42] & b[25])^(a[41] & b[26])^(a[40] & b[27])^(a[39] & b[28])^(a[38] & b[29])^(a[37] & b[30])^(a[36] & b[31])^(a[35] & b[32])^(a[34] & b[33])^(a[33] & b[34])^(a[32] & b[35])^(a[31] & b[36])^(a[30] & b[37])^(a[29] & b[38])^(a[28] & b[39])^(a[27] & b[40])^(a[26] & b[41])^(a[25] & b[42])^(a[24] & b[43])^(a[23] & b[44])^(a[22] & b[45])^(a[21] & b[46])^(a[20] & b[47])^(a[19] & b[48])^(a[18] & b[49])^(a[17] & b[50])^(a[16] & b[51])^(a[15] & b[52])^(a[14] & b[53])^(a[13] & b[54])^(a[12] & b[55])^(a[11] & b[56])^(a[10] & b[57])^(a[9] & b[58])^(a[8] & b[59])^(a[7] & b[60])^(a[6] & b[61])^(a[5] & b[62])^(a[4] & b[63])^(a[3] & b[64])^(a[2] & b[65])^(a[1] & b[66])^(a[0] & b[67]);
assign y[68] = (a[68] & b[0])^(a[67] & b[1])^(a[66] & b[2])^(a[65] & b[3])^(a[64] & b[4])^(a[63] & b[5])^(a[62] & b[6])^(a[61] & b[7])^(a[60] & b[8])^(a[59] & b[9])^(a[58] & b[10])^(a[57] & b[11])^(a[56] & b[12])^(a[55] & b[13])^(a[54] & b[14])^(a[53] & b[15])^(a[52] & b[16])^(a[51] & b[17])^(a[50] & b[18])^(a[49] & b[19])^(a[48] & b[20])^(a[47] & b[21])^(a[46] & b[22])^(a[45] & b[23])^(a[44] & b[24])^(a[43] & b[25])^(a[42] & b[26])^(a[41] & b[27])^(a[40] & b[28])^(a[39] & b[29])^(a[38] & b[30])^(a[37] & b[31])^(a[36] & b[32])^(a[35] & b[33])^(a[34] & b[34])^(a[33] & b[35])^(a[32] & b[36])^(a[31] & b[37])^(a[30] & b[38])^(a[29] & b[39])^(a[28] & b[40])^(a[27] & b[41])^(a[26] & b[42])^(a[25] & b[43])^(a[24] & b[44])^(a[23] & b[45])^(a[22] & b[46])^(a[21] & b[47])^(a[20] & b[48])^(a[19] & b[49])^(a[18] & b[50])^(a[17] & b[51])^(a[16] & b[52])^(a[15] & b[53])^(a[14] & b[54])^(a[13] & b[55])^(a[12] & b[56])^(a[11] & b[57])^(a[10] & b[58])^(a[9] & b[59])^(a[8] & b[60])^(a[7] & b[61])^(a[6] & b[62])^(a[5] & b[63])^(a[4] & b[64])^(a[3] & b[65])^(a[2] & b[66])^(a[1] & b[67])^(a[0] & b[68]);
assign y[69] = (a[69] & b[0])^(a[68] & b[1])^(a[67] & b[2])^(a[66] & b[3])^(a[65] & b[4])^(a[64] & b[5])^(a[63] & b[6])^(a[62] & b[7])^(a[61] & b[8])^(a[60] & b[9])^(a[59] & b[10])^(a[58] & b[11])^(a[57] & b[12])^(a[56] & b[13])^(a[55] & b[14])^(a[54] & b[15])^(a[53] & b[16])^(a[52] & b[17])^(a[51] & b[18])^(a[50] & b[19])^(a[49] & b[20])^(a[48] & b[21])^(a[47] & b[22])^(a[46] & b[23])^(a[45] & b[24])^(a[44] & b[25])^(a[43] & b[26])^(a[42] & b[27])^(a[41] & b[28])^(a[40] & b[29])^(a[39] & b[30])^(a[38] & b[31])^(a[37] & b[32])^(a[36] & b[33])^(a[35] & b[34])^(a[34] & b[35])^(a[33] & b[36])^(a[32] & b[37])^(a[31] & b[38])^(a[30] & b[39])^(a[29] & b[40])^(a[28] & b[41])^(a[27] & b[42])^(a[26] & b[43])^(a[25] & b[44])^(a[24] & b[45])^(a[23] & b[46])^(a[22] & b[47])^(a[21] & b[48])^(a[20] & b[49])^(a[19] & b[50])^(a[18] & b[51])^(a[17] & b[52])^(a[16] & b[53])^(a[15] & b[54])^(a[14] & b[55])^(a[13] & b[56])^(a[12] & b[57])^(a[11] & b[58])^(a[10] & b[59])^(a[9] & b[60])^(a[8] & b[61])^(a[7] & b[62])^(a[6] & b[63])^(a[5] & b[64])^(a[4] & b[65])^(a[3] & b[66])^(a[2] & b[67])^(a[1] & b[68])^(a[0] & b[69]);
assign y[70] = (a[70] & b[0])^(a[69] & b[1])^(a[68] & b[2])^(a[67] & b[3])^(a[66] & b[4])^(a[65] & b[5])^(a[64] & b[6])^(a[63] & b[7])^(a[62] & b[8])^(a[61] & b[9])^(a[60] & b[10])^(a[59] & b[11])^(a[58] & b[12])^(a[57] & b[13])^(a[56] & b[14])^(a[55] & b[15])^(a[54] & b[16])^(a[53] & b[17])^(a[52] & b[18])^(a[51] & b[19])^(a[50] & b[20])^(a[49] & b[21])^(a[48] & b[22])^(a[47] & b[23])^(a[46] & b[24])^(a[45] & b[25])^(a[44] & b[26])^(a[43] & b[27])^(a[42] & b[28])^(a[41] & b[29])^(a[40] & b[30])^(a[39] & b[31])^(a[38] & b[32])^(a[37] & b[33])^(a[36] & b[34])^(a[35] & b[35])^(a[34] & b[36])^(a[33] & b[37])^(a[32] & b[38])^(a[31] & b[39])^(a[30] & b[40])^(a[29] & b[41])^(a[28] & b[42])^(a[27] & b[43])^(a[26] & b[44])^(a[25] & b[45])^(a[24] & b[46])^(a[23] & b[47])^(a[22] & b[48])^(a[21] & b[49])^(a[20] & b[50])^(a[19] & b[51])^(a[18] & b[52])^(a[17] & b[53])^(a[16] & b[54])^(a[15] & b[55])^(a[14] & b[56])^(a[13] & b[57])^(a[12] & b[58])^(a[11] & b[59])^(a[10] & b[60])^(a[9] & b[61])^(a[8] & b[62])^(a[7] & b[63])^(a[6] & b[64])^(a[5] & b[65])^(a[4] & b[66])^(a[3] & b[67])^(a[2] & b[68])^(a[1] & b[69])^(a[0] & b[70]);
assign y[71] = (a[71] & b[0])^(a[70] & b[1])^(a[69] & b[2])^(a[68] & b[3])^(a[67] & b[4])^(a[66] & b[5])^(a[65] & b[6])^(a[64] & b[7])^(a[63] & b[8])^(a[62] & b[9])^(a[61] & b[10])^(a[60] & b[11])^(a[59] & b[12])^(a[58] & b[13])^(a[57] & b[14])^(a[56] & b[15])^(a[55] & b[16])^(a[54] & b[17])^(a[53] & b[18])^(a[52] & b[19])^(a[51] & b[20])^(a[50] & b[21])^(a[49] & b[22])^(a[48] & b[23])^(a[47] & b[24])^(a[46] & b[25])^(a[45] & b[26])^(a[44] & b[27])^(a[43] & b[28])^(a[42] & b[29])^(a[41] & b[30])^(a[40] & b[31])^(a[39] & b[32])^(a[38] & b[33])^(a[37] & b[34])^(a[36] & b[35])^(a[35] & b[36])^(a[34] & b[37])^(a[33] & b[38])^(a[32] & b[39])^(a[31] & b[40])^(a[30] & b[41])^(a[29] & b[42])^(a[28] & b[43])^(a[27] & b[44])^(a[26] & b[45])^(a[25] & b[46])^(a[24] & b[47])^(a[23] & b[48])^(a[22] & b[49])^(a[21] & b[50])^(a[20] & b[51])^(a[19] & b[52])^(a[18] & b[53])^(a[17] & b[54])^(a[16] & b[55])^(a[15] & b[56])^(a[14] & b[57])^(a[13] & b[58])^(a[12] & b[59])^(a[11] & b[60])^(a[10] & b[61])^(a[9] & b[62])^(a[8] & b[63])^(a[7] & b[64])^(a[6] & b[65])^(a[5] & b[66])^(a[4] & b[67])^(a[3] & b[68])^(a[2] & b[69])^(a[1] & b[70])^(a[0] & b[71]);
assign y[72] = (a[72] & b[0])^(a[71] & b[1])^(a[70] & b[2])^(a[69] & b[3])^(a[68] & b[4])^(a[67] & b[5])^(a[66] & b[6])^(a[65] & b[7])^(a[64] & b[8])^(a[63] & b[9])^(a[62] & b[10])^(a[61] & b[11])^(a[60] & b[12])^(a[59] & b[13])^(a[58] & b[14])^(a[57] & b[15])^(a[56] & b[16])^(a[55] & b[17])^(a[54] & b[18])^(a[53] & b[19])^(a[52] & b[20])^(a[51] & b[21])^(a[50] & b[22])^(a[49] & b[23])^(a[48] & b[24])^(a[47] & b[25])^(a[46] & b[26])^(a[45] & b[27])^(a[44] & b[28])^(a[43] & b[29])^(a[42] & b[30])^(a[41] & b[31])^(a[40] & b[32])^(a[39] & b[33])^(a[38] & b[34])^(a[37] & b[35])^(a[36] & b[36])^(a[35] & b[37])^(a[34] & b[38])^(a[33] & b[39])^(a[32] & b[40])^(a[31] & b[41])^(a[30] & b[42])^(a[29] & b[43])^(a[28] & b[44])^(a[27] & b[45])^(a[26] & b[46])^(a[25] & b[47])^(a[24] & b[48])^(a[23] & b[49])^(a[22] & b[50])^(a[21] & b[51])^(a[20] & b[52])^(a[19] & b[53])^(a[18] & b[54])^(a[17] & b[55])^(a[16] & b[56])^(a[15] & b[57])^(a[14] & b[58])^(a[13] & b[59])^(a[12] & b[60])^(a[11] & b[61])^(a[10] & b[62])^(a[9] & b[63])^(a[8] & b[64])^(a[7] & b[65])^(a[6] & b[66])^(a[5] & b[67])^(a[4] & b[68])^(a[3] & b[69])^(a[2] & b[70])^(a[1] & b[71])^(a[0] & b[72]);
assign y[73] = (a[73] & b[0])^(a[72] & b[1])^(a[71] & b[2])^(a[70] & b[3])^(a[69] & b[4])^(a[68] & b[5])^(a[67] & b[6])^(a[66] & b[7])^(a[65] & b[8])^(a[64] & b[9])^(a[63] & b[10])^(a[62] & b[11])^(a[61] & b[12])^(a[60] & b[13])^(a[59] & b[14])^(a[58] & b[15])^(a[57] & b[16])^(a[56] & b[17])^(a[55] & b[18])^(a[54] & b[19])^(a[53] & b[20])^(a[52] & b[21])^(a[51] & b[22])^(a[50] & b[23])^(a[49] & b[24])^(a[48] & b[25])^(a[47] & b[26])^(a[46] & b[27])^(a[45] & b[28])^(a[44] & b[29])^(a[43] & b[30])^(a[42] & b[31])^(a[41] & b[32])^(a[40] & b[33])^(a[39] & b[34])^(a[38] & b[35])^(a[37] & b[36])^(a[36] & b[37])^(a[35] & b[38])^(a[34] & b[39])^(a[33] & b[40])^(a[32] & b[41])^(a[31] & b[42])^(a[30] & b[43])^(a[29] & b[44])^(a[28] & b[45])^(a[27] & b[46])^(a[26] & b[47])^(a[25] & b[48])^(a[24] & b[49])^(a[23] & b[50])^(a[22] & b[51])^(a[21] & b[52])^(a[20] & b[53])^(a[19] & b[54])^(a[18] & b[55])^(a[17] & b[56])^(a[16] & b[57])^(a[15] & b[58])^(a[14] & b[59])^(a[13] & b[60])^(a[12] & b[61])^(a[11] & b[62])^(a[10] & b[63])^(a[9] & b[64])^(a[8] & b[65])^(a[7] & b[66])^(a[6] & b[67])^(a[5] & b[68])^(a[4] & b[69])^(a[3] & b[70])^(a[2] & b[71])^(a[1] & b[72])^(a[0] & b[73]);
assign y[74] = (a[74] & b[0])^(a[73] & b[1])^(a[72] & b[2])^(a[71] & b[3])^(a[70] & b[4])^(a[69] & b[5])^(a[68] & b[6])^(a[67] & b[7])^(a[66] & b[8])^(a[65] & b[9])^(a[64] & b[10])^(a[63] & b[11])^(a[62] & b[12])^(a[61] & b[13])^(a[60] & b[14])^(a[59] & b[15])^(a[58] & b[16])^(a[57] & b[17])^(a[56] & b[18])^(a[55] & b[19])^(a[54] & b[20])^(a[53] & b[21])^(a[52] & b[22])^(a[51] & b[23])^(a[50] & b[24])^(a[49] & b[25])^(a[48] & b[26])^(a[47] & b[27])^(a[46] & b[28])^(a[45] & b[29])^(a[44] & b[30])^(a[43] & b[31])^(a[42] & b[32])^(a[41] & b[33])^(a[40] & b[34])^(a[39] & b[35])^(a[38] & b[36])^(a[37] & b[37])^(a[36] & b[38])^(a[35] & b[39])^(a[34] & b[40])^(a[33] & b[41])^(a[32] & b[42])^(a[31] & b[43])^(a[30] & b[44])^(a[29] & b[45])^(a[28] & b[46])^(a[27] & b[47])^(a[26] & b[48])^(a[25] & b[49])^(a[24] & b[50])^(a[23] & b[51])^(a[22] & b[52])^(a[21] & b[53])^(a[20] & b[54])^(a[19] & b[55])^(a[18] & b[56])^(a[17] & b[57])^(a[16] & b[58])^(a[15] & b[59])^(a[14] & b[60])^(a[13] & b[61])^(a[12] & b[62])^(a[11] & b[63])^(a[10] & b[64])^(a[9] & b[65])^(a[8] & b[66])^(a[7] & b[67])^(a[6] & b[68])^(a[5] & b[69])^(a[4] & b[70])^(a[3] & b[71])^(a[2] & b[72])^(a[1] & b[73])^(a[0] & b[74]);
assign y[75] = (a[75] & b[0])^(a[74] & b[1])^(a[73] & b[2])^(a[72] & b[3])^(a[71] & b[4])^(a[70] & b[5])^(a[69] & b[6])^(a[68] & b[7])^(a[67] & b[8])^(a[66] & b[9])^(a[65] & b[10])^(a[64] & b[11])^(a[63] & b[12])^(a[62] & b[13])^(a[61] & b[14])^(a[60] & b[15])^(a[59] & b[16])^(a[58] & b[17])^(a[57] & b[18])^(a[56] & b[19])^(a[55] & b[20])^(a[54] & b[21])^(a[53] & b[22])^(a[52] & b[23])^(a[51] & b[24])^(a[50] & b[25])^(a[49] & b[26])^(a[48] & b[27])^(a[47] & b[28])^(a[46] & b[29])^(a[45] & b[30])^(a[44] & b[31])^(a[43] & b[32])^(a[42] & b[33])^(a[41] & b[34])^(a[40] & b[35])^(a[39] & b[36])^(a[38] & b[37])^(a[37] & b[38])^(a[36] & b[39])^(a[35] & b[40])^(a[34] & b[41])^(a[33] & b[42])^(a[32] & b[43])^(a[31] & b[44])^(a[30] & b[45])^(a[29] & b[46])^(a[28] & b[47])^(a[27] & b[48])^(a[26] & b[49])^(a[25] & b[50])^(a[24] & b[51])^(a[23] & b[52])^(a[22] & b[53])^(a[21] & b[54])^(a[20] & b[55])^(a[19] & b[56])^(a[18] & b[57])^(a[17] & b[58])^(a[16] & b[59])^(a[15] & b[60])^(a[14] & b[61])^(a[13] & b[62])^(a[12] & b[63])^(a[11] & b[64])^(a[10] & b[65])^(a[9] & b[66])^(a[8] & b[67])^(a[7] & b[68])^(a[6] & b[69])^(a[5] & b[70])^(a[4] & b[71])^(a[3] & b[72])^(a[2] & b[73])^(a[1] & b[74])^(a[0] & b[75]);
assign y[76] = (a[76] & b[0])^(a[75] & b[1])^(a[74] & b[2])^(a[73] & b[3])^(a[72] & b[4])^(a[71] & b[5])^(a[70] & b[6])^(a[69] & b[7])^(a[68] & b[8])^(a[67] & b[9])^(a[66] & b[10])^(a[65] & b[11])^(a[64] & b[12])^(a[63] & b[13])^(a[62] & b[14])^(a[61] & b[15])^(a[60] & b[16])^(a[59] & b[17])^(a[58] & b[18])^(a[57] & b[19])^(a[56] & b[20])^(a[55] & b[21])^(a[54] & b[22])^(a[53] & b[23])^(a[52] & b[24])^(a[51] & b[25])^(a[50] & b[26])^(a[49] & b[27])^(a[48] & b[28])^(a[47] & b[29])^(a[46] & b[30])^(a[45] & b[31])^(a[44] & b[32])^(a[43] & b[33])^(a[42] & b[34])^(a[41] & b[35])^(a[40] & b[36])^(a[39] & b[37])^(a[38] & b[38])^(a[37] & b[39])^(a[36] & b[40])^(a[35] & b[41])^(a[34] & b[42])^(a[33] & b[43])^(a[32] & b[44])^(a[31] & b[45])^(a[30] & b[46])^(a[29] & b[47])^(a[28] & b[48])^(a[27] & b[49])^(a[26] & b[50])^(a[25] & b[51])^(a[24] & b[52])^(a[23] & b[53])^(a[22] & b[54])^(a[21] & b[55])^(a[20] & b[56])^(a[19] & b[57])^(a[18] & b[58])^(a[17] & b[59])^(a[16] & b[60])^(a[15] & b[61])^(a[14] & b[62])^(a[13] & b[63])^(a[12] & b[64])^(a[11] & b[65])^(a[10] & b[66])^(a[9] & b[67])^(a[8] & b[68])^(a[7] & b[69])^(a[6] & b[70])^(a[5] & b[71])^(a[4] & b[72])^(a[3] & b[73])^(a[2] & b[74])^(a[1] & b[75])^(a[0] & b[76]);
assign y[77] = (a[77] & b[0])^(a[76] & b[1])^(a[75] & b[2])^(a[74] & b[3])^(a[73] & b[4])^(a[72] & b[5])^(a[71] & b[6])^(a[70] & b[7])^(a[69] & b[8])^(a[68] & b[9])^(a[67] & b[10])^(a[66] & b[11])^(a[65] & b[12])^(a[64] & b[13])^(a[63] & b[14])^(a[62] & b[15])^(a[61] & b[16])^(a[60] & b[17])^(a[59] & b[18])^(a[58] & b[19])^(a[57] & b[20])^(a[56] & b[21])^(a[55] & b[22])^(a[54] & b[23])^(a[53] & b[24])^(a[52] & b[25])^(a[51] & b[26])^(a[50] & b[27])^(a[49] & b[28])^(a[48] & b[29])^(a[47] & b[30])^(a[46] & b[31])^(a[45] & b[32])^(a[44] & b[33])^(a[43] & b[34])^(a[42] & b[35])^(a[41] & b[36])^(a[40] & b[37])^(a[39] & b[38])^(a[38] & b[39])^(a[37] & b[40])^(a[36] & b[41])^(a[35] & b[42])^(a[34] & b[43])^(a[33] & b[44])^(a[32] & b[45])^(a[31] & b[46])^(a[30] & b[47])^(a[29] & b[48])^(a[28] & b[49])^(a[27] & b[50])^(a[26] & b[51])^(a[25] & b[52])^(a[24] & b[53])^(a[23] & b[54])^(a[22] & b[55])^(a[21] & b[56])^(a[20] & b[57])^(a[19] & b[58])^(a[18] & b[59])^(a[17] & b[60])^(a[16] & b[61])^(a[15] & b[62])^(a[14] & b[63])^(a[13] & b[64])^(a[12] & b[65])^(a[11] & b[66])^(a[10] & b[67])^(a[9] & b[68])^(a[8] & b[69])^(a[7] & b[70])^(a[6] & b[71])^(a[5] & b[72])^(a[4] & b[73])^(a[3] & b[74])^(a[2] & b[75])^(a[1] & b[76])^(a[0] & b[77]);
assign y[78] = (a[78] & b[0])^(a[77] & b[1])^(a[76] & b[2])^(a[75] & b[3])^(a[74] & b[4])^(a[73] & b[5])^(a[72] & b[6])^(a[71] & b[7])^(a[70] & b[8])^(a[69] & b[9])^(a[68] & b[10])^(a[67] & b[11])^(a[66] & b[12])^(a[65] & b[13])^(a[64] & b[14])^(a[63] & b[15])^(a[62] & b[16])^(a[61] & b[17])^(a[60] & b[18])^(a[59] & b[19])^(a[58] & b[20])^(a[57] & b[21])^(a[56] & b[22])^(a[55] & b[23])^(a[54] & b[24])^(a[53] & b[25])^(a[52] & b[26])^(a[51] & b[27])^(a[50] & b[28])^(a[49] & b[29])^(a[48] & b[30])^(a[47] & b[31])^(a[46] & b[32])^(a[45] & b[33])^(a[44] & b[34])^(a[43] & b[35])^(a[42] & b[36])^(a[41] & b[37])^(a[40] & b[38])^(a[39] & b[39])^(a[38] & b[40])^(a[37] & b[41])^(a[36] & b[42])^(a[35] & b[43])^(a[34] & b[44])^(a[33] & b[45])^(a[32] & b[46])^(a[31] & b[47])^(a[30] & b[48])^(a[29] & b[49])^(a[28] & b[50])^(a[27] & b[51])^(a[26] & b[52])^(a[25] & b[53])^(a[24] & b[54])^(a[23] & b[55])^(a[22] & b[56])^(a[21] & b[57])^(a[20] & b[58])^(a[19] & b[59])^(a[18] & b[60])^(a[17] & b[61])^(a[16] & b[62])^(a[15] & b[63])^(a[14] & b[64])^(a[13] & b[65])^(a[12] & b[66])^(a[11] & b[67])^(a[10] & b[68])^(a[9] & b[69])^(a[8] & b[70])^(a[7] & b[71])^(a[6] & b[72])^(a[5] & b[73])^(a[4] & b[74])^(a[3] & b[75])^(a[2] & b[76])^(a[1] & b[77])^(a[0] & b[78]);
assign y[79] = (a[79] & b[0])^(a[78] & b[1])^(a[77] & b[2])^(a[76] & b[3])^(a[75] & b[4])^(a[74] & b[5])^(a[73] & b[6])^(a[72] & b[7])^(a[71] & b[8])^(a[70] & b[9])^(a[69] & b[10])^(a[68] & b[11])^(a[67] & b[12])^(a[66] & b[13])^(a[65] & b[14])^(a[64] & b[15])^(a[63] & b[16])^(a[62] & b[17])^(a[61] & b[18])^(a[60] & b[19])^(a[59] & b[20])^(a[58] & b[21])^(a[57] & b[22])^(a[56] & b[23])^(a[55] & b[24])^(a[54] & b[25])^(a[53] & b[26])^(a[52] & b[27])^(a[51] & b[28])^(a[50] & b[29])^(a[49] & b[30])^(a[48] & b[31])^(a[47] & b[32])^(a[46] & b[33])^(a[45] & b[34])^(a[44] & b[35])^(a[43] & b[36])^(a[42] & b[37])^(a[41] & b[38])^(a[40] & b[39])^(a[39] & b[40])^(a[38] & b[41])^(a[37] & b[42])^(a[36] & b[43])^(a[35] & b[44])^(a[34] & b[45])^(a[33] & b[46])^(a[32] & b[47])^(a[31] & b[48])^(a[30] & b[49])^(a[29] & b[50])^(a[28] & b[51])^(a[27] & b[52])^(a[26] & b[53])^(a[25] & b[54])^(a[24] & b[55])^(a[23] & b[56])^(a[22] & b[57])^(a[21] & b[58])^(a[20] & b[59])^(a[19] & b[60])^(a[18] & b[61])^(a[17] & b[62])^(a[16] & b[63])^(a[15] & b[64])^(a[14] & b[65])^(a[13] & b[66])^(a[12] & b[67])^(a[11] & b[68])^(a[10] & b[69])^(a[9] & b[70])^(a[8] & b[71])^(a[7] & b[72])^(a[6] & b[73])^(a[5] & b[74])^(a[4] & b[75])^(a[3] & b[76])^(a[2] & b[77])^(a[1] & b[78])^(a[0] & b[79]);
assign y[80] = (a[80] & b[0])^(a[79] & b[1])^(a[78] & b[2])^(a[77] & b[3])^(a[76] & b[4])^(a[75] & b[5])^(a[74] & b[6])^(a[73] & b[7])^(a[72] & b[8])^(a[71] & b[9])^(a[70] & b[10])^(a[69] & b[11])^(a[68] & b[12])^(a[67] & b[13])^(a[66] & b[14])^(a[65] & b[15])^(a[64] & b[16])^(a[63] & b[17])^(a[62] & b[18])^(a[61] & b[19])^(a[60] & b[20])^(a[59] & b[21])^(a[58] & b[22])^(a[57] & b[23])^(a[56] & b[24])^(a[55] & b[25])^(a[54] & b[26])^(a[53] & b[27])^(a[52] & b[28])^(a[51] & b[29])^(a[50] & b[30])^(a[49] & b[31])^(a[48] & b[32])^(a[47] & b[33])^(a[46] & b[34])^(a[45] & b[35])^(a[44] & b[36])^(a[43] & b[37])^(a[42] & b[38])^(a[41] & b[39])^(a[40] & b[40])^(a[39] & b[41])^(a[38] & b[42])^(a[37] & b[43])^(a[36] & b[44])^(a[35] & b[45])^(a[34] & b[46])^(a[33] & b[47])^(a[32] & b[48])^(a[31] & b[49])^(a[30] & b[50])^(a[29] & b[51])^(a[28] & b[52])^(a[27] & b[53])^(a[26] & b[54])^(a[25] & b[55])^(a[24] & b[56])^(a[23] & b[57])^(a[22] & b[58])^(a[21] & b[59])^(a[20] & b[60])^(a[19] & b[61])^(a[18] & b[62])^(a[17] & b[63])^(a[16] & b[64])^(a[15] & b[65])^(a[14] & b[66])^(a[13] & b[67])^(a[12] & b[68])^(a[11] & b[69])^(a[10] & b[70])^(a[9] & b[71])^(a[8] & b[72])^(a[7] & b[73])^(a[6] & b[74])^(a[5] & b[75])^(a[4] & b[76])^(a[3] & b[77])^(a[2] & b[78])^(a[1] & b[79])^(a[0] & b[80]);
assign y[81] = (a[81] & b[0])^(a[80] & b[1])^(a[79] & b[2])^(a[78] & b[3])^(a[77] & b[4])^(a[76] & b[5])^(a[75] & b[6])^(a[74] & b[7])^(a[73] & b[8])^(a[72] & b[9])^(a[71] & b[10])^(a[70] & b[11])^(a[69] & b[12])^(a[68] & b[13])^(a[67] & b[14])^(a[66] & b[15])^(a[65] & b[16])^(a[64] & b[17])^(a[63] & b[18])^(a[62] & b[19])^(a[61] & b[20])^(a[60] & b[21])^(a[59] & b[22])^(a[58] & b[23])^(a[57] & b[24])^(a[56] & b[25])^(a[55] & b[26])^(a[54] & b[27])^(a[53] & b[28])^(a[52] & b[29])^(a[51] & b[30])^(a[50] & b[31])^(a[49] & b[32])^(a[48] & b[33])^(a[47] & b[34])^(a[46] & b[35])^(a[45] & b[36])^(a[44] & b[37])^(a[43] & b[38])^(a[42] & b[39])^(a[41] & b[40])^(a[40] & b[41])^(a[39] & b[42])^(a[38] & b[43])^(a[37] & b[44])^(a[36] & b[45])^(a[35] & b[46])^(a[34] & b[47])^(a[33] & b[48])^(a[32] & b[49])^(a[31] & b[50])^(a[30] & b[51])^(a[29] & b[52])^(a[28] & b[53])^(a[27] & b[54])^(a[26] & b[55])^(a[25] & b[56])^(a[24] & b[57])^(a[23] & b[58])^(a[22] & b[59])^(a[21] & b[60])^(a[20] & b[61])^(a[19] & b[62])^(a[18] & b[63])^(a[17] & b[64])^(a[16] & b[65])^(a[15] & b[66])^(a[14] & b[67])^(a[13] & b[68])^(a[12] & b[69])^(a[11] & b[70])^(a[10] & b[71])^(a[9] & b[72])^(a[8] & b[73])^(a[7] & b[74])^(a[6] & b[75])^(a[5] & b[76])^(a[4] & b[77])^(a[3] & b[78])^(a[2] & b[79])^(a[1] & b[80])^(a[0] & b[81]);
assign y[82] = (a[82] & b[0])^(a[81] & b[1])^(a[80] & b[2])^(a[79] & b[3])^(a[78] & b[4])^(a[77] & b[5])^(a[76] & b[6])^(a[75] & b[7])^(a[74] & b[8])^(a[73] & b[9])^(a[72] & b[10])^(a[71] & b[11])^(a[70] & b[12])^(a[69] & b[13])^(a[68] & b[14])^(a[67] & b[15])^(a[66] & b[16])^(a[65] & b[17])^(a[64] & b[18])^(a[63] & b[19])^(a[62] & b[20])^(a[61] & b[21])^(a[60] & b[22])^(a[59] & b[23])^(a[58] & b[24])^(a[57] & b[25])^(a[56] & b[26])^(a[55] & b[27])^(a[54] & b[28])^(a[53] & b[29])^(a[52] & b[30])^(a[51] & b[31])^(a[50] & b[32])^(a[49] & b[33])^(a[48] & b[34])^(a[47] & b[35])^(a[46] & b[36])^(a[45] & b[37])^(a[44] & b[38])^(a[43] & b[39])^(a[42] & b[40])^(a[41] & b[41])^(a[40] & b[42])^(a[39] & b[43])^(a[38] & b[44])^(a[37] & b[45])^(a[36] & b[46])^(a[35] & b[47])^(a[34] & b[48])^(a[33] & b[49])^(a[32] & b[50])^(a[31] & b[51])^(a[30] & b[52])^(a[29] & b[53])^(a[28] & b[54])^(a[27] & b[55])^(a[26] & b[56])^(a[25] & b[57])^(a[24] & b[58])^(a[23] & b[59])^(a[22] & b[60])^(a[21] & b[61])^(a[20] & b[62])^(a[19] & b[63])^(a[18] & b[64])^(a[17] & b[65])^(a[16] & b[66])^(a[15] & b[67])^(a[14] & b[68])^(a[13] & b[69])^(a[12] & b[70])^(a[11] & b[71])^(a[10] & b[72])^(a[9] & b[73])^(a[8] & b[74])^(a[7] & b[75])^(a[6] & b[76])^(a[5] & b[77])^(a[4] & b[78])^(a[3] & b[79])^(a[2] & b[80])^(a[1] & b[81])^(a[0] & b[82]);
assign y[83] = (a[83] & b[0])^(a[82] & b[1])^(a[81] & b[2])^(a[80] & b[3])^(a[79] & b[4])^(a[78] & b[5])^(a[77] & b[6])^(a[76] & b[7])^(a[75] & b[8])^(a[74] & b[9])^(a[73] & b[10])^(a[72] & b[11])^(a[71] & b[12])^(a[70] & b[13])^(a[69] & b[14])^(a[68] & b[15])^(a[67] & b[16])^(a[66] & b[17])^(a[65] & b[18])^(a[64] & b[19])^(a[63] & b[20])^(a[62] & b[21])^(a[61] & b[22])^(a[60] & b[23])^(a[59] & b[24])^(a[58] & b[25])^(a[57] & b[26])^(a[56] & b[27])^(a[55] & b[28])^(a[54] & b[29])^(a[53] & b[30])^(a[52] & b[31])^(a[51] & b[32])^(a[50] & b[33])^(a[49] & b[34])^(a[48] & b[35])^(a[47] & b[36])^(a[46] & b[37])^(a[45] & b[38])^(a[44] & b[39])^(a[43] & b[40])^(a[42] & b[41])^(a[41] & b[42])^(a[40] & b[43])^(a[39] & b[44])^(a[38] & b[45])^(a[37] & b[46])^(a[36] & b[47])^(a[35] & b[48])^(a[34] & b[49])^(a[33] & b[50])^(a[32] & b[51])^(a[31] & b[52])^(a[30] & b[53])^(a[29] & b[54])^(a[28] & b[55])^(a[27] & b[56])^(a[26] & b[57])^(a[25] & b[58])^(a[24] & b[59])^(a[23] & b[60])^(a[22] & b[61])^(a[21] & b[62])^(a[20] & b[63])^(a[19] & b[64])^(a[18] & b[65])^(a[17] & b[66])^(a[16] & b[67])^(a[15] & b[68])^(a[14] & b[69])^(a[13] & b[70])^(a[12] & b[71])^(a[11] & b[72])^(a[10] & b[73])^(a[9] & b[74])^(a[8] & b[75])^(a[7] & b[76])^(a[6] & b[77])^(a[5] & b[78])^(a[4] & b[79])^(a[3] & b[80])^(a[2] & b[81])^(a[1] & b[82])^(a[0] & b[83]);
assign y[84] = (a[84] & b[0])^(a[83] & b[1])^(a[82] & b[2])^(a[81] & b[3])^(a[80] & b[4])^(a[79] & b[5])^(a[78] & b[6])^(a[77] & b[7])^(a[76] & b[8])^(a[75] & b[9])^(a[74] & b[10])^(a[73] & b[11])^(a[72] & b[12])^(a[71] & b[13])^(a[70] & b[14])^(a[69] & b[15])^(a[68] & b[16])^(a[67] & b[17])^(a[66] & b[18])^(a[65] & b[19])^(a[64] & b[20])^(a[63] & b[21])^(a[62] & b[22])^(a[61] & b[23])^(a[60] & b[24])^(a[59] & b[25])^(a[58] & b[26])^(a[57] & b[27])^(a[56] & b[28])^(a[55] & b[29])^(a[54] & b[30])^(a[53] & b[31])^(a[52] & b[32])^(a[51] & b[33])^(a[50] & b[34])^(a[49] & b[35])^(a[48] & b[36])^(a[47] & b[37])^(a[46] & b[38])^(a[45] & b[39])^(a[44] & b[40])^(a[43] & b[41])^(a[42] & b[42])^(a[41] & b[43])^(a[40] & b[44])^(a[39] & b[45])^(a[38] & b[46])^(a[37] & b[47])^(a[36] & b[48])^(a[35] & b[49])^(a[34] & b[50])^(a[33] & b[51])^(a[32] & b[52])^(a[31] & b[53])^(a[30] & b[54])^(a[29] & b[55])^(a[28] & b[56])^(a[27] & b[57])^(a[26] & b[58])^(a[25] & b[59])^(a[24] & b[60])^(a[23] & b[61])^(a[22] & b[62])^(a[21] & b[63])^(a[20] & b[64])^(a[19] & b[65])^(a[18] & b[66])^(a[17] & b[67])^(a[16] & b[68])^(a[15] & b[69])^(a[14] & b[70])^(a[13] & b[71])^(a[12] & b[72])^(a[11] & b[73])^(a[10] & b[74])^(a[9] & b[75])^(a[8] & b[76])^(a[7] & b[77])^(a[6] & b[78])^(a[5] & b[79])^(a[4] & b[80])^(a[3] & b[81])^(a[2] & b[82])^(a[1] & b[83])^(a[0] & b[84]);
assign y[85] = (a[85] & b[0])^(a[84] & b[1])^(a[83] & b[2])^(a[82] & b[3])^(a[81] & b[4])^(a[80] & b[5])^(a[79] & b[6])^(a[78] & b[7])^(a[77] & b[8])^(a[76] & b[9])^(a[75] & b[10])^(a[74] & b[11])^(a[73] & b[12])^(a[72] & b[13])^(a[71] & b[14])^(a[70] & b[15])^(a[69] & b[16])^(a[68] & b[17])^(a[67] & b[18])^(a[66] & b[19])^(a[65] & b[20])^(a[64] & b[21])^(a[63] & b[22])^(a[62] & b[23])^(a[61] & b[24])^(a[60] & b[25])^(a[59] & b[26])^(a[58] & b[27])^(a[57] & b[28])^(a[56] & b[29])^(a[55] & b[30])^(a[54] & b[31])^(a[53] & b[32])^(a[52] & b[33])^(a[51] & b[34])^(a[50] & b[35])^(a[49] & b[36])^(a[48] & b[37])^(a[47] & b[38])^(a[46] & b[39])^(a[45] & b[40])^(a[44] & b[41])^(a[43] & b[42])^(a[42] & b[43])^(a[41] & b[44])^(a[40] & b[45])^(a[39] & b[46])^(a[38] & b[47])^(a[37] & b[48])^(a[36] & b[49])^(a[35] & b[50])^(a[34] & b[51])^(a[33] & b[52])^(a[32] & b[53])^(a[31] & b[54])^(a[30] & b[55])^(a[29] & b[56])^(a[28] & b[57])^(a[27] & b[58])^(a[26] & b[59])^(a[25] & b[60])^(a[24] & b[61])^(a[23] & b[62])^(a[22] & b[63])^(a[21] & b[64])^(a[20] & b[65])^(a[19] & b[66])^(a[18] & b[67])^(a[17] & b[68])^(a[16] & b[69])^(a[15] & b[70])^(a[14] & b[71])^(a[13] & b[72])^(a[12] & b[73])^(a[11] & b[74])^(a[10] & b[75])^(a[9] & b[76])^(a[8] & b[77])^(a[7] & b[78])^(a[6] & b[79])^(a[5] & b[80])^(a[4] & b[81])^(a[3] & b[82])^(a[2] & b[83])^(a[1] & b[84])^(a[0] & b[85]);
assign y[86] = (a[86] & b[0])^(a[85] & b[1])^(a[84] & b[2])^(a[83] & b[3])^(a[82] & b[4])^(a[81] & b[5])^(a[80] & b[6])^(a[79] & b[7])^(a[78] & b[8])^(a[77] & b[9])^(a[76] & b[10])^(a[75] & b[11])^(a[74] & b[12])^(a[73] & b[13])^(a[72] & b[14])^(a[71] & b[15])^(a[70] & b[16])^(a[69] & b[17])^(a[68] & b[18])^(a[67] & b[19])^(a[66] & b[20])^(a[65] & b[21])^(a[64] & b[22])^(a[63] & b[23])^(a[62] & b[24])^(a[61] & b[25])^(a[60] & b[26])^(a[59] & b[27])^(a[58] & b[28])^(a[57] & b[29])^(a[56] & b[30])^(a[55] & b[31])^(a[54] & b[32])^(a[53] & b[33])^(a[52] & b[34])^(a[51] & b[35])^(a[50] & b[36])^(a[49] & b[37])^(a[48] & b[38])^(a[47] & b[39])^(a[46] & b[40])^(a[45] & b[41])^(a[44] & b[42])^(a[43] & b[43])^(a[42] & b[44])^(a[41] & b[45])^(a[40] & b[46])^(a[39] & b[47])^(a[38] & b[48])^(a[37] & b[49])^(a[36] & b[50])^(a[35] & b[51])^(a[34] & b[52])^(a[33] & b[53])^(a[32] & b[54])^(a[31] & b[55])^(a[30] & b[56])^(a[29] & b[57])^(a[28] & b[58])^(a[27] & b[59])^(a[26] & b[60])^(a[25] & b[61])^(a[24] & b[62])^(a[23] & b[63])^(a[22] & b[64])^(a[21] & b[65])^(a[20] & b[66])^(a[19] & b[67])^(a[18] & b[68])^(a[17] & b[69])^(a[16] & b[70])^(a[15] & b[71])^(a[14] & b[72])^(a[13] & b[73])^(a[12] & b[74])^(a[11] & b[75])^(a[10] & b[76])^(a[9] & b[77])^(a[8] & b[78])^(a[7] & b[79])^(a[6] & b[80])^(a[5] & b[81])^(a[4] & b[82])^(a[3] & b[83])^(a[2] & b[84])^(a[1] & b[85])^(a[0] & b[86]);
assign y[87] = (a[87] & b[0])^(a[86] & b[1])^(a[85] & b[2])^(a[84] & b[3])^(a[83] & b[4])^(a[82] & b[5])^(a[81] & b[6])^(a[80] & b[7])^(a[79] & b[8])^(a[78] & b[9])^(a[77] & b[10])^(a[76] & b[11])^(a[75] & b[12])^(a[74] & b[13])^(a[73] & b[14])^(a[72] & b[15])^(a[71] & b[16])^(a[70] & b[17])^(a[69] & b[18])^(a[68] & b[19])^(a[67] & b[20])^(a[66] & b[21])^(a[65] & b[22])^(a[64] & b[23])^(a[63] & b[24])^(a[62] & b[25])^(a[61] & b[26])^(a[60] & b[27])^(a[59] & b[28])^(a[58] & b[29])^(a[57] & b[30])^(a[56] & b[31])^(a[55] & b[32])^(a[54] & b[33])^(a[53] & b[34])^(a[52] & b[35])^(a[51] & b[36])^(a[50] & b[37])^(a[49] & b[38])^(a[48] & b[39])^(a[47] & b[40])^(a[46] & b[41])^(a[45] & b[42])^(a[44] & b[43])^(a[43] & b[44])^(a[42] & b[45])^(a[41] & b[46])^(a[40] & b[47])^(a[39] & b[48])^(a[38] & b[49])^(a[37] & b[50])^(a[36] & b[51])^(a[35] & b[52])^(a[34] & b[53])^(a[33] & b[54])^(a[32] & b[55])^(a[31] & b[56])^(a[30] & b[57])^(a[29] & b[58])^(a[28] & b[59])^(a[27] & b[60])^(a[26] & b[61])^(a[25] & b[62])^(a[24] & b[63])^(a[23] & b[64])^(a[22] & b[65])^(a[21] & b[66])^(a[20] & b[67])^(a[19] & b[68])^(a[18] & b[69])^(a[17] & b[70])^(a[16] & b[71])^(a[15] & b[72])^(a[14] & b[73])^(a[13] & b[74])^(a[12] & b[75])^(a[11] & b[76])^(a[10] & b[77])^(a[9] & b[78])^(a[8] & b[79])^(a[7] & b[80])^(a[6] & b[81])^(a[5] & b[82])^(a[4] & b[83])^(a[3] & b[84])^(a[2] & b[85])^(a[1] & b[86])^(a[0] & b[87]);
assign y[88] = (a[88] & b[0])^(a[87] & b[1])^(a[86] & b[2])^(a[85] & b[3])^(a[84] & b[4])^(a[83] & b[5])^(a[82] & b[6])^(a[81] & b[7])^(a[80] & b[8])^(a[79] & b[9])^(a[78] & b[10])^(a[77] & b[11])^(a[76] & b[12])^(a[75] & b[13])^(a[74] & b[14])^(a[73] & b[15])^(a[72] & b[16])^(a[71] & b[17])^(a[70] & b[18])^(a[69] & b[19])^(a[68] & b[20])^(a[67] & b[21])^(a[66] & b[22])^(a[65] & b[23])^(a[64] & b[24])^(a[63] & b[25])^(a[62] & b[26])^(a[61] & b[27])^(a[60] & b[28])^(a[59] & b[29])^(a[58] & b[30])^(a[57] & b[31])^(a[56] & b[32])^(a[55] & b[33])^(a[54] & b[34])^(a[53] & b[35])^(a[52] & b[36])^(a[51] & b[37])^(a[50] & b[38])^(a[49] & b[39])^(a[48] & b[40])^(a[47] & b[41])^(a[46] & b[42])^(a[45] & b[43])^(a[44] & b[44])^(a[43] & b[45])^(a[42] & b[46])^(a[41] & b[47])^(a[40] & b[48])^(a[39] & b[49])^(a[38] & b[50])^(a[37] & b[51])^(a[36] & b[52])^(a[35] & b[53])^(a[34] & b[54])^(a[33] & b[55])^(a[32] & b[56])^(a[31] & b[57])^(a[30] & b[58])^(a[29] & b[59])^(a[28] & b[60])^(a[27] & b[61])^(a[26] & b[62])^(a[25] & b[63])^(a[24] & b[64])^(a[23] & b[65])^(a[22] & b[66])^(a[21] & b[67])^(a[20] & b[68])^(a[19] & b[69])^(a[18] & b[70])^(a[17] & b[71])^(a[16] & b[72])^(a[15] & b[73])^(a[14] & b[74])^(a[13] & b[75])^(a[12] & b[76])^(a[11] & b[77])^(a[10] & b[78])^(a[9] & b[79])^(a[8] & b[80])^(a[7] & b[81])^(a[6] & b[82])^(a[5] & b[83])^(a[4] & b[84])^(a[3] & b[85])^(a[2] & b[86])^(a[1] & b[87])^(a[0] & b[88]);
assign y[89] = (a[89] & b[0])^(a[88] & b[1])^(a[87] & b[2])^(a[86] & b[3])^(a[85] & b[4])^(a[84] & b[5])^(a[83] & b[6])^(a[82] & b[7])^(a[81] & b[8])^(a[80] & b[9])^(a[79] & b[10])^(a[78] & b[11])^(a[77] & b[12])^(a[76] & b[13])^(a[75] & b[14])^(a[74] & b[15])^(a[73] & b[16])^(a[72] & b[17])^(a[71] & b[18])^(a[70] & b[19])^(a[69] & b[20])^(a[68] & b[21])^(a[67] & b[22])^(a[66] & b[23])^(a[65] & b[24])^(a[64] & b[25])^(a[63] & b[26])^(a[62] & b[27])^(a[61] & b[28])^(a[60] & b[29])^(a[59] & b[30])^(a[58] & b[31])^(a[57] & b[32])^(a[56] & b[33])^(a[55] & b[34])^(a[54] & b[35])^(a[53] & b[36])^(a[52] & b[37])^(a[51] & b[38])^(a[50] & b[39])^(a[49] & b[40])^(a[48] & b[41])^(a[47] & b[42])^(a[46] & b[43])^(a[45] & b[44])^(a[44] & b[45])^(a[43] & b[46])^(a[42] & b[47])^(a[41] & b[48])^(a[40] & b[49])^(a[39] & b[50])^(a[38] & b[51])^(a[37] & b[52])^(a[36] & b[53])^(a[35] & b[54])^(a[34] & b[55])^(a[33] & b[56])^(a[32] & b[57])^(a[31] & b[58])^(a[30] & b[59])^(a[29] & b[60])^(a[28] & b[61])^(a[27] & b[62])^(a[26] & b[63])^(a[25] & b[64])^(a[24] & b[65])^(a[23] & b[66])^(a[22] & b[67])^(a[21] & b[68])^(a[20] & b[69])^(a[19] & b[70])^(a[18] & b[71])^(a[17] & b[72])^(a[16] & b[73])^(a[15] & b[74])^(a[14] & b[75])^(a[13] & b[76])^(a[12] & b[77])^(a[11] & b[78])^(a[10] & b[79])^(a[9] & b[80])^(a[8] & b[81])^(a[7] & b[82])^(a[6] & b[83])^(a[5] & b[84])^(a[4] & b[85])^(a[3] & b[86])^(a[2] & b[87])^(a[1] & b[88])^(a[0] & b[89]);
assign y[90] = (a[90] & b[0])^(a[89] & b[1])^(a[88] & b[2])^(a[87] & b[3])^(a[86] & b[4])^(a[85] & b[5])^(a[84] & b[6])^(a[83] & b[7])^(a[82] & b[8])^(a[81] & b[9])^(a[80] & b[10])^(a[79] & b[11])^(a[78] & b[12])^(a[77] & b[13])^(a[76] & b[14])^(a[75] & b[15])^(a[74] & b[16])^(a[73] & b[17])^(a[72] & b[18])^(a[71] & b[19])^(a[70] & b[20])^(a[69] & b[21])^(a[68] & b[22])^(a[67] & b[23])^(a[66] & b[24])^(a[65] & b[25])^(a[64] & b[26])^(a[63] & b[27])^(a[62] & b[28])^(a[61] & b[29])^(a[60] & b[30])^(a[59] & b[31])^(a[58] & b[32])^(a[57] & b[33])^(a[56] & b[34])^(a[55] & b[35])^(a[54] & b[36])^(a[53] & b[37])^(a[52] & b[38])^(a[51] & b[39])^(a[50] & b[40])^(a[49] & b[41])^(a[48] & b[42])^(a[47] & b[43])^(a[46] & b[44])^(a[45] & b[45])^(a[44] & b[46])^(a[43] & b[47])^(a[42] & b[48])^(a[41] & b[49])^(a[40] & b[50])^(a[39] & b[51])^(a[38] & b[52])^(a[37] & b[53])^(a[36] & b[54])^(a[35] & b[55])^(a[34] & b[56])^(a[33] & b[57])^(a[32] & b[58])^(a[31] & b[59])^(a[30] & b[60])^(a[29] & b[61])^(a[28] & b[62])^(a[27] & b[63])^(a[26] & b[64])^(a[25] & b[65])^(a[24] & b[66])^(a[23] & b[67])^(a[22] & b[68])^(a[21] & b[69])^(a[20] & b[70])^(a[19] & b[71])^(a[18] & b[72])^(a[17] & b[73])^(a[16] & b[74])^(a[15] & b[75])^(a[14] & b[76])^(a[13] & b[77])^(a[12] & b[78])^(a[11] & b[79])^(a[10] & b[80])^(a[9] & b[81])^(a[8] & b[82])^(a[7] & b[83])^(a[6] & b[84])^(a[5] & b[85])^(a[4] & b[86])^(a[3] & b[87])^(a[2] & b[88])^(a[1] & b[89])^(a[0] & b[90]);
assign y[91] = (a[91] & b[0])^(a[90] & b[1])^(a[89] & b[2])^(a[88] & b[3])^(a[87] & b[4])^(a[86] & b[5])^(a[85] & b[6])^(a[84] & b[7])^(a[83] & b[8])^(a[82] & b[9])^(a[81] & b[10])^(a[80] & b[11])^(a[79] & b[12])^(a[78] & b[13])^(a[77] & b[14])^(a[76] & b[15])^(a[75] & b[16])^(a[74] & b[17])^(a[73] & b[18])^(a[72] & b[19])^(a[71] & b[20])^(a[70] & b[21])^(a[69] & b[22])^(a[68] & b[23])^(a[67] & b[24])^(a[66] & b[25])^(a[65] & b[26])^(a[64] & b[27])^(a[63] & b[28])^(a[62] & b[29])^(a[61] & b[30])^(a[60] & b[31])^(a[59] & b[32])^(a[58] & b[33])^(a[57] & b[34])^(a[56] & b[35])^(a[55] & b[36])^(a[54] & b[37])^(a[53] & b[38])^(a[52] & b[39])^(a[51] & b[40])^(a[50] & b[41])^(a[49] & b[42])^(a[48] & b[43])^(a[47] & b[44])^(a[46] & b[45])^(a[45] & b[46])^(a[44] & b[47])^(a[43] & b[48])^(a[42] & b[49])^(a[41] & b[50])^(a[40] & b[51])^(a[39] & b[52])^(a[38] & b[53])^(a[37] & b[54])^(a[36] & b[55])^(a[35] & b[56])^(a[34] & b[57])^(a[33] & b[58])^(a[32] & b[59])^(a[31] & b[60])^(a[30] & b[61])^(a[29] & b[62])^(a[28] & b[63])^(a[27] & b[64])^(a[26] & b[65])^(a[25] & b[66])^(a[24] & b[67])^(a[23] & b[68])^(a[22] & b[69])^(a[21] & b[70])^(a[20] & b[71])^(a[19] & b[72])^(a[18] & b[73])^(a[17] & b[74])^(a[16] & b[75])^(a[15] & b[76])^(a[14] & b[77])^(a[13] & b[78])^(a[12] & b[79])^(a[11] & b[80])^(a[10] & b[81])^(a[9] & b[82])^(a[8] & b[83])^(a[7] & b[84])^(a[6] & b[85])^(a[5] & b[86])^(a[4] & b[87])^(a[3] & b[88])^(a[2] & b[89])^(a[1] & b[90])^(a[0] & b[91]);
assign y[92] = (a[92] & b[0])^(a[91] & b[1])^(a[90] & b[2])^(a[89] & b[3])^(a[88] & b[4])^(a[87] & b[5])^(a[86] & b[6])^(a[85] & b[7])^(a[84] & b[8])^(a[83] & b[9])^(a[82] & b[10])^(a[81] & b[11])^(a[80] & b[12])^(a[79] & b[13])^(a[78] & b[14])^(a[77] & b[15])^(a[76] & b[16])^(a[75] & b[17])^(a[74] & b[18])^(a[73] & b[19])^(a[72] & b[20])^(a[71] & b[21])^(a[70] & b[22])^(a[69] & b[23])^(a[68] & b[24])^(a[67] & b[25])^(a[66] & b[26])^(a[65] & b[27])^(a[64] & b[28])^(a[63] & b[29])^(a[62] & b[30])^(a[61] & b[31])^(a[60] & b[32])^(a[59] & b[33])^(a[58] & b[34])^(a[57] & b[35])^(a[56] & b[36])^(a[55] & b[37])^(a[54] & b[38])^(a[53] & b[39])^(a[52] & b[40])^(a[51] & b[41])^(a[50] & b[42])^(a[49] & b[43])^(a[48] & b[44])^(a[47] & b[45])^(a[46] & b[46])^(a[45] & b[47])^(a[44] & b[48])^(a[43] & b[49])^(a[42] & b[50])^(a[41] & b[51])^(a[40] & b[52])^(a[39] & b[53])^(a[38] & b[54])^(a[37] & b[55])^(a[36] & b[56])^(a[35] & b[57])^(a[34] & b[58])^(a[33] & b[59])^(a[32] & b[60])^(a[31] & b[61])^(a[30] & b[62])^(a[29] & b[63])^(a[28] & b[64])^(a[27] & b[65])^(a[26] & b[66])^(a[25] & b[67])^(a[24] & b[68])^(a[23] & b[69])^(a[22] & b[70])^(a[21] & b[71])^(a[20] & b[72])^(a[19] & b[73])^(a[18] & b[74])^(a[17] & b[75])^(a[16] & b[76])^(a[15] & b[77])^(a[14] & b[78])^(a[13] & b[79])^(a[12] & b[80])^(a[11] & b[81])^(a[10] & b[82])^(a[9] & b[83])^(a[8] & b[84])^(a[7] & b[85])^(a[6] & b[86])^(a[5] & b[87])^(a[4] & b[88])^(a[3] & b[89])^(a[2] & b[90])^(a[1] & b[91])^(a[0] & b[92]);
assign y[93] = (a[93] & b[0])^(a[92] & b[1])^(a[91] & b[2])^(a[90] & b[3])^(a[89] & b[4])^(a[88] & b[5])^(a[87] & b[6])^(a[86] & b[7])^(a[85] & b[8])^(a[84] & b[9])^(a[83] & b[10])^(a[82] & b[11])^(a[81] & b[12])^(a[80] & b[13])^(a[79] & b[14])^(a[78] & b[15])^(a[77] & b[16])^(a[76] & b[17])^(a[75] & b[18])^(a[74] & b[19])^(a[73] & b[20])^(a[72] & b[21])^(a[71] & b[22])^(a[70] & b[23])^(a[69] & b[24])^(a[68] & b[25])^(a[67] & b[26])^(a[66] & b[27])^(a[65] & b[28])^(a[64] & b[29])^(a[63] & b[30])^(a[62] & b[31])^(a[61] & b[32])^(a[60] & b[33])^(a[59] & b[34])^(a[58] & b[35])^(a[57] & b[36])^(a[56] & b[37])^(a[55] & b[38])^(a[54] & b[39])^(a[53] & b[40])^(a[52] & b[41])^(a[51] & b[42])^(a[50] & b[43])^(a[49] & b[44])^(a[48] & b[45])^(a[47] & b[46])^(a[46] & b[47])^(a[45] & b[48])^(a[44] & b[49])^(a[43] & b[50])^(a[42] & b[51])^(a[41] & b[52])^(a[40] & b[53])^(a[39] & b[54])^(a[38] & b[55])^(a[37] & b[56])^(a[36] & b[57])^(a[35] & b[58])^(a[34] & b[59])^(a[33] & b[60])^(a[32] & b[61])^(a[31] & b[62])^(a[30] & b[63])^(a[29] & b[64])^(a[28] & b[65])^(a[27] & b[66])^(a[26] & b[67])^(a[25] & b[68])^(a[24] & b[69])^(a[23] & b[70])^(a[22] & b[71])^(a[21] & b[72])^(a[20] & b[73])^(a[19] & b[74])^(a[18] & b[75])^(a[17] & b[76])^(a[16] & b[77])^(a[15] & b[78])^(a[14] & b[79])^(a[13] & b[80])^(a[12] & b[81])^(a[11] & b[82])^(a[10] & b[83])^(a[9] & b[84])^(a[8] & b[85])^(a[7] & b[86])^(a[6] & b[87])^(a[5] & b[88])^(a[4] & b[89])^(a[3] & b[90])^(a[2] & b[91])^(a[1] & b[92])^(a[0] & b[93]);
assign y[94] = (a[94] & b[0])^(a[93] & b[1])^(a[92] & b[2])^(a[91] & b[3])^(a[90] & b[4])^(a[89] & b[5])^(a[88] & b[6])^(a[87] & b[7])^(a[86] & b[8])^(a[85] & b[9])^(a[84] & b[10])^(a[83] & b[11])^(a[82] & b[12])^(a[81] & b[13])^(a[80] & b[14])^(a[79] & b[15])^(a[78] & b[16])^(a[77] & b[17])^(a[76] & b[18])^(a[75] & b[19])^(a[74] & b[20])^(a[73] & b[21])^(a[72] & b[22])^(a[71] & b[23])^(a[70] & b[24])^(a[69] & b[25])^(a[68] & b[26])^(a[67] & b[27])^(a[66] & b[28])^(a[65] & b[29])^(a[64] & b[30])^(a[63] & b[31])^(a[62] & b[32])^(a[61] & b[33])^(a[60] & b[34])^(a[59] & b[35])^(a[58] & b[36])^(a[57] & b[37])^(a[56] & b[38])^(a[55] & b[39])^(a[54] & b[40])^(a[53] & b[41])^(a[52] & b[42])^(a[51] & b[43])^(a[50] & b[44])^(a[49] & b[45])^(a[48] & b[46])^(a[47] & b[47])^(a[46] & b[48])^(a[45] & b[49])^(a[44] & b[50])^(a[43] & b[51])^(a[42] & b[52])^(a[41] & b[53])^(a[40] & b[54])^(a[39] & b[55])^(a[38] & b[56])^(a[37] & b[57])^(a[36] & b[58])^(a[35] & b[59])^(a[34] & b[60])^(a[33] & b[61])^(a[32] & b[62])^(a[31] & b[63])^(a[30] & b[64])^(a[29] & b[65])^(a[28] & b[66])^(a[27] & b[67])^(a[26] & b[68])^(a[25] & b[69])^(a[24] & b[70])^(a[23] & b[71])^(a[22] & b[72])^(a[21] & b[73])^(a[20] & b[74])^(a[19] & b[75])^(a[18] & b[76])^(a[17] & b[77])^(a[16] & b[78])^(a[15] & b[79])^(a[14] & b[80])^(a[13] & b[81])^(a[12] & b[82])^(a[11] & b[83])^(a[10] & b[84])^(a[9] & b[85])^(a[8] & b[86])^(a[7] & b[87])^(a[6] & b[88])^(a[5] & b[89])^(a[4] & b[90])^(a[3] & b[91])^(a[2] & b[92])^(a[1] & b[93])^(a[0] & b[94]);
assign y[95] = (a[95] & b[0])^(a[94] & b[1])^(a[93] & b[2])^(a[92] & b[3])^(a[91] & b[4])^(a[90] & b[5])^(a[89] & b[6])^(a[88] & b[7])^(a[87] & b[8])^(a[86] & b[9])^(a[85] & b[10])^(a[84] & b[11])^(a[83] & b[12])^(a[82] & b[13])^(a[81] & b[14])^(a[80] & b[15])^(a[79] & b[16])^(a[78] & b[17])^(a[77] & b[18])^(a[76] & b[19])^(a[75] & b[20])^(a[74] & b[21])^(a[73] & b[22])^(a[72] & b[23])^(a[71] & b[24])^(a[70] & b[25])^(a[69] & b[26])^(a[68] & b[27])^(a[67] & b[28])^(a[66] & b[29])^(a[65] & b[30])^(a[64] & b[31])^(a[63] & b[32])^(a[62] & b[33])^(a[61] & b[34])^(a[60] & b[35])^(a[59] & b[36])^(a[58] & b[37])^(a[57] & b[38])^(a[56] & b[39])^(a[55] & b[40])^(a[54] & b[41])^(a[53] & b[42])^(a[52] & b[43])^(a[51] & b[44])^(a[50] & b[45])^(a[49] & b[46])^(a[48] & b[47])^(a[47] & b[48])^(a[46] & b[49])^(a[45] & b[50])^(a[44] & b[51])^(a[43] & b[52])^(a[42] & b[53])^(a[41] & b[54])^(a[40] & b[55])^(a[39] & b[56])^(a[38] & b[57])^(a[37] & b[58])^(a[36] & b[59])^(a[35] & b[60])^(a[34] & b[61])^(a[33] & b[62])^(a[32] & b[63])^(a[31] & b[64])^(a[30] & b[65])^(a[29] & b[66])^(a[28] & b[67])^(a[27] & b[68])^(a[26] & b[69])^(a[25] & b[70])^(a[24] & b[71])^(a[23] & b[72])^(a[22] & b[73])^(a[21] & b[74])^(a[20] & b[75])^(a[19] & b[76])^(a[18] & b[77])^(a[17] & b[78])^(a[16] & b[79])^(a[15] & b[80])^(a[14] & b[81])^(a[13] & b[82])^(a[12] & b[83])^(a[11] & b[84])^(a[10] & b[85])^(a[9] & b[86])^(a[8] & b[87])^(a[7] & b[88])^(a[6] & b[89])^(a[5] & b[90])^(a[4] & b[91])^(a[3] & b[92])^(a[2] & b[93])^(a[1] & b[94])^(a[0] & b[95]);
assign y[96] = (a[96] & b[0])^(a[95] & b[1])^(a[94] & b[2])^(a[93] & b[3])^(a[92] & b[4])^(a[91] & b[5])^(a[90] & b[6])^(a[89] & b[7])^(a[88] & b[8])^(a[87] & b[9])^(a[86] & b[10])^(a[85] & b[11])^(a[84] & b[12])^(a[83] & b[13])^(a[82] & b[14])^(a[81] & b[15])^(a[80] & b[16])^(a[79] & b[17])^(a[78] & b[18])^(a[77] & b[19])^(a[76] & b[20])^(a[75] & b[21])^(a[74] & b[22])^(a[73] & b[23])^(a[72] & b[24])^(a[71] & b[25])^(a[70] & b[26])^(a[69] & b[27])^(a[68] & b[28])^(a[67] & b[29])^(a[66] & b[30])^(a[65] & b[31])^(a[64] & b[32])^(a[63] & b[33])^(a[62] & b[34])^(a[61] & b[35])^(a[60] & b[36])^(a[59] & b[37])^(a[58] & b[38])^(a[57] & b[39])^(a[56] & b[40])^(a[55] & b[41])^(a[54] & b[42])^(a[53] & b[43])^(a[52] & b[44])^(a[51] & b[45])^(a[50] & b[46])^(a[49] & b[47])^(a[48] & b[48])^(a[47] & b[49])^(a[46] & b[50])^(a[45] & b[51])^(a[44] & b[52])^(a[43] & b[53])^(a[42] & b[54])^(a[41] & b[55])^(a[40] & b[56])^(a[39] & b[57])^(a[38] & b[58])^(a[37] & b[59])^(a[36] & b[60])^(a[35] & b[61])^(a[34] & b[62])^(a[33] & b[63])^(a[32] & b[64])^(a[31] & b[65])^(a[30] & b[66])^(a[29] & b[67])^(a[28] & b[68])^(a[27] & b[69])^(a[26] & b[70])^(a[25] & b[71])^(a[24] & b[72])^(a[23] & b[73])^(a[22] & b[74])^(a[21] & b[75])^(a[20] & b[76])^(a[19] & b[77])^(a[18] & b[78])^(a[17] & b[79])^(a[16] & b[80])^(a[15] & b[81])^(a[14] & b[82])^(a[13] & b[83])^(a[12] & b[84])^(a[11] & b[85])^(a[10] & b[86])^(a[9] & b[87])^(a[8] & b[88])^(a[7] & b[89])^(a[6] & b[90])^(a[5] & b[91])^(a[4] & b[92])^(a[3] & b[93])^(a[2] & b[94])^(a[1] & b[95])^(a[0] & b[96]);
assign y[97] = (a[97] & b[0])^(a[96] & b[1])^(a[95] & b[2])^(a[94] & b[3])^(a[93] & b[4])^(a[92] & b[5])^(a[91] & b[6])^(a[90] & b[7])^(a[89] & b[8])^(a[88] & b[9])^(a[87] & b[10])^(a[86] & b[11])^(a[85] & b[12])^(a[84] & b[13])^(a[83] & b[14])^(a[82] & b[15])^(a[81] & b[16])^(a[80] & b[17])^(a[79] & b[18])^(a[78] & b[19])^(a[77] & b[20])^(a[76] & b[21])^(a[75] & b[22])^(a[74] & b[23])^(a[73] & b[24])^(a[72] & b[25])^(a[71] & b[26])^(a[70] & b[27])^(a[69] & b[28])^(a[68] & b[29])^(a[67] & b[30])^(a[66] & b[31])^(a[65] & b[32])^(a[64] & b[33])^(a[63] & b[34])^(a[62] & b[35])^(a[61] & b[36])^(a[60] & b[37])^(a[59] & b[38])^(a[58] & b[39])^(a[57] & b[40])^(a[56] & b[41])^(a[55] & b[42])^(a[54] & b[43])^(a[53] & b[44])^(a[52] & b[45])^(a[51] & b[46])^(a[50] & b[47])^(a[49] & b[48])^(a[48] & b[49])^(a[47] & b[50])^(a[46] & b[51])^(a[45] & b[52])^(a[44] & b[53])^(a[43] & b[54])^(a[42] & b[55])^(a[41] & b[56])^(a[40] & b[57])^(a[39] & b[58])^(a[38] & b[59])^(a[37] & b[60])^(a[36] & b[61])^(a[35] & b[62])^(a[34] & b[63])^(a[33] & b[64])^(a[32] & b[65])^(a[31] & b[66])^(a[30] & b[67])^(a[29] & b[68])^(a[28] & b[69])^(a[27] & b[70])^(a[26] & b[71])^(a[25] & b[72])^(a[24] & b[73])^(a[23] & b[74])^(a[22] & b[75])^(a[21] & b[76])^(a[20] & b[77])^(a[19] & b[78])^(a[18] & b[79])^(a[17] & b[80])^(a[16] & b[81])^(a[15] & b[82])^(a[14] & b[83])^(a[13] & b[84])^(a[12] & b[85])^(a[11] & b[86])^(a[10] & b[87])^(a[9] & b[88])^(a[8] & b[89])^(a[7] & b[90])^(a[6] & b[91])^(a[5] & b[92])^(a[4] & b[93])^(a[3] & b[94])^(a[2] & b[95])^(a[1] & b[96])^(a[0] & b[97]);
assign y[98] = (a[98] & b[0])^(a[97] & b[1])^(a[96] & b[2])^(a[95] & b[3])^(a[94] & b[4])^(a[93] & b[5])^(a[92] & b[6])^(a[91] & b[7])^(a[90] & b[8])^(a[89] & b[9])^(a[88] & b[10])^(a[87] & b[11])^(a[86] & b[12])^(a[85] & b[13])^(a[84] & b[14])^(a[83] & b[15])^(a[82] & b[16])^(a[81] & b[17])^(a[80] & b[18])^(a[79] & b[19])^(a[78] & b[20])^(a[77] & b[21])^(a[76] & b[22])^(a[75] & b[23])^(a[74] & b[24])^(a[73] & b[25])^(a[72] & b[26])^(a[71] & b[27])^(a[70] & b[28])^(a[69] & b[29])^(a[68] & b[30])^(a[67] & b[31])^(a[66] & b[32])^(a[65] & b[33])^(a[64] & b[34])^(a[63] & b[35])^(a[62] & b[36])^(a[61] & b[37])^(a[60] & b[38])^(a[59] & b[39])^(a[58] & b[40])^(a[57] & b[41])^(a[56] & b[42])^(a[55] & b[43])^(a[54] & b[44])^(a[53] & b[45])^(a[52] & b[46])^(a[51] & b[47])^(a[50] & b[48])^(a[49] & b[49])^(a[48] & b[50])^(a[47] & b[51])^(a[46] & b[52])^(a[45] & b[53])^(a[44] & b[54])^(a[43] & b[55])^(a[42] & b[56])^(a[41] & b[57])^(a[40] & b[58])^(a[39] & b[59])^(a[38] & b[60])^(a[37] & b[61])^(a[36] & b[62])^(a[35] & b[63])^(a[34] & b[64])^(a[33] & b[65])^(a[32] & b[66])^(a[31] & b[67])^(a[30] & b[68])^(a[29] & b[69])^(a[28] & b[70])^(a[27] & b[71])^(a[26] & b[72])^(a[25] & b[73])^(a[24] & b[74])^(a[23] & b[75])^(a[22] & b[76])^(a[21] & b[77])^(a[20] & b[78])^(a[19] & b[79])^(a[18] & b[80])^(a[17] & b[81])^(a[16] & b[82])^(a[15] & b[83])^(a[14] & b[84])^(a[13] & b[85])^(a[12] & b[86])^(a[11] & b[87])^(a[10] & b[88])^(a[9] & b[89])^(a[8] & b[90])^(a[7] & b[91])^(a[6] & b[92])^(a[5] & b[93])^(a[4] & b[94])^(a[3] & b[95])^(a[2] & b[96])^(a[1] & b[97])^(a[0] & b[98]);
assign y[99] = (a[99] & b[0])^(a[98] & b[1])^(a[97] & b[2])^(a[96] & b[3])^(a[95] & b[4])^(a[94] & b[5])^(a[93] & b[6])^(a[92] & b[7])^(a[91] & b[8])^(a[90] & b[9])^(a[89] & b[10])^(a[88] & b[11])^(a[87] & b[12])^(a[86] & b[13])^(a[85] & b[14])^(a[84] & b[15])^(a[83] & b[16])^(a[82] & b[17])^(a[81] & b[18])^(a[80] & b[19])^(a[79] & b[20])^(a[78] & b[21])^(a[77] & b[22])^(a[76] & b[23])^(a[75] & b[24])^(a[74] & b[25])^(a[73] & b[26])^(a[72] & b[27])^(a[71] & b[28])^(a[70] & b[29])^(a[69] & b[30])^(a[68] & b[31])^(a[67] & b[32])^(a[66] & b[33])^(a[65] & b[34])^(a[64] & b[35])^(a[63] & b[36])^(a[62] & b[37])^(a[61] & b[38])^(a[60] & b[39])^(a[59] & b[40])^(a[58] & b[41])^(a[57] & b[42])^(a[56] & b[43])^(a[55] & b[44])^(a[54] & b[45])^(a[53] & b[46])^(a[52] & b[47])^(a[51] & b[48])^(a[50] & b[49])^(a[49] & b[50])^(a[48] & b[51])^(a[47] & b[52])^(a[46] & b[53])^(a[45] & b[54])^(a[44] & b[55])^(a[43] & b[56])^(a[42] & b[57])^(a[41] & b[58])^(a[40] & b[59])^(a[39] & b[60])^(a[38] & b[61])^(a[37] & b[62])^(a[36] & b[63])^(a[35] & b[64])^(a[34] & b[65])^(a[33] & b[66])^(a[32] & b[67])^(a[31] & b[68])^(a[30] & b[69])^(a[29] & b[70])^(a[28] & b[71])^(a[27] & b[72])^(a[26] & b[73])^(a[25] & b[74])^(a[24] & b[75])^(a[23] & b[76])^(a[22] & b[77])^(a[21] & b[78])^(a[20] & b[79])^(a[19] & b[80])^(a[18] & b[81])^(a[17] & b[82])^(a[16] & b[83])^(a[15] & b[84])^(a[14] & b[85])^(a[13] & b[86])^(a[12] & b[87])^(a[11] & b[88])^(a[10] & b[89])^(a[9] & b[90])^(a[8] & b[91])^(a[7] & b[92])^(a[6] & b[93])^(a[5] & b[94])^(a[4] & b[95])^(a[3] & b[96])^(a[2] & b[97])^(a[1] & b[98])^(a[0] & b[99]);
assign y[100] = (a[100] & b[0])^(a[99] & b[1])^(a[98] & b[2])^(a[97] & b[3])^(a[96] & b[4])^(a[95] & b[5])^(a[94] & b[6])^(a[93] & b[7])^(a[92] & b[8])^(a[91] & b[9])^(a[90] & b[10])^(a[89] & b[11])^(a[88] & b[12])^(a[87] & b[13])^(a[86] & b[14])^(a[85] & b[15])^(a[84] & b[16])^(a[83] & b[17])^(a[82] & b[18])^(a[81] & b[19])^(a[80] & b[20])^(a[79] & b[21])^(a[78] & b[22])^(a[77] & b[23])^(a[76] & b[24])^(a[75] & b[25])^(a[74] & b[26])^(a[73] & b[27])^(a[72] & b[28])^(a[71] & b[29])^(a[70] & b[30])^(a[69] & b[31])^(a[68] & b[32])^(a[67] & b[33])^(a[66] & b[34])^(a[65] & b[35])^(a[64] & b[36])^(a[63] & b[37])^(a[62] & b[38])^(a[61] & b[39])^(a[60] & b[40])^(a[59] & b[41])^(a[58] & b[42])^(a[57] & b[43])^(a[56] & b[44])^(a[55] & b[45])^(a[54] & b[46])^(a[53] & b[47])^(a[52] & b[48])^(a[51] & b[49])^(a[50] & b[50])^(a[49] & b[51])^(a[48] & b[52])^(a[47] & b[53])^(a[46] & b[54])^(a[45] & b[55])^(a[44] & b[56])^(a[43] & b[57])^(a[42] & b[58])^(a[41] & b[59])^(a[40] & b[60])^(a[39] & b[61])^(a[38] & b[62])^(a[37] & b[63])^(a[36] & b[64])^(a[35] & b[65])^(a[34] & b[66])^(a[33] & b[67])^(a[32] & b[68])^(a[31] & b[69])^(a[30] & b[70])^(a[29] & b[71])^(a[28] & b[72])^(a[27] & b[73])^(a[26] & b[74])^(a[25] & b[75])^(a[24] & b[76])^(a[23] & b[77])^(a[22] & b[78])^(a[21] & b[79])^(a[20] & b[80])^(a[19] & b[81])^(a[18] & b[82])^(a[17] & b[83])^(a[16] & b[84])^(a[15] & b[85])^(a[14] & b[86])^(a[13] & b[87])^(a[12] & b[88])^(a[11] & b[89])^(a[10] & b[90])^(a[9] & b[91])^(a[8] & b[92])^(a[7] & b[93])^(a[6] & b[94])^(a[5] & b[95])^(a[4] & b[96])^(a[3] & b[97])^(a[2] & b[98])^(a[1] & b[99])^(a[0] & b[100]);
assign y[101] = (a[101] & b[0])^(a[100] & b[1])^(a[99] & b[2])^(a[98] & b[3])^(a[97] & b[4])^(a[96] & b[5])^(a[95] & b[6])^(a[94] & b[7])^(a[93] & b[8])^(a[92] & b[9])^(a[91] & b[10])^(a[90] & b[11])^(a[89] & b[12])^(a[88] & b[13])^(a[87] & b[14])^(a[86] & b[15])^(a[85] & b[16])^(a[84] & b[17])^(a[83] & b[18])^(a[82] & b[19])^(a[81] & b[20])^(a[80] & b[21])^(a[79] & b[22])^(a[78] & b[23])^(a[77] & b[24])^(a[76] & b[25])^(a[75] & b[26])^(a[74] & b[27])^(a[73] & b[28])^(a[72] & b[29])^(a[71] & b[30])^(a[70] & b[31])^(a[69] & b[32])^(a[68] & b[33])^(a[67] & b[34])^(a[66] & b[35])^(a[65] & b[36])^(a[64] & b[37])^(a[63] & b[38])^(a[62] & b[39])^(a[61] & b[40])^(a[60] & b[41])^(a[59] & b[42])^(a[58] & b[43])^(a[57] & b[44])^(a[56] & b[45])^(a[55] & b[46])^(a[54] & b[47])^(a[53] & b[48])^(a[52] & b[49])^(a[51] & b[50])^(a[50] & b[51])^(a[49] & b[52])^(a[48] & b[53])^(a[47] & b[54])^(a[46] & b[55])^(a[45] & b[56])^(a[44] & b[57])^(a[43] & b[58])^(a[42] & b[59])^(a[41] & b[60])^(a[40] & b[61])^(a[39] & b[62])^(a[38] & b[63])^(a[37] & b[64])^(a[36] & b[65])^(a[35] & b[66])^(a[34] & b[67])^(a[33] & b[68])^(a[32] & b[69])^(a[31] & b[70])^(a[30] & b[71])^(a[29] & b[72])^(a[28] & b[73])^(a[27] & b[74])^(a[26] & b[75])^(a[25] & b[76])^(a[24] & b[77])^(a[23] & b[78])^(a[22] & b[79])^(a[21] & b[80])^(a[20] & b[81])^(a[19] & b[82])^(a[18] & b[83])^(a[17] & b[84])^(a[16] & b[85])^(a[15] & b[86])^(a[14] & b[87])^(a[13] & b[88])^(a[12] & b[89])^(a[11] & b[90])^(a[10] & b[91])^(a[9] & b[92])^(a[8] & b[93])^(a[7] & b[94])^(a[6] & b[95])^(a[5] & b[96])^(a[4] & b[97])^(a[3] & b[98])^(a[2] & b[99])^(a[1] & b[100])^(a[0] & b[101]);
assign y[102] = (a[102] & b[0])^(a[101] & b[1])^(a[100] & b[2])^(a[99] & b[3])^(a[98] & b[4])^(a[97] & b[5])^(a[96] & b[6])^(a[95] & b[7])^(a[94] & b[8])^(a[93] & b[9])^(a[92] & b[10])^(a[91] & b[11])^(a[90] & b[12])^(a[89] & b[13])^(a[88] & b[14])^(a[87] & b[15])^(a[86] & b[16])^(a[85] & b[17])^(a[84] & b[18])^(a[83] & b[19])^(a[82] & b[20])^(a[81] & b[21])^(a[80] & b[22])^(a[79] & b[23])^(a[78] & b[24])^(a[77] & b[25])^(a[76] & b[26])^(a[75] & b[27])^(a[74] & b[28])^(a[73] & b[29])^(a[72] & b[30])^(a[71] & b[31])^(a[70] & b[32])^(a[69] & b[33])^(a[68] & b[34])^(a[67] & b[35])^(a[66] & b[36])^(a[65] & b[37])^(a[64] & b[38])^(a[63] & b[39])^(a[62] & b[40])^(a[61] & b[41])^(a[60] & b[42])^(a[59] & b[43])^(a[58] & b[44])^(a[57] & b[45])^(a[56] & b[46])^(a[55] & b[47])^(a[54] & b[48])^(a[53] & b[49])^(a[52] & b[50])^(a[51] & b[51])^(a[50] & b[52])^(a[49] & b[53])^(a[48] & b[54])^(a[47] & b[55])^(a[46] & b[56])^(a[45] & b[57])^(a[44] & b[58])^(a[43] & b[59])^(a[42] & b[60])^(a[41] & b[61])^(a[40] & b[62])^(a[39] & b[63])^(a[38] & b[64])^(a[37] & b[65])^(a[36] & b[66])^(a[35] & b[67])^(a[34] & b[68])^(a[33] & b[69])^(a[32] & b[70])^(a[31] & b[71])^(a[30] & b[72])^(a[29] & b[73])^(a[28] & b[74])^(a[27] & b[75])^(a[26] & b[76])^(a[25] & b[77])^(a[24] & b[78])^(a[23] & b[79])^(a[22] & b[80])^(a[21] & b[81])^(a[20] & b[82])^(a[19] & b[83])^(a[18] & b[84])^(a[17] & b[85])^(a[16] & b[86])^(a[15] & b[87])^(a[14] & b[88])^(a[13] & b[89])^(a[12] & b[90])^(a[11] & b[91])^(a[10] & b[92])^(a[9] & b[93])^(a[8] & b[94])^(a[7] & b[95])^(a[6] & b[96])^(a[5] & b[97])^(a[4] & b[98])^(a[3] & b[99])^(a[2] & b[100])^(a[1] & b[101])^(a[0] & b[102]);
assign y[103] = (a[103] & b[0])^(a[102] & b[1])^(a[101] & b[2])^(a[100] & b[3])^(a[99] & b[4])^(a[98] & b[5])^(a[97] & b[6])^(a[96] & b[7])^(a[95] & b[8])^(a[94] & b[9])^(a[93] & b[10])^(a[92] & b[11])^(a[91] & b[12])^(a[90] & b[13])^(a[89] & b[14])^(a[88] & b[15])^(a[87] & b[16])^(a[86] & b[17])^(a[85] & b[18])^(a[84] & b[19])^(a[83] & b[20])^(a[82] & b[21])^(a[81] & b[22])^(a[80] & b[23])^(a[79] & b[24])^(a[78] & b[25])^(a[77] & b[26])^(a[76] & b[27])^(a[75] & b[28])^(a[74] & b[29])^(a[73] & b[30])^(a[72] & b[31])^(a[71] & b[32])^(a[70] & b[33])^(a[69] & b[34])^(a[68] & b[35])^(a[67] & b[36])^(a[66] & b[37])^(a[65] & b[38])^(a[64] & b[39])^(a[63] & b[40])^(a[62] & b[41])^(a[61] & b[42])^(a[60] & b[43])^(a[59] & b[44])^(a[58] & b[45])^(a[57] & b[46])^(a[56] & b[47])^(a[55] & b[48])^(a[54] & b[49])^(a[53] & b[50])^(a[52] & b[51])^(a[51] & b[52])^(a[50] & b[53])^(a[49] & b[54])^(a[48] & b[55])^(a[47] & b[56])^(a[46] & b[57])^(a[45] & b[58])^(a[44] & b[59])^(a[43] & b[60])^(a[42] & b[61])^(a[41] & b[62])^(a[40] & b[63])^(a[39] & b[64])^(a[38] & b[65])^(a[37] & b[66])^(a[36] & b[67])^(a[35] & b[68])^(a[34] & b[69])^(a[33] & b[70])^(a[32] & b[71])^(a[31] & b[72])^(a[30] & b[73])^(a[29] & b[74])^(a[28] & b[75])^(a[27] & b[76])^(a[26] & b[77])^(a[25] & b[78])^(a[24] & b[79])^(a[23] & b[80])^(a[22] & b[81])^(a[21] & b[82])^(a[20] & b[83])^(a[19] & b[84])^(a[18] & b[85])^(a[17] & b[86])^(a[16] & b[87])^(a[15] & b[88])^(a[14] & b[89])^(a[13] & b[90])^(a[12] & b[91])^(a[11] & b[92])^(a[10] & b[93])^(a[9] & b[94])^(a[8] & b[95])^(a[7] & b[96])^(a[6] & b[97])^(a[5] & b[98])^(a[4] & b[99])^(a[3] & b[100])^(a[2] & b[101])^(a[1] & b[102])^(a[0] & b[103]);
assign y[104] = (a[104] & b[0])^(a[103] & b[1])^(a[102] & b[2])^(a[101] & b[3])^(a[100] & b[4])^(a[99] & b[5])^(a[98] & b[6])^(a[97] & b[7])^(a[96] & b[8])^(a[95] & b[9])^(a[94] & b[10])^(a[93] & b[11])^(a[92] & b[12])^(a[91] & b[13])^(a[90] & b[14])^(a[89] & b[15])^(a[88] & b[16])^(a[87] & b[17])^(a[86] & b[18])^(a[85] & b[19])^(a[84] & b[20])^(a[83] & b[21])^(a[82] & b[22])^(a[81] & b[23])^(a[80] & b[24])^(a[79] & b[25])^(a[78] & b[26])^(a[77] & b[27])^(a[76] & b[28])^(a[75] & b[29])^(a[74] & b[30])^(a[73] & b[31])^(a[72] & b[32])^(a[71] & b[33])^(a[70] & b[34])^(a[69] & b[35])^(a[68] & b[36])^(a[67] & b[37])^(a[66] & b[38])^(a[65] & b[39])^(a[64] & b[40])^(a[63] & b[41])^(a[62] & b[42])^(a[61] & b[43])^(a[60] & b[44])^(a[59] & b[45])^(a[58] & b[46])^(a[57] & b[47])^(a[56] & b[48])^(a[55] & b[49])^(a[54] & b[50])^(a[53] & b[51])^(a[52] & b[52])^(a[51] & b[53])^(a[50] & b[54])^(a[49] & b[55])^(a[48] & b[56])^(a[47] & b[57])^(a[46] & b[58])^(a[45] & b[59])^(a[44] & b[60])^(a[43] & b[61])^(a[42] & b[62])^(a[41] & b[63])^(a[40] & b[64])^(a[39] & b[65])^(a[38] & b[66])^(a[37] & b[67])^(a[36] & b[68])^(a[35] & b[69])^(a[34] & b[70])^(a[33] & b[71])^(a[32] & b[72])^(a[31] & b[73])^(a[30] & b[74])^(a[29] & b[75])^(a[28] & b[76])^(a[27] & b[77])^(a[26] & b[78])^(a[25] & b[79])^(a[24] & b[80])^(a[23] & b[81])^(a[22] & b[82])^(a[21] & b[83])^(a[20] & b[84])^(a[19] & b[85])^(a[18] & b[86])^(a[17] & b[87])^(a[16] & b[88])^(a[15] & b[89])^(a[14] & b[90])^(a[13] & b[91])^(a[12] & b[92])^(a[11] & b[93])^(a[10] & b[94])^(a[9] & b[95])^(a[8] & b[96])^(a[7] & b[97])^(a[6] & b[98])^(a[5] & b[99])^(a[4] & b[100])^(a[3] & b[101])^(a[2] & b[102])^(a[1] & b[103])^(a[0] & b[104]);
assign y[105] = (a[105] & b[0])^(a[104] & b[1])^(a[103] & b[2])^(a[102] & b[3])^(a[101] & b[4])^(a[100] & b[5])^(a[99] & b[6])^(a[98] & b[7])^(a[97] & b[8])^(a[96] & b[9])^(a[95] & b[10])^(a[94] & b[11])^(a[93] & b[12])^(a[92] & b[13])^(a[91] & b[14])^(a[90] & b[15])^(a[89] & b[16])^(a[88] & b[17])^(a[87] & b[18])^(a[86] & b[19])^(a[85] & b[20])^(a[84] & b[21])^(a[83] & b[22])^(a[82] & b[23])^(a[81] & b[24])^(a[80] & b[25])^(a[79] & b[26])^(a[78] & b[27])^(a[77] & b[28])^(a[76] & b[29])^(a[75] & b[30])^(a[74] & b[31])^(a[73] & b[32])^(a[72] & b[33])^(a[71] & b[34])^(a[70] & b[35])^(a[69] & b[36])^(a[68] & b[37])^(a[67] & b[38])^(a[66] & b[39])^(a[65] & b[40])^(a[64] & b[41])^(a[63] & b[42])^(a[62] & b[43])^(a[61] & b[44])^(a[60] & b[45])^(a[59] & b[46])^(a[58] & b[47])^(a[57] & b[48])^(a[56] & b[49])^(a[55] & b[50])^(a[54] & b[51])^(a[53] & b[52])^(a[52] & b[53])^(a[51] & b[54])^(a[50] & b[55])^(a[49] & b[56])^(a[48] & b[57])^(a[47] & b[58])^(a[46] & b[59])^(a[45] & b[60])^(a[44] & b[61])^(a[43] & b[62])^(a[42] & b[63])^(a[41] & b[64])^(a[40] & b[65])^(a[39] & b[66])^(a[38] & b[67])^(a[37] & b[68])^(a[36] & b[69])^(a[35] & b[70])^(a[34] & b[71])^(a[33] & b[72])^(a[32] & b[73])^(a[31] & b[74])^(a[30] & b[75])^(a[29] & b[76])^(a[28] & b[77])^(a[27] & b[78])^(a[26] & b[79])^(a[25] & b[80])^(a[24] & b[81])^(a[23] & b[82])^(a[22] & b[83])^(a[21] & b[84])^(a[20] & b[85])^(a[19] & b[86])^(a[18] & b[87])^(a[17] & b[88])^(a[16] & b[89])^(a[15] & b[90])^(a[14] & b[91])^(a[13] & b[92])^(a[12] & b[93])^(a[11] & b[94])^(a[10] & b[95])^(a[9] & b[96])^(a[8] & b[97])^(a[7] & b[98])^(a[6] & b[99])^(a[5] & b[100])^(a[4] & b[101])^(a[3] & b[102])^(a[2] & b[103])^(a[1] & b[104])^(a[0] & b[105]);
assign y[106] = (a[106] & b[0])^(a[105] & b[1])^(a[104] & b[2])^(a[103] & b[3])^(a[102] & b[4])^(a[101] & b[5])^(a[100] & b[6])^(a[99] & b[7])^(a[98] & b[8])^(a[97] & b[9])^(a[96] & b[10])^(a[95] & b[11])^(a[94] & b[12])^(a[93] & b[13])^(a[92] & b[14])^(a[91] & b[15])^(a[90] & b[16])^(a[89] & b[17])^(a[88] & b[18])^(a[87] & b[19])^(a[86] & b[20])^(a[85] & b[21])^(a[84] & b[22])^(a[83] & b[23])^(a[82] & b[24])^(a[81] & b[25])^(a[80] & b[26])^(a[79] & b[27])^(a[78] & b[28])^(a[77] & b[29])^(a[76] & b[30])^(a[75] & b[31])^(a[74] & b[32])^(a[73] & b[33])^(a[72] & b[34])^(a[71] & b[35])^(a[70] & b[36])^(a[69] & b[37])^(a[68] & b[38])^(a[67] & b[39])^(a[66] & b[40])^(a[65] & b[41])^(a[64] & b[42])^(a[63] & b[43])^(a[62] & b[44])^(a[61] & b[45])^(a[60] & b[46])^(a[59] & b[47])^(a[58] & b[48])^(a[57] & b[49])^(a[56] & b[50])^(a[55] & b[51])^(a[54] & b[52])^(a[53] & b[53])^(a[52] & b[54])^(a[51] & b[55])^(a[50] & b[56])^(a[49] & b[57])^(a[48] & b[58])^(a[47] & b[59])^(a[46] & b[60])^(a[45] & b[61])^(a[44] & b[62])^(a[43] & b[63])^(a[42] & b[64])^(a[41] & b[65])^(a[40] & b[66])^(a[39] & b[67])^(a[38] & b[68])^(a[37] & b[69])^(a[36] & b[70])^(a[35] & b[71])^(a[34] & b[72])^(a[33] & b[73])^(a[32] & b[74])^(a[31] & b[75])^(a[30] & b[76])^(a[29] & b[77])^(a[28] & b[78])^(a[27] & b[79])^(a[26] & b[80])^(a[25] & b[81])^(a[24] & b[82])^(a[23] & b[83])^(a[22] & b[84])^(a[21] & b[85])^(a[20] & b[86])^(a[19] & b[87])^(a[18] & b[88])^(a[17] & b[89])^(a[16] & b[90])^(a[15] & b[91])^(a[14] & b[92])^(a[13] & b[93])^(a[12] & b[94])^(a[11] & b[95])^(a[10] & b[96])^(a[9] & b[97])^(a[8] & b[98])^(a[7] & b[99])^(a[6] & b[100])^(a[5] & b[101])^(a[4] & b[102])^(a[3] & b[103])^(a[2] & b[104])^(a[1] & b[105])^(a[0] & b[106]);
assign y[107] = (a[107] & b[0])^(a[106] & b[1])^(a[105] & b[2])^(a[104] & b[3])^(a[103] & b[4])^(a[102] & b[5])^(a[101] & b[6])^(a[100] & b[7])^(a[99] & b[8])^(a[98] & b[9])^(a[97] & b[10])^(a[96] & b[11])^(a[95] & b[12])^(a[94] & b[13])^(a[93] & b[14])^(a[92] & b[15])^(a[91] & b[16])^(a[90] & b[17])^(a[89] & b[18])^(a[88] & b[19])^(a[87] & b[20])^(a[86] & b[21])^(a[85] & b[22])^(a[84] & b[23])^(a[83] & b[24])^(a[82] & b[25])^(a[81] & b[26])^(a[80] & b[27])^(a[79] & b[28])^(a[78] & b[29])^(a[77] & b[30])^(a[76] & b[31])^(a[75] & b[32])^(a[74] & b[33])^(a[73] & b[34])^(a[72] & b[35])^(a[71] & b[36])^(a[70] & b[37])^(a[69] & b[38])^(a[68] & b[39])^(a[67] & b[40])^(a[66] & b[41])^(a[65] & b[42])^(a[64] & b[43])^(a[63] & b[44])^(a[62] & b[45])^(a[61] & b[46])^(a[60] & b[47])^(a[59] & b[48])^(a[58] & b[49])^(a[57] & b[50])^(a[56] & b[51])^(a[55] & b[52])^(a[54] & b[53])^(a[53] & b[54])^(a[52] & b[55])^(a[51] & b[56])^(a[50] & b[57])^(a[49] & b[58])^(a[48] & b[59])^(a[47] & b[60])^(a[46] & b[61])^(a[45] & b[62])^(a[44] & b[63])^(a[43] & b[64])^(a[42] & b[65])^(a[41] & b[66])^(a[40] & b[67])^(a[39] & b[68])^(a[38] & b[69])^(a[37] & b[70])^(a[36] & b[71])^(a[35] & b[72])^(a[34] & b[73])^(a[33] & b[74])^(a[32] & b[75])^(a[31] & b[76])^(a[30] & b[77])^(a[29] & b[78])^(a[28] & b[79])^(a[27] & b[80])^(a[26] & b[81])^(a[25] & b[82])^(a[24] & b[83])^(a[23] & b[84])^(a[22] & b[85])^(a[21] & b[86])^(a[20] & b[87])^(a[19] & b[88])^(a[18] & b[89])^(a[17] & b[90])^(a[16] & b[91])^(a[15] & b[92])^(a[14] & b[93])^(a[13] & b[94])^(a[12] & b[95])^(a[11] & b[96])^(a[10] & b[97])^(a[9] & b[98])^(a[8] & b[99])^(a[7] & b[100])^(a[6] & b[101])^(a[5] & b[102])^(a[4] & b[103])^(a[3] & b[104])^(a[2] & b[105])^(a[1] & b[106])^(a[0] & b[107]);
assign y[108] = (a[108] & b[0])^(a[107] & b[1])^(a[106] & b[2])^(a[105] & b[3])^(a[104] & b[4])^(a[103] & b[5])^(a[102] & b[6])^(a[101] & b[7])^(a[100] & b[8])^(a[99] & b[9])^(a[98] & b[10])^(a[97] & b[11])^(a[96] & b[12])^(a[95] & b[13])^(a[94] & b[14])^(a[93] & b[15])^(a[92] & b[16])^(a[91] & b[17])^(a[90] & b[18])^(a[89] & b[19])^(a[88] & b[20])^(a[87] & b[21])^(a[86] & b[22])^(a[85] & b[23])^(a[84] & b[24])^(a[83] & b[25])^(a[82] & b[26])^(a[81] & b[27])^(a[80] & b[28])^(a[79] & b[29])^(a[78] & b[30])^(a[77] & b[31])^(a[76] & b[32])^(a[75] & b[33])^(a[74] & b[34])^(a[73] & b[35])^(a[72] & b[36])^(a[71] & b[37])^(a[70] & b[38])^(a[69] & b[39])^(a[68] & b[40])^(a[67] & b[41])^(a[66] & b[42])^(a[65] & b[43])^(a[64] & b[44])^(a[63] & b[45])^(a[62] & b[46])^(a[61] & b[47])^(a[60] & b[48])^(a[59] & b[49])^(a[58] & b[50])^(a[57] & b[51])^(a[56] & b[52])^(a[55] & b[53])^(a[54] & b[54])^(a[53] & b[55])^(a[52] & b[56])^(a[51] & b[57])^(a[50] & b[58])^(a[49] & b[59])^(a[48] & b[60])^(a[47] & b[61])^(a[46] & b[62])^(a[45] & b[63])^(a[44] & b[64])^(a[43] & b[65])^(a[42] & b[66])^(a[41] & b[67])^(a[40] & b[68])^(a[39] & b[69])^(a[38] & b[70])^(a[37] & b[71])^(a[36] & b[72])^(a[35] & b[73])^(a[34] & b[74])^(a[33] & b[75])^(a[32] & b[76])^(a[31] & b[77])^(a[30] & b[78])^(a[29] & b[79])^(a[28] & b[80])^(a[27] & b[81])^(a[26] & b[82])^(a[25] & b[83])^(a[24] & b[84])^(a[23] & b[85])^(a[22] & b[86])^(a[21] & b[87])^(a[20] & b[88])^(a[19] & b[89])^(a[18] & b[90])^(a[17] & b[91])^(a[16] & b[92])^(a[15] & b[93])^(a[14] & b[94])^(a[13] & b[95])^(a[12] & b[96])^(a[11] & b[97])^(a[10] & b[98])^(a[9] & b[99])^(a[8] & b[100])^(a[7] & b[101])^(a[6] & b[102])^(a[5] & b[103])^(a[4] & b[104])^(a[3] & b[105])^(a[2] & b[106])^(a[1] & b[107])^(a[0] & b[108]);
assign y[109] = (a[109] & b[0])^(a[108] & b[1])^(a[107] & b[2])^(a[106] & b[3])^(a[105] & b[4])^(a[104] & b[5])^(a[103] & b[6])^(a[102] & b[7])^(a[101] & b[8])^(a[100] & b[9])^(a[99] & b[10])^(a[98] & b[11])^(a[97] & b[12])^(a[96] & b[13])^(a[95] & b[14])^(a[94] & b[15])^(a[93] & b[16])^(a[92] & b[17])^(a[91] & b[18])^(a[90] & b[19])^(a[89] & b[20])^(a[88] & b[21])^(a[87] & b[22])^(a[86] & b[23])^(a[85] & b[24])^(a[84] & b[25])^(a[83] & b[26])^(a[82] & b[27])^(a[81] & b[28])^(a[80] & b[29])^(a[79] & b[30])^(a[78] & b[31])^(a[77] & b[32])^(a[76] & b[33])^(a[75] & b[34])^(a[74] & b[35])^(a[73] & b[36])^(a[72] & b[37])^(a[71] & b[38])^(a[70] & b[39])^(a[69] & b[40])^(a[68] & b[41])^(a[67] & b[42])^(a[66] & b[43])^(a[65] & b[44])^(a[64] & b[45])^(a[63] & b[46])^(a[62] & b[47])^(a[61] & b[48])^(a[60] & b[49])^(a[59] & b[50])^(a[58] & b[51])^(a[57] & b[52])^(a[56] & b[53])^(a[55] & b[54])^(a[54] & b[55])^(a[53] & b[56])^(a[52] & b[57])^(a[51] & b[58])^(a[50] & b[59])^(a[49] & b[60])^(a[48] & b[61])^(a[47] & b[62])^(a[46] & b[63])^(a[45] & b[64])^(a[44] & b[65])^(a[43] & b[66])^(a[42] & b[67])^(a[41] & b[68])^(a[40] & b[69])^(a[39] & b[70])^(a[38] & b[71])^(a[37] & b[72])^(a[36] & b[73])^(a[35] & b[74])^(a[34] & b[75])^(a[33] & b[76])^(a[32] & b[77])^(a[31] & b[78])^(a[30] & b[79])^(a[29] & b[80])^(a[28] & b[81])^(a[27] & b[82])^(a[26] & b[83])^(a[25] & b[84])^(a[24] & b[85])^(a[23] & b[86])^(a[22] & b[87])^(a[21] & b[88])^(a[20] & b[89])^(a[19] & b[90])^(a[18] & b[91])^(a[17] & b[92])^(a[16] & b[93])^(a[15] & b[94])^(a[14] & b[95])^(a[13] & b[96])^(a[12] & b[97])^(a[11] & b[98])^(a[10] & b[99])^(a[9] & b[100])^(a[8] & b[101])^(a[7] & b[102])^(a[6] & b[103])^(a[5] & b[104])^(a[4] & b[105])^(a[3] & b[106])^(a[2] & b[107])^(a[1] & b[108])^(a[0] & b[109]);
assign y[110] = (a[110] & b[0])^(a[109] & b[1])^(a[108] & b[2])^(a[107] & b[3])^(a[106] & b[4])^(a[105] & b[5])^(a[104] & b[6])^(a[103] & b[7])^(a[102] & b[8])^(a[101] & b[9])^(a[100] & b[10])^(a[99] & b[11])^(a[98] & b[12])^(a[97] & b[13])^(a[96] & b[14])^(a[95] & b[15])^(a[94] & b[16])^(a[93] & b[17])^(a[92] & b[18])^(a[91] & b[19])^(a[90] & b[20])^(a[89] & b[21])^(a[88] & b[22])^(a[87] & b[23])^(a[86] & b[24])^(a[85] & b[25])^(a[84] & b[26])^(a[83] & b[27])^(a[82] & b[28])^(a[81] & b[29])^(a[80] & b[30])^(a[79] & b[31])^(a[78] & b[32])^(a[77] & b[33])^(a[76] & b[34])^(a[75] & b[35])^(a[74] & b[36])^(a[73] & b[37])^(a[72] & b[38])^(a[71] & b[39])^(a[70] & b[40])^(a[69] & b[41])^(a[68] & b[42])^(a[67] & b[43])^(a[66] & b[44])^(a[65] & b[45])^(a[64] & b[46])^(a[63] & b[47])^(a[62] & b[48])^(a[61] & b[49])^(a[60] & b[50])^(a[59] & b[51])^(a[58] & b[52])^(a[57] & b[53])^(a[56] & b[54])^(a[55] & b[55])^(a[54] & b[56])^(a[53] & b[57])^(a[52] & b[58])^(a[51] & b[59])^(a[50] & b[60])^(a[49] & b[61])^(a[48] & b[62])^(a[47] & b[63])^(a[46] & b[64])^(a[45] & b[65])^(a[44] & b[66])^(a[43] & b[67])^(a[42] & b[68])^(a[41] & b[69])^(a[40] & b[70])^(a[39] & b[71])^(a[38] & b[72])^(a[37] & b[73])^(a[36] & b[74])^(a[35] & b[75])^(a[34] & b[76])^(a[33] & b[77])^(a[32] & b[78])^(a[31] & b[79])^(a[30] & b[80])^(a[29] & b[81])^(a[28] & b[82])^(a[27] & b[83])^(a[26] & b[84])^(a[25] & b[85])^(a[24] & b[86])^(a[23] & b[87])^(a[22] & b[88])^(a[21] & b[89])^(a[20] & b[90])^(a[19] & b[91])^(a[18] & b[92])^(a[17] & b[93])^(a[16] & b[94])^(a[15] & b[95])^(a[14] & b[96])^(a[13] & b[97])^(a[12] & b[98])^(a[11] & b[99])^(a[10] & b[100])^(a[9] & b[101])^(a[8] & b[102])^(a[7] & b[103])^(a[6] & b[104])^(a[5] & b[105])^(a[4] & b[106])^(a[3] & b[107])^(a[2] & b[108])^(a[1] & b[109])^(a[0] & b[110]);
assign y[111] = (a[111] & b[0])^(a[110] & b[1])^(a[109] & b[2])^(a[108] & b[3])^(a[107] & b[4])^(a[106] & b[5])^(a[105] & b[6])^(a[104] & b[7])^(a[103] & b[8])^(a[102] & b[9])^(a[101] & b[10])^(a[100] & b[11])^(a[99] & b[12])^(a[98] & b[13])^(a[97] & b[14])^(a[96] & b[15])^(a[95] & b[16])^(a[94] & b[17])^(a[93] & b[18])^(a[92] & b[19])^(a[91] & b[20])^(a[90] & b[21])^(a[89] & b[22])^(a[88] & b[23])^(a[87] & b[24])^(a[86] & b[25])^(a[85] & b[26])^(a[84] & b[27])^(a[83] & b[28])^(a[82] & b[29])^(a[81] & b[30])^(a[80] & b[31])^(a[79] & b[32])^(a[78] & b[33])^(a[77] & b[34])^(a[76] & b[35])^(a[75] & b[36])^(a[74] & b[37])^(a[73] & b[38])^(a[72] & b[39])^(a[71] & b[40])^(a[70] & b[41])^(a[69] & b[42])^(a[68] & b[43])^(a[67] & b[44])^(a[66] & b[45])^(a[65] & b[46])^(a[64] & b[47])^(a[63] & b[48])^(a[62] & b[49])^(a[61] & b[50])^(a[60] & b[51])^(a[59] & b[52])^(a[58] & b[53])^(a[57] & b[54])^(a[56] & b[55])^(a[55] & b[56])^(a[54] & b[57])^(a[53] & b[58])^(a[52] & b[59])^(a[51] & b[60])^(a[50] & b[61])^(a[49] & b[62])^(a[48] & b[63])^(a[47] & b[64])^(a[46] & b[65])^(a[45] & b[66])^(a[44] & b[67])^(a[43] & b[68])^(a[42] & b[69])^(a[41] & b[70])^(a[40] & b[71])^(a[39] & b[72])^(a[38] & b[73])^(a[37] & b[74])^(a[36] & b[75])^(a[35] & b[76])^(a[34] & b[77])^(a[33] & b[78])^(a[32] & b[79])^(a[31] & b[80])^(a[30] & b[81])^(a[29] & b[82])^(a[28] & b[83])^(a[27] & b[84])^(a[26] & b[85])^(a[25] & b[86])^(a[24] & b[87])^(a[23] & b[88])^(a[22] & b[89])^(a[21] & b[90])^(a[20] & b[91])^(a[19] & b[92])^(a[18] & b[93])^(a[17] & b[94])^(a[16] & b[95])^(a[15] & b[96])^(a[14] & b[97])^(a[13] & b[98])^(a[12] & b[99])^(a[11] & b[100])^(a[10] & b[101])^(a[9] & b[102])^(a[8] & b[103])^(a[7] & b[104])^(a[6] & b[105])^(a[5] & b[106])^(a[4] & b[107])^(a[3] & b[108])^(a[2] & b[109])^(a[1] & b[110])^(a[0] & b[111]);
assign y[112] = (a[112] & b[0])^(a[111] & b[1])^(a[110] & b[2])^(a[109] & b[3])^(a[108] & b[4])^(a[107] & b[5])^(a[106] & b[6])^(a[105] & b[7])^(a[104] & b[8])^(a[103] & b[9])^(a[102] & b[10])^(a[101] & b[11])^(a[100] & b[12])^(a[99] & b[13])^(a[98] & b[14])^(a[97] & b[15])^(a[96] & b[16])^(a[95] & b[17])^(a[94] & b[18])^(a[93] & b[19])^(a[92] & b[20])^(a[91] & b[21])^(a[90] & b[22])^(a[89] & b[23])^(a[88] & b[24])^(a[87] & b[25])^(a[86] & b[26])^(a[85] & b[27])^(a[84] & b[28])^(a[83] & b[29])^(a[82] & b[30])^(a[81] & b[31])^(a[80] & b[32])^(a[79] & b[33])^(a[78] & b[34])^(a[77] & b[35])^(a[76] & b[36])^(a[75] & b[37])^(a[74] & b[38])^(a[73] & b[39])^(a[72] & b[40])^(a[71] & b[41])^(a[70] & b[42])^(a[69] & b[43])^(a[68] & b[44])^(a[67] & b[45])^(a[66] & b[46])^(a[65] & b[47])^(a[64] & b[48])^(a[63] & b[49])^(a[62] & b[50])^(a[61] & b[51])^(a[60] & b[52])^(a[59] & b[53])^(a[58] & b[54])^(a[57] & b[55])^(a[56] & b[56])^(a[55] & b[57])^(a[54] & b[58])^(a[53] & b[59])^(a[52] & b[60])^(a[51] & b[61])^(a[50] & b[62])^(a[49] & b[63])^(a[48] & b[64])^(a[47] & b[65])^(a[46] & b[66])^(a[45] & b[67])^(a[44] & b[68])^(a[43] & b[69])^(a[42] & b[70])^(a[41] & b[71])^(a[40] & b[72])^(a[39] & b[73])^(a[38] & b[74])^(a[37] & b[75])^(a[36] & b[76])^(a[35] & b[77])^(a[34] & b[78])^(a[33] & b[79])^(a[32] & b[80])^(a[31] & b[81])^(a[30] & b[82])^(a[29] & b[83])^(a[28] & b[84])^(a[27] & b[85])^(a[26] & b[86])^(a[25] & b[87])^(a[24] & b[88])^(a[23] & b[89])^(a[22] & b[90])^(a[21] & b[91])^(a[20] & b[92])^(a[19] & b[93])^(a[18] & b[94])^(a[17] & b[95])^(a[16] & b[96])^(a[15] & b[97])^(a[14] & b[98])^(a[13] & b[99])^(a[12] & b[100])^(a[11] & b[101])^(a[10] & b[102])^(a[9] & b[103])^(a[8] & b[104])^(a[7] & b[105])^(a[6] & b[106])^(a[5] & b[107])^(a[4] & b[108])^(a[3] & b[109])^(a[2] & b[110])^(a[1] & b[111])^(a[0] & b[112]);
assign y[113] = (a[113] & b[0])^(a[112] & b[1])^(a[111] & b[2])^(a[110] & b[3])^(a[109] & b[4])^(a[108] & b[5])^(a[107] & b[6])^(a[106] & b[7])^(a[105] & b[8])^(a[104] & b[9])^(a[103] & b[10])^(a[102] & b[11])^(a[101] & b[12])^(a[100] & b[13])^(a[99] & b[14])^(a[98] & b[15])^(a[97] & b[16])^(a[96] & b[17])^(a[95] & b[18])^(a[94] & b[19])^(a[93] & b[20])^(a[92] & b[21])^(a[91] & b[22])^(a[90] & b[23])^(a[89] & b[24])^(a[88] & b[25])^(a[87] & b[26])^(a[86] & b[27])^(a[85] & b[28])^(a[84] & b[29])^(a[83] & b[30])^(a[82] & b[31])^(a[81] & b[32])^(a[80] & b[33])^(a[79] & b[34])^(a[78] & b[35])^(a[77] & b[36])^(a[76] & b[37])^(a[75] & b[38])^(a[74] & b[39])^(a[73] & b[40])^(a[72] & b[41])^(a[71] & b[42])^(a[70] & b[43])^(a[69] & b[44])^(a[68] & b[45])^(a[67] & b[46])^(a[66] & b[47])^(a[65] & b[48])^(a[64] & b[49])^(a[63] & b[50])^(a[62] & b[51])^(a[61] & b[52])^(a[60] & b[53])^(a[59] & b[54])^(a[58] & b[55])^(a[57] & b[56])^(a[56] & b[57])^(a[55] & b[58])^(a[54] & b[59])^(a[53] & b[60])^(a[52] & b[61])^(a[51] & b[62])^(a[50] & b[63])^(a[49] & b[64])^(a[48] & b[65])^(a[47] & b[66])^(a[46] & b[67])^(a[45] & b[68])^(a[44] & b[69])^(a[43] & b[70])^(a[42] & b[71])^(a[41] & b[72])^(a[40] & b[73])^(a[39] & b[74])^(a[38] & b[75])^(a[37] & b[76])^(a[36] & b[77])^(a[35] & b[78])^(a[34] & b[79])^(a[33] & b[80])^(a[32] & b[81])^(a[31] & b[82])^(a[30] & b[83])^(a[29] & b[84])^(a[28] & b[85])^(a[27] & b[86])^(a[26] & b[87])^(a[25] & b[88])^(a[24] & b[89])^(a[23] & b[90])^(a[22] & b[91])^(a[21] & b[92])^(a[20] & b[93])^(a[19] & b[94])^(a[18] & b[95])^(a[17] & b[96])^(a[16] & b[97])^(a[15] & b[98])^(a[14] & b[99])^(a[13] & b[100])^(a[12] & b[101])^(a[11] & b[102])^(a[10] & b[103])^(a[9] & b[104])^(a[8] & b[105])^(a[7] & b[106])^(a[6] & b[107])^(a[5] & b[108])^(a[4] & b[109])^(a[3] & b[110])^(a[2] & b[111])^(a[1] & b[112])^(a[0] & b[113]);
assign y[114] = (a[114] & b[0])^(a[113] & b[1])^(a[112] & b[2])^(a[111] & b[3])^(a[110] & b[4])^(a[109] & b[5])^(a[108] & b[6])^(a[107] & b[7])^(a[106] & b[8])^(a[105] & b[9])^(a[104] & b[10])^(a[103] & b[11])^(a[102] & b[12])^(a[101] & b[13])^(a[100] & b[14])^(a[99] & b[15])^(a[98] & b[16])^(a[97] & b[17])^(a[96] & b[18])^(a[95] & b[19])^(a[94] & b[20])^(a[93] & b[21])^(a[92] & b[22])^(a[91] & b[23])^(a[90] & b[24])^(a[89] & b[25])^(a[88] & b[26])^(a[87] & b[27])^(a[86] & b[28])^(a[85] & b[29])^(a[84] & b[30])^(a[83] & b[31])^(a[82] & b[32])^(a[81] & b[33])^(a[80] & b[34])^(a[79] & b[35])^(a[78] & b[36])^(a[77] & b[37])^(a[76] & b[38])^(a[75] & b[39])^(a[74] & b[40])^(a[73] & b[41])^(a[72] & b[42])^(a[71] & b[43])^(a[70] & b[44])^(a[69] & b[45])^(a[68] & b[46])^(a[67] & b[47])^(a[66] & b[48])^(a[65] & b[49])^(a[64] & b[50])^(a[63] & b[51])^(a[62] & b[52])^(a[61] & b[53])^(a[60] & b[54])^(a[59] & b[55])^(a[58] & b[56])^(a[57] & b[57])^(a[56] & b[58])^(a[55] & b[59])^(a[54] & b[60])^(a[53] & b[61])^(a[52] & b[62])^(a[51] & b[63])^(a[50] & b[64])^(a[49] & b[65])^(a[48] & b[66])^(a[47] & b[67])^(a[46] & b[68])^(a[45] & b[69])^(a[44] & b[70])^(a[43] & b[71])^(a[42] & b[72])^(a[41] & b[73])^(a[40] & b[74])^(a[39] & b[75])^(a[38] & b[76])^(a[37] & b[77])^(a[36] & b[78])^(a[35] & b[79])^(a[34] & b[80])^(a[33] & b[81])^(a[32] & b[82])^(a[31] & b[83])^(a[30] & b[84])^(a[29] & b[85])^(a[28] & b[86])^(a[27] & b[87])^(a[26] & b[88])^(a[25] & b[89])^(a[24] & b[90])^(a[23] & b[91])^(a[22] & b[92])^(a[21] & b[93])^(a[20] & b[94])^(a[19] & b[95])^(a[18] & b[96])^(a[17] & b[97])^(a[16] & b[98])^(a[15] & b[99])^(a[14] & b[100])^(a[13] & b[101])^(a[12] & b[102])^(a[11] & b[103])^(a[10] & b[104])^(a[9] & b[105])^(a[8] & b[106])^(a[7] & b[107])^(a[6] & b[108])^(a[5] & b[109])^(a[4] & b[110])^(a[3] & b[111])^(a[2] & b[112])^(a[1] & b[113])^(a[0] & b[114]);
assign y[115] = (a[115] & b[0])^(a[114] & b[1])^(a[113] & b[2])^(a[112] & b[3])^(a[111] & b[4])^(a[110] & b[5])^(a[109] & b[6])^(a[108] & b[7])^(a[107] & b[8])^(a[106] & b[9])^(a[105] & b[10])^(a[104] & b[11])^(a[103] & b[12])^(a[102] & b[13])^(a[101] & b[14])^(a[100] & b[15])^(a[99] & b[16])^(a[98] & b[17])^(a[97] & b[18])^(a[96] & b[19])^(a[95] & b[20])^(a[94] & b[21])^(a[93] & b[22])^(a[92] & b[23])^(a[91] & b[24])^(a[90] & b[25])^(a[89] & b[26])^(a[88] & b[27])^(a[87] & b[28])^(a[86] & b[29])^(a[85] & b[30])^(a[84] & b[31])^(a[83] & b[32])^(a[82] & b[33])^(a[81] & b[34])^(a[80] & b[35])^(a[79] & b[36])^(a[78] & b[37])^(a[77] & b[38])^(a[76] & b[39])^(a[75] & b[40])^(a[74] & b[41])^(a[73] & b[42])^(a[72] & b[43])^(a[71] & b[44])^(a[70] & b[45])^(a[69] & b[46])^(a[68] & b[47])^(a[67] & b[48])^(a[66] & b[49])^(a[65] & b[50])^(a[64] & b[51])^(a[63] & b[52])^(a[62] & b[53])^(a[61] & b[54])^(a[60] & b[55])^(a[59] & b[56])^(a[58] & b[57])^(a[57] & b[58])^(a[56] & b[59])^(a[55] & b[60])^(a[54] & b[61])^(a[53] & b[62])^(a[52] & b[63])^(a[51] & b[64])^(a[50] & b[65])^(a[49] & b[66])^(a[48] & b[67])^(a[47] & b[68])^(a[46] & b[69])^(a[45] & b[70])^(a[44] & b[71])^(a[43] & b[72])^(a[42] & b[73])^(a[41] & b[74])^(a[40] & b[75])^(a[39] & b[76])^(a[38] & b[77])^(a[37] & b[78])^(a[36] & b[79])^(a[35] & b[80])^(a[34] & b[81])^(a[33] & b[82])^(a[32] & b[83])^(a[31] & b[84])^(a[30] & b[85])^(a[29] & b[86])^(a[28] & b[87])^(a[27] & b[88])^(a[26] & b[89])^(a[25] & b[90])^(a[24] & b[91])^(a[23] & b[92])^(a[22] & b[93])^(a[21] & b[94])^(a[20] & b[95])^(a[19] & b[96])^(a[18] & b[97])^(a[17] & b[98])^(a[16] & b[99])^(a[15] & b[100])^(a[14] & b[101])^(a[13] & b[102])^(a[12] & b[103])^(a[11] & b[104])^(a[10] & b[105])^(a[9] & b[106])^(a[8] & b[107])^(a[7] & b[108])^(a[6] & b[109])^(a[5] & b[110])^(a[4] & b[111])^(a[3] & b[112])^(a[2] & b[113])^(a[1] & b[114])^(a[0] & b[115]);
assign y[116] = (a[116] & b[0])^(a[115] & b[1])^(a[114] & b[2])^(a[113] & b[3])^(a[112] & b[4])^(a[111] & b[5])^(a[110] & b[6])^(a[109] & b[7])^(a[108] & b[8])^(a[107] & b[9])^(a[106] & b[10])^(a[105] & b[11])^(a[104] & b[12])^(a[103] & b[13])^(a[102] & b[14])^(a[101] & b[15])^(a[100] & b[16])^(a[99] & b[17])^(a[98] & b[18])^(a[97] & b[19])^(a[96] & b[20])^(a[95] & b[21])^(a[94] & b[22])^(a[93] & b[23])^(a[92] & b[24])^(a[91] & b[25])^(a[90] & b[26])^(a[89] & b[27])^(a[88] & b[28])^(a[87] & b[29])^(a[86] & b[30])^(a[85] & b[31])^(a[84] & b[32])^(a[83] & b[33])^(a[82] & b[34])^(a[81] & b[35])^(a[80] & b[36])^(a[79] & b[37])^(a[78] & b[38])^(a[77] & b[39])^(a[76] & b[40])^(a[75] & b[41])^(a[74] & b[42])^(a[73] & b[43])^(a[72] & b[44])^(a[71] & b[45])^(a[70] & b[46])^(a[69] & b[47])^(a[68] & b[48])^(a[67] & b[49])^(a[66] & b[50])^(a[65] & b[51])^(a[64] & b[52])^(a[63] & b[53])^(a[62] & b[54])^(a[61] & b[55])^(a[60] & b[56])^(a[59] & b[57])^(a[58] & b[58])^(a[57] & b[59])^(a[56] & b[60])^(a[55] & b[61])^(a[54] & b[62])^(a[53] & b[63])^(a[52] & b[64])^(a[51] & b[65])^(a[50] & b[66])^(a[49] & b[67])^(a[48] & b[68])^(a[47] & b[69])^(a[46] & b[70])^(a[45] & b[71])^(a[44] & b[72])^(a[43] & b[73])^(a[42] & b[74])^(a[41] & b[75])^(a[40] & b[76])^(a[39] & b[77])^(a[38] & b[78])^(a[37] & b[79])^(a[36] & b[80])^(a[35] & b[81])^(a[34] & b[82])^(a[33] & b[83])^(a[32] & b[84])^(a[31] & b[85])^(a[30] & b[86])^(a[29] & b[87])^(a[28] & b[88])^(a[27] & b[89])^(a[26] & b[90])^(a[25] & b[91])^(a[24] & b[92])^(a[23] & b[93])^(a[22] & b[94])^(a[21] & b[95])^(a[20] & b[96])^(a[19] & b[97])^(a[18] & b[98])^(a[17] & b[99])^(a[16] & b[100])^(a[15] & b[101])^(a[14] & b[102])^(a[13] & b[103])^(a[12] & b[104])^(a[11] & b[105])^(a[10] & b[106])^(a[9] & b[107])^(a[8] & b[108])^(a[7] & b[109])^(a[6] & b[110])^(a[5] & b[111])^(a[4] & b[112])^(a[3] & b[113])^(a[2] & b[114])^(a[1] & b[115])^(a[0] & b[116]);
assign y[117] = (a[117] & b[0])^(a[116] & b[1])^(a[115] & b[2])^(a[114] & b[3])^(a[113] & b[4])^(a[112] & b[5])^(a[111] & b[6])^(a[110] & b[7])^(a[109] & b[8])^(a[108] & b[9])^(a[107] & b[10])^(a[106] & b[11])^(a[105] & b[12])^(a[104] & b[13])^(a[103] & b[14])^(a[102] & b[15])^(a[101] & b[16])^(a[100] & b[17])^(a[99] & b[18])^(a[98] & b[19])^(a[97] & b[20])^(a[96] & b[21])^(a[95] & b[22])^(a[94] & b[23])^(a[93] & b[24])^(a[92] & b[25])^(a[91] & b[26])^(a[90] & b[27])^(a[89] & b[28])^(a[88] & b[29])^(a[87] & b[30])^(a[86] & b[31])^(a[85] & b[32])^(a[84] & b[33])^(a[83] & b[34])^(a[82] & b[35])^(a[81] & b[36])^(a[80] & b[37])^(a[79] & b[38])^(a[78] & b[39])^(a[77] & b[40])^(a[76] & b[41])^(a[75] & b[42])^(a[74] & b[43])^(a[73] & b[44])^(a[72] & b[45])^(a[71] & b[46])^(a[70] & b[47])^(a[69] & b[48])^(a[68] & b[49])^(a[67] & b[50])^(a[66] & b[51])^(a[65] & b[52])^(a[64] & b[53])^(a[63] & b[54])^(a[62] & b[55])^(a[61] & b[56])^(a[60] & b[57])^(a[59] & b[58])^(a[58] & b[59])^(a[57] & b[60])^(a[56] & b[61])^(a[55] & b[62])^(a[54] & b[63])^(a[53] & b[64])^(a[52] & b[65])^(a[51] & b[66])^(a[50] & b[67])^(a[49] & b[68])^(a[48] & b[69])^(a[47] & b[70])^(a[46] & b[71])^(a[45] & b[72])^(a[44] & b[73])^(a[43] & b[74])^(a[42] & b[75])^(a[41] & b[76])^(a[40] & b[77])^(a[39] & b[78])^(a[38] & b[79])^(a[37] & b[80])^(a[36] & b[81])^(a[35] & b[82])^(a[34] & b[83])^(a[33] & b[84])^(a[32] & b[85])^(a[31] & b[86])^(a[30] & b[87])^(a[29] & b[88])^(a[28] & b[89])^(a[27] & b[90])^(a[26] & b[91])^(a[25] & b[92])^(a[24] & b[93])^(a[23] & b[94])^(a[22] & b[95])^(a[21] & b[96])^(a[20] & b[97])^(a[19] & b[98])^(a[18] & b[99])^(a[17] & b[100])^(a[16] & b[101])^(a[15] & b[102])^(a[14] & b[103])^(a[13] & b[104])^(a[12] & b[105])^(a[11] & b[106])^(a[10] & b[107])^(a[9] & b[108])^(a[8] & b[109])^(a[7] & b[110])^(a[6] & b[111])^(a[5] & b[112])^(a[4] & b[113])^(a[3] & b[114])^(a[2] & b[115])^(a[1] & b[116])^(a[0] & b[117]);
assign y[118] = (a[118] & b[0])^(a[117] & b[1])^(a[116] & b[2])^(a[115] & b[3])^(a[114] & b[4])^(a[113] & b[5])^(a[112] & b[6])^(a[111] & b[7])^(a[110] & b[8])^(a[109] & b[9])^(a[108] & b[10])^(a[107] & b[11])^(a[106] & b[12])^(a[105] & b[13])^(a[104] & b[14])^(a[103] & b[15])^(a[102] & b[16])^(a[101] & b[17])^(a[100] & b[18])^(a[99] & b[19])^(a[98] & b[20])^(a[97] & b[21])^(a[96] & b[22])^(a[95] & b[23])^(a[94] & b[24])^(a[93] & b[25])^(a[92] & b[26])^(a[91] & b[27])^(a[90] & b[28])^(a[89] & b[29])^(a[88] & b[30])^(a[87] & b[31])^(a[86] & b[32])^(a[85] & b[33])^(a[84] & b[34])^(a[83] & b[35])^(a[82] & b[36])^(a[81] & b[37])^(a[80] & b[38])^(a[79] & b[39])^(a[78] & b[40])^(a[77] & b[41])^(a[76] & b[42])^(a[75] & b[43])^(a[74] & b[44])^(a[73] & b[45])^(a[72] & b[46])^(a[71] & b[47])^(a[70] & b[48])^(a[69] & b[49])^(a[68] & b[50])^(a[67] & b[51])^(a[66] & b[52])^(a[65] & b[53])^(a[64] & b[54])^(a[63] & b[55])^(a[62] & b[56])^(a[61] & b[57])^(a[60] & b[58])^(a[59] & b[59])^(a[58] & b[60])^(a[57] & b[61])^(a[56] & b[62])^(a[55] & b[63])^(a[54] & b[64])^(a[53] & b[65])^(a[52] & b[66])^(a[51] & b[67])^(a[50] & b[68])^(a[49] & b[69])^(a[48] & b[70])^(a[47] & b[71])^(a[46] & b[72])^(a[45] & b[73])^(a[44] & b[74])^(a[43] & b[75])^(a[42] & b[76])^(a[41] & b[77])^(a[40] & b[78])^(a[39] & b[79])^(a[38] & b[80])^(a[37] & b[81])^(a[36] & b[82])^(a[35] & b[83])^(a[34] & b[84])^(a[33] & b[85])^(a[32] & b[86])^(a[31] & b[87])^(a[30] & b[88])^(a[29] & b[89])^(a[28] & b[90])^(a[27] & b[91])^(a[26] & b[92])^(a[25] & b[93])^(a[24] & b[94])^(a[23] & b[95])^(a[22] & b[96])^(a[21] & b[97])^(a[20] & b[98])^(a[19] & b[99])^(a[18] & b[100])^(a[17] & b[101])^(a[16] & b[102])^(a[15] & b[103])^(a[14] & b[104])^(a[13] & b[105])^(a[12] & b[106])^(a[11] & b[107])^(a[10] & b[108])^(a[9] & b[109])^(a[8] & b[110])^(a[7] & b[111])^(a[6] & b[112])^(a[5] & b[113])^(a[4] & b[114])^(a[3] & b[115])^(a[2] & b[116])^(a[1] & b[117])^(a[0] & b[118]);
assign y[119] = (a[119] & b[0])^(a[118] & b[1])^(a[117] & b[2])^(a[116] & b[3])^(a[115] & b[4])^(a[114] & b[5])^(a[113] & b[6])^(a[112] & b[7])^(a[111] & b[8])^(a[110] & b[9])^(a[109] & b[10])^(a[108] & b[11])^(a[107] & b[12])^(a[106] & b[13])^(a[105] & b[14])^(a[104] & b[15])^(a[103] & b[16])^(a[102] & b[17])^(a[101] & b[18])^(a[100] & b[19])^(a[99] & b[20])^(a[98] & b[21])^(a[97] & b[22])^(a[96] & b[23])^(a[95] & b[24])^(a[94] & b[25])^(a[93] & b[26])^(a[92] & b[27])^(a[91] & b[28])^(a[90] & b[29])^(a[89] & b[30])^(a[88] & b[31])^(a[87] & b[32])^(a[86] & b[33])^(a[85] & b[34])^(a[84] & b[35])^(a[83] & b[36])^(a[82] & b[37])^(a[81] & b[38])^(a[80] & b[39])^(a[79] & b[40])^(a[78] & b[41])^(a[77] & b[42])^(a[76] & b[43])^(a[75] & b[44])^(a[74] & b[45])^(a[73] & b[46])^(a[72] & b[47])^(a[71] & b[48])^(a[70] & b[49])^(a[69] & b[50])^(a[68] & b[51])^(a[67] & b[52])^(a[66] & b[53])^(a[65] & b[54])^(a[64] & b[55])^(a[63] & b[56])^(a[62] & b[57])^(a[61] & b[58])^(a[60] & b[59])^(a[59] & b[60])^(a[58] & b[61])^(a[57] & b[62])^(a[56] & b[63])^(a[55] & b[64])^(a[54] & b[65])^(a[53] & b[66])^(a[52] & b[67])^(a[51] & b[68])^(a[50] & b[69])^(a[49] & b[70])^(a[48] & b[71])^(a[47] & b[72])^(a[46] & b[73])^(a[45] & b[74])^(a[44] & b[75])^(a[43] & b[76])^(a[42] & b[77])^(a[41] & b[78])^(a[40] & b[79])^(a[39] & b[80])^(a[38] & b[81])^(a[37] & b[82])^(a[36] & b[83])^(a[35] & b[84])^(a[34] & b[85])^(a[33] & b[86])^(a[32] & b[87])^(a[31] & b[88])^(a[30] & b[89])^(a[29] & b[90])^(a[28] & b[91])^(a[27] & b[92])^(a[26] & b[93])^(a[25] & b[94])^(a[24] & b[95])^(a[23] & b[96])^(a[22] & b[97])^(a[21] & b[98])^(a[20] & b[99])^(a[19] & b[100])^(a[18] & b[101])^(a[17] & b[102])^(a[16] & b[103])^(a[15] & b[104])^(a[14] & b[105])^(a[13] & b[106])^(a[12] & b[107])^(a[11] & b[108])^(a[10] & b[109])^(a[9] & b[110])^(a[8] & b[111])^(a[7] & b[112])^(a[6] & b[113])^(a[5] & b[114])^(a[4] & b[115])^(a[3] & b[116])^(a[2] & b[117])^(a[1] & b[118])^(a[0] & b[119]);
assign y[120] = (a[120] & b[0])^(a[119] & b[1])^(a[118] & b[2])^(a[117] & b[3])^(a[116] & b[4])^(a[115] & b[5])^(a[114] & b[6])^(a[113] & b[7])^(a[112] & b[8])^(a[111] & b[9])^(a[110] & b[10])^(a[109] & b[11])^(a[108] & b[12])^(a[107] & b[13])^(a[106] & b[14])^(a[105] & b[15])^(a[104] & b[16])^(a[103] & b[17])^(a[102] & b[18])^(a[101] & b[19])^(a[100] & b[20])^(a[99] & b[21])^(a[98] & b[22])^(a[97] & b[23])^(a[96] & b[24])^(a[95] & b[25])^(a[94] & b[26])^(a[93] & b[27])^(a[92] & b[28])^(a[91] & b[29])^(a[90] & b[30])^(a[89] & b[31])^(a[88] & b[32])^(a[87] & b[33])^(a[86] & b[34])^(a[85] & b[35])^(a[84] & b[36])^(a[83] & b[37])^(a[82] & b[38])^(a[81] & b[39])^(a[80] & b[40])^(a[79] & b[41])^(a[78] & b[42])^(a[77] & b[43])^(a[76] & b[44])^(a[75] & b[45])^(a[74] & b[46])^(a[73] & b[47])^(a[72] & b[48])^(a[71] & b[49])^(a[70] & b[50])^(a[69] & b[51])^(a[68] & b[52])^(a[67] & b[53])^(a[66] & b[54])^(a[65] & b[55])^(a[64] & b[56])^(a[63] & b[57])^(a[62] & b[58])^(a[61] & b[59])^(a[60] & b[60])^(a[59] & b[61])^(a[58] & b[62])^(a[57] & b[63])^(a[56] & b[64])^(a[55] & b[65])^(a[54] & b[66])^(a[53] & b[67])^(a[52] & b[68])^(a[51] & b[69])^(a[50] & b[70])^(a[49] & b[71])^(a[48] & b[72])^(a[47] & b[73])^(a[46] & b[74])^(a[45] & b[75])^(a[44] & b[76])^(a[43] & b[77])^(a[42] & b[78])^(a[41] & b[79])^(a[40] & b[80])^(a[39] & b[81])^(a[38] & b[82])^(a[37] & b[83])^(a[36] & b[84])^(a[35] & b[85])^(a[34] & b[86])^(a[33] & b[87])^(a[32] & b[88])^(a[31] & b[89])^(a[30] & b[90])^(a[29] & b[91])^(a[28] & b[92])^(a[27] & b[93])^(a[26] & b[94])^(a[25] & b[95])^(a[24] & b[96])^(a[23] & b[97])^(a[22] & b[98])^(a[21] & b[99])^(a[20] & b[100])^(a[19] & b[101])^(a[18] & b[102])^(a[17] & b[103])^(a[16] & b[104])^(a[15] & b[105])^(a[14] & b[106])^(a[13] & b[107])^(a[12] & b[108])^(a[11] & b[109])^(a[10] & b[110])^(a[9] & b[111])^(a[8] & b[112])^(a[7] & b[113])^(a[6] & b[114])^(a[5] & b[115])^(a[4] & b[116])^(a[3] & b[117])^(a[2] & b[118])^(a[1] & b[119])^(a[0] & b[120]);
assign y[121] = (a[121] & b[0])^(a[120] & b[1])^(a[119] & b[2])^(a[118] & b[3])^(a[117] & b[4])^(a[116] & b[5])^(a[115] & b[6])^(a[114] & b[7])^(a[113] & b[8])^(a[112] & b[9])^(a[111] & b[10])^(a[110] & b[11])^(a[109] & b[12])^(a[108] & b[13])^(a[107] & b[14])^(a[106] & b[15])^(a[105] & b[16])^(a[104] & b[17])^(a[103] & b[18])^(a[102] & b[19])^(a[101] & b[20])^(a[100] & b[21])^(a[99] & b[22])^(a[98] & b[23])^(a[97] & b[24])^(a[96] & b[25])^(a[95] & b[26])^(a[94] & b[27])^(a[93] & b[28])^(a[92] & b[29])^(a[91] & b[30])^(a[90] & b[31])^(a[89] & b[32])^(a[88] & b[33])^(a[87] & b[34])^(a[86] & b[35])^(a[85] & b[36])^(a[84] & b[37])^(a[83] & b[38])^(a[82] & b[39])^(a[81] & b[40])^(a[80] & b[41])^(a[79] & b[42])^(a[78] & b[43])^(a[77] & b[44])^(a[76] & b[45])^(a[75] & b[46])^(a[74] & b[47])^(a[73] & b[48])^(a[72] & b[49])^(a[71] & b[50])^(a[70] & b[51])^(a[69] & b[52])^(a[68] & b[53])^(a[67] & b[54])^(a[66] & b[55])^(a[65] & b[56])^(a[64] & b[57])^(a[63] & b[58])^(a[62] & b[59])^(a[61] & b[60])^(a[60] & b[61])^(a[59] & b[62])^(a[58] & b[63])^(a[57] & b[64])^(a[56] & b[65])^(a[55] & b[66])^(a[54] & b[67])^(a[53] & b[68])^(a[52] & b[69])^(a[51] & b[70])^(a[50] & b[71])^(a[49] & b[72])^(a[48] & b[73])^(a[47] & b[74])^(a[46] & b[75])^(a[45] & b[76])^(a[44] & b[77])^(a[43] & b[78])^(a[42] & b[79])^(a[41] & b[80])^(a[40] & b[81])^(a[39] & b[82])^(a[38] & b[83])^(a[37] & b[84])^(a[36] & b[85])^(a[35] & b[86])^(a[34] & b[87])^(a[33] & b[88])^(a[32] & b[89])^(a[31] & b[90])^(a[30] & b[91])^(a[29] & b[92])^(a[28] & b[93])^(a[27] & b[94])^(a[26] & b[95])^(a[25] & b[96])^(a[24] & b[97])^(a[23] & b[98])^(a[22] & b[99])^(a[21] & b[100])^(a[20] & b[101])^(a[19] & b[102])^(a[18] & b[103])^(a[17] & b[104])^(a[16] & b[105])^(a[15] & b[106])^(a[14] & b[107])^(a[13] & b[108])^(a[12] & b[109])^(a[11] & b[110])^(a[10] & b[111])^(a[9] & b[112])^(a[8] & b[113])^(a[7] & b[114])^(a[6] & b[115])^(a[5] & b[116])^(a[4] & b[117])^(a[3] & b[118])^(a[2] & b[119])^(a[1] & b[120])^(a[0] & b[121]);
assign y[122] = (a[122] & b[0])^(a[121] & b[1])^(a[120] & b[2])^(a[119] & b[3])^(a[118] & b[4])^(a[117] & b[5])^(a[116] & b[6])^(a[115] & b[7])^(a[114] & b[8])^(a[113] & b[9])^(a[112] & b[10])^(a[111] & b[11])^(a[110] & b[12])^(a[109] & b[13])^(a[108] & b[14])^(a[107] & b[15])^(a[106] & b[16])^(a[105] & b[17])^(a[104] & b[18])^(a[103] & b[19])^(a[102] & b[20])^(a[101] & b[21])^(a[100] & b[22])^(a[99] & b[23])^(a[98] & b[24])^(a[97] & b[25])^(a[96] & b[26])^(a[95] & b[27])^(a[94] & b[28])^(a[93] & b[29])^(a[92] & b[30])^(a[91] & b[31])^(a[90] & b[32])^(a[89] & b[33])^(a[88] & b[34])^(a[87] & b[35])^(a[86] & b[36])^(a[85] & b[37])^(a[84] & b[38])^(a[83] & b[39])^(a[82] & b[40])^(a[81] & b[41])^(a[80] & b[42])^(a[79] & b[43])^(a[78] & b[44])^(a[77] & b[45])^(a[76] & b[46])^(a[75] & b[47])^(a[74] & b[48])^(a[73] & b[49])^(a[72] & b[50])^(a[71] & b[51])^(a[70] & b[52])^(a[69] & b[53])^(a[68] & b[54])^(a[67] & b[55])^(a[66] & b[56])^(a[65] & b[57])^(a[64] & b[58])^(a[63] & b[59])^(a[62] & b[60])^(a[61] & b[61])^(a[60] & b[62])^(a[59] & b[63])^(a[58] & b[64])^(a[57] & b[65])^(a[56] & b[66])^(a[55] & b[67])^(a[54] & b[68])^(a[53] & b[69])^(a[52] & b[70])^(a[51] & b[71])^(a[50] & b[72])^(a[49] & b[73])^(a[48] & b[74])^(a[47] & b[75])^(a[46] & b[76])^(a[45] & b[77])^(a[44] & b[78])^(a[43] & b[79])^(a[42] & b[80])^(a[41] & b[81])^(a[40] & b[82])^(a[39] & b[83])^(a[38] & b[84])^(a[37] & b[85])^(a[36] & b[86])^(a[35] & b[87])^(a[34] & b[88])^(a[33] & b[89])^(a[32] & b[90])^(a[31] & b[91])^(a[30] & b[92])^(a[29] & b[93])^(a[28] & b[94])^(a[27] & b[95])^(a[26] & b[96])^(a[25] & b[97])^(a[24] & b[98])^(a[23] & b[99])^(a[22] & b[100])^(a[21] & b[101])^(a[20] & b[102])^(a[19] & b[103])^(a[18] & b[104])^(a[17] & b[105])^(a[16] & b[106])^(a[15] & b[107])^(a[14] & b[108])^(a[13] & b[109])^(a[12] & b[110])^(a[11] & b[111])^(a[10] & b[112])^(a[9] & b[113])^(a[8] & b[114])^(a[7] & b[115])^(a[6] & b[116])^(a[5] & b[117])^(a[4] & b[118])^(a[3] & b[119])^(a[2] & b[120])^(a[1] & b[121])^(a[0] & b[122]);
assign y[123] = (a[123] & b[0])^(a[122] & b[1])^(a[121] & b[2])^(a[120] & b[3])^(a[119] & b[4])^(a[118] & b[5])^(a[117] & b[6])^(a[116] & b[7])^(a[115] & b[8])^(a[114] & b[9])^(a[113] & b[10])^(a[112] & b[11])^(a[111] & b[12])^(a[110] & b[13])^(a[109] & b[14])^(a[108] & b[15])^(a[107] & b[16])^(a[106] & b[17])^(a[105] & b[18])^(a[104] & b[19])^(a[103] & b[20])^(a[102] & b[21])^(a[101] & b[22])^(a[100] & b[23])^(a[99] & b[24])^(a[98] & b[25])^(a[97] & b[26])^(a[96] & b[27])^(a[95] & b[28])^(a[94] & b[29])^(a[93] & b[30])^(a[92] & b[31])^(a[91] & b[32])^(a[90] & b[33])^(a[89] & b[34])^(a[88] & b[35])^(a[87] & b[36])^(a[86] & b[37])^(a[85] & b[38])^(a[84] & b[39])^(a[83] & b[40])^(a[82] & b[41])^(a[81] & b[42])^(a[80] & b[43])^(a[79] & b[44])^(a[78] & b[45])^(a[77] & b[46])^(a[76] & b[47])^(a[75] & b[48])^(a[74] & b[49])^(a[73] & b[50])^(a[72] & b[51])^(a[71] & b[52])^(a[70] & b[53])^(a[69] & b[54])^(a[68] & b[55])^(a[67] & b[56])^(a[66] & b[57])^(a[65] & b[58])^(a[64] & b[59])^(a[63] & b[60])^(a[62] & b[61])^(a[61] & b[62])^(a[60] & b[63])^(a[59] & b[64])^(a[58] & b[65])^(a[57] & b[66])^(a[56] & b[67])^(a[55] & b[68])^(a[54] & b[69])^(a[53] & b[70])^(a[52] & b[71])^(a[51] & b[72])^(a[50] & b[73])^(a[49] & b[74])^(a[48] & b[75])^(a[47] & b[76])^(a[46] & b[77])^(a[45] & b[78])^(a[44] & b[79])^(a[43] & b[80])^(a[42] & b[81])^(a[41] & b[82])^(a[40] & b[83])^(a[39] & b[84])^(a[38] & b[85])^(a[37] & b[86])^(a[36] & b[87])^(a[35] & b[88])^(a[34] & b[89])^(a[33] & b[90])^(a[32] & b[91])^(a[31] & b[92])^(a[30] & b[93])^(a[29] & b[94])^(a[28] & b[95])^(a[27] & b[96])^(a[26] & b[97])^(a[25] & b[98])^(a[24] & b[99])^(a[23] & b[100])^(a[22] & b[101])^(a[21] & b[102])^(a[20] & b[103])^(a[19] & b[104])^(a[18] & b[105])^(a[17] & b[106])^(a[16] & b[107])^(a[15] & b[108])^(a[14] & b[109])^(a[13] & b[110])^(a[12] & b[111])^(a[11] & b[112])^(a[10] & b[113])^(a[9] & b[114])^(a[8] & b[115])^(a[7] & b[116])^(a[6] & b[117])^(a[5] & b[118])^(a[4] & b[119])^(a[3] & b[120])^(a[2] & b[121])^(a[1] & b[122])^(a[0] & b[123]);
assign y[124] = (a[124] & b[0])^(a[123] & b[1])^(a[122] & b[2])^(a[121] & b[3])^(a[120] & b[4])^(a[119] & b[5])^(a[118] & b[6])^(a[117] & b[7])^(a[116] & b[8])^(a[115] & b[9])^(a[114] & b[10])^(a[113] & b[11])^(a[112] & b[12])^(a[111] & b[13])^(a[110] & b[14])^(a[109] & b[15])^(a[108] & b[16])^(a[107] & b[17])^(a[106] & b[18])^(a[105] & b[19])^(a[104] & b[20])^(a[103] & b[21])^(a[102] & b[22])^(a[101] & b[23])^(a[100] & b[24])^(a[99] & b[25])^(a[98] & b[26])^(a[97] & b[27])^(a[96] & b[28])^(a[95] & b[29])^(a[94] & b[30])^(a[93] & b[31])^(a[92] & b[32])^(a[91] & b[33])^(a[90] & b[34])^(a[89] & b[35])^(a[88] & b[36])^(a[87] & b[37])^(a[86] & b[38])^(a[85] & b[39])^(a[84] & b[40])^(a[83] & b[41])^(a[82] & b[42])^(a[81] & b[43])^(a[80] & b[44])^(a[79] & b[45])^(a[78] & b[46])^(a[77] & b[47])^(a[76] & b[48])^(a[75] & b[49])^(a[74] & b[50])^(a[73] & b[51])^(a[72] & b[52])^(a[71] & b[53])^(a[70] & b[54])^(a[69] & b[55])^(a[68] & b[56])^(a[67] & b[57])^(a[66] & b[58])^(a[65] & b[59])^(a[64] & b[60])^(a[63] & b[61])^(a[62] & b[62])^(a[61] & b[63])^(a[60] & b[64])^(a[59] & b[65])^(a[58] & b[66])^(a[57] & b[67])^(a[56] & b[68])^(a[55] & b[69])^(a[54] & b[70])^(a[53] & b[71])^(a[52] & b[72])^(a[51] & b[73])^(a[50] & b[74])^(a[49] & b[75])^(a[48] & b[76])^(a[47] & b[77])^(a[46] & b[78])^(a[45] & b[79])^(a[44] & b[80])^(a[43] & b[81])^(a[42] & b[82])^(a[41] & b[83])^(a[40] & b[84])^(a[39] & b[85])^(a[38] & b[86])^(a[37] & b[87])^(a[36] & b[88])^(a[35] & b[89])^(a[34] & b[90])^(a[33] & b[91])^(a[32] & b[92])^(a[31] & b[93])^(a[30] & b[94])^(a[29] & b[95])^(a[28] & b[96])^(a[27] & b[97])^(a[26] & b[98])^(a[25] & b[99])^(a[24] & b[100])^(a[23] & b[101])^(a[22] & b[102])^(a[21] & b[103])^(a[20] & b[104])^(a[19] & b[105])^(a[18] & b[106])^(a[17] & b[107])^(a[16] & b[108])^(a[15] & b[109])^(a[14] & b[110])^(a[13] & b[111])^(a[12] & b[112])^(a[11] & b[113])^(a[10] & b[114])^(a[9] & b[115])^(a[8] & b[116])^(a[7] & b[117])^(a[6] & b[118])^(a[5] & b[119])^(a[4] & b[120])^(a[3] & b[121])^(a[2] & b[122])^(a[1] & b[123])^(a[0] & b[124]);
assign y[125] = (a[125] & b[0])^(a[124] & b[1])^(a[123] & b[2])^(a[122] & b[3])^(a[121] & b[4])^(a[120] & b[5])^(a[119] & b[6])^(a[118] & b[7])^(a[117] & b[8])^(a[116] & b[9])^(a[115] & b[10])^(a[114] & b[11])^(a[113] & b[12])^(a[112] & b[13])^(a[111] & b[14])^(a[110] & b[15])^(a[109] & b[16])^(a[108] & b[17])^(a[107] & b[18])^(a[106] & b[19])^(a[105] & b[20])^(a[104] & b[21])^(a[103] & b[22])^(a[102] & b[23])^(a[101] & b[24])^(a[100] & b[25])^(a[99] & b[26])^(a[98] & b[27])^(a[97] & b[28])^(a[96] & b[29])^(a[95] & b[30])^(a[94] & b[31])^(a[93] & b[32])^(a[92] & b[33])^(a[91] & b[34])^(a[90] & b[35])^(a[89] & b[36])^(a[88] & b[37])^(a[87] & b[38])^(a[86] & b[39])^(a[85] & b[40])^(a[84] & b[41])^(a[83] & b[42])^(a[82] & b[43])^(a[81] & b[44])^(a[80] & b[45])^(a[79] & b[46])^(a[78] & b[47])^(a[77] & b[48])^(a[76] & b[49])^(a[75] & b[50])^(a[74] & b[51])^(a[73] & b[52])^(a[72] & b[53])^(a[71] & b[54])^(a[70] & b[55])^(a[69] & b[56])^(a[68] & b[57])^(a[67] & b[58])^(a[66] & b[59])^(a[65] & b[60])^(a[64] & b[61])^(a[63] & b[62])^(a[62] & b[63])^(a[61] & b[64])^(a[60] & b[65])^(a[59] & b[66])^(a[58] & b[67])^(a[57] & b[68])^(a[56] & b[69])^(a[55] & b[70])^(a[54] & b[71])^(a[53] & b[72])^(a[52] & b[73])^(a[51] & b[74])^(a[50] & b[75])^(a[49] & b[76])^(a[48] & b[77])^(a[47] & b[78])^(a[46] & b[79])^(a[45] & b[80])^(a[44] & b[81])^(a[43] & b[82])^(a[42] & b[83])^(a[41] & b[84])^(a[40] & b[85])^(a[39] & b[86])^(a[38] & b[87])^(a[37] & b[88])^(a[36] & b[89])^(a[35] & b[90])^(a[34] & b[91])^(a[33] & b[92])^(a[32] & b[93])^(a[31] & b[94])^(a[30] & b[95])^(a[29] & b[96])^(a[28] & b[97])^(a[27] & b[98])^(a[26] & b[99])^(a[25] & b[100])^(a[24] & b[101])^(a[23] & b[102])^(a[22] & b[103])^(a[21] & b[104])^(a[20] & b[105])^(a[19] & b[106])^(a[18] & b[107])^(a[17] & b[108])^(a[16] & b[109])^(a[15] & b[110])^(a[14] & b[111])^(a[13] & b[112])^(a[12] & b[113])^(a[11] & b[114])^(a[10] & b[115])^(a[9] & b[116])^(a[8] & b[117])^(a[7] & b[118])^(a[6] & b[119])^(a[5] & b[120])^(a[4] & b[121])^(a[3] & b[122])^(a[2] & b[123])^(a[1] & b[124])^(a[0] & b[125]);
assign y[126] = (a[126] & b[0])^(a[125] & b[1])^(a[124] & b[2])^(a[123] & b[3])^(a[122] & b[4])^(a[121] & b[5])^(a[120] & b[6])^(a[119] & b[7])^(a[118] & b[8])^(a[117] & b[9])^(a[116] & b[10])^(a[115] & b[11])^(a[114] & b[12])^(a[113] & b[13])^(a[112] & b[14])^(a[111] & b[15])^(a[110] & b[16])^(a[109] & b[17])^(a[108] & b[18])^(a[107] & b[19])^(a[106] & b[20])^(a[105] & b[21])^(a[104] & b[22])^(a[103] & b[23])^(a[102] & b[24])^(a[101] & b[25])^(a[100] & b[26])^(a[99] & b[27])^(a[98] & b[28])^(a[97] & b[29])^(a[96] & b[30])^(a[95] & b[31])^(a[94] & b[32])^(a[93] & b[33])^(a[92] & b[34])^(a[91] & b[35])^(a[90] & b[36])^(a[89] & b[37])^(a[88] & b[38])^(a[87] & b[39])^(a[86] & b[40])^(a[85] & b[41])^(a[84] & b[42])^(a[83] & b[43])^(a[82] & b[44])^(a[81] & b[45])^(a[80] & b[46])^(a[79] & b[47])^(a[78] & b[48])^(a[77] & b[49])^(a[76] & b[50])^(a[75] & b[51])^(a[74] & b[52])^(a[73] & b[53])^(a[72] & b[54])^(a[71] & b[55])^(a[70] & b[56])^(a[69] & b[57])^(a[68] & b[58])^(a[67] & b[59])^(a[66] & b[60])^(a[65] & b[61])^(a[64] & b[62])^(a[63] & b[63])^(a[62] & b[64])^(a[61] & b[65])^(a[60] & b[66])^(a[59] & b[67])^(a[58] & b[68])^(a[57] & b[69])^(a[56] & b[70])^(a[55] & b[71])^(a[54] & b[72])^(a[53] & b[73])^(a[52] & b[74])^(a[51] & b[75])^(a[50] & b[76])^(a[49] & b[77])^(a[48] & b[78])^(a[47] & b[79])^(a[46] & b[80])^(a[45] & b[81])^(a[44] & b[82])^(a[43] & b[83])^(a[42] & b[84])^(a[41] & b[85])^(a[40] & b[86])^(a[39] & b[87])^(a[38] & b[88])^(a[37] & b[89])^(a[36] & b[90])^(a[35] & b[91])^(a[34] & b[92])^(a[33] & b[93])^(a[32] & b[94])^(a[31] & b[95])^(a[30] & b[96])^(a[29] & b[97])^(a[28] & b[98])^(a[27] & b[99])^(a[26] & b[100])^(a[25] & b[101])^(a[24] & b[102])^(a[23] & b[103])^(a[22] & b[104])^(a[21] & b[105])^(a[20] & b[106])^(a[19] & b[107])^(a[18] & b[108])^(a[17] & b[109])^(a[16] & b[110])^(a[15] & b[111])^(a[14] & b[112])^(a[13] & b[113])^(a[12] & b[114])^(a[11] & b[115])^(a[10] & b[116])^(a[9] & b[117])^(a[8] & b[118])^(a[7] & b[119])^(a[6] & b[120])^(a[5] & b[121])^(a[4] & b[122])^(a[3] & b[123])^(a[2] & b[124])^(a[1] & b[125])^(a[0] & b[126]);
assign y[127] = (a[127] & b[0])^(a[126] & b[1])^(a[125] & b[2])^(a[124] & b[3])^(a[123] & b[4])^(a[122] & b[5])^(a[121] & b[6])^(a[120] & b[7])^(a[119] & b[8])^(a[118] & b[9])^(a[117] & b[10])^(a[116] & b[11])^(a[115] & b[12])^(a[114] & b[13])^(a[113] & b[14])^(a[112] & b[15])^(a[111] & b[16])^(a[110] & b[17])^(a[109] & b[18])^(a[108] & b[19])^(a[107] & b[20])^(a[106] & b[21])^(a[105] & b[22])^(a[104] & b[23])^(a[103] & b[24])^(a[102] & b[25])^(a[101] & b[26])^(a[100] & b[27])^(a[99] & b[28])^(a[98] & b[29])^(a[97] & b[30])^(a[96] & b[31])^(a[95] & b[32])^(a[94] & b[33])^(a[93] & b[34])^(a[92] & b[35])^(a[91] & b[36])^(a[90] & b[37])^(a[89] & b[38])^(a[88] & b[39])^(a[87] & b[40])^(a[86] & b[41])^(a[85] & b[42])^(a[84] & b[43])^(a[83] & b[44])^(a[82] & b[45])^(a[81] & b[46])^(a[80] & b[47])^(a[79] & b[48])^(a[78] & b[49])^(a[77] & b[50])^(a[76] & b[51])^(a[75] & b[52])^(a[74] & b[53])^(a[73] & b[54])^(a[72] & b[55])^(a[71] & b[56])^(a[70] & b[57])^(a[69] & b[58])^(a[68] & b[59])^(a[67] & b[60])^(a[66] & b[61])^(a[65] & b[62])^(a[64] & b[63])^(a[63] & b[64])^(a[62] & b[65])^(a[61] & b[66])^(a[60] & b[67])^(a[59] & b[68])^(a[58] & b[69])^(a[57] & b[70])^(a[56] & b[71])^(a[55] & b[72])^(a[54] & b[73])^(a[53] & b[74])^(a[52] & b[75])^(a[51] & b[76])^(a[50] & b[77])^(a[49] & b[78])^(a[48] & b[79])^(a[47] & b[80])^(a[46] & b[81])^(a[45] & b[82])^(a[44] & b[83])^(a[43] & b[84])^(a[42] & b[85])^(a[41] & b[86])^(a[40] & b[87])^(a[39] & b[88])^(a[38] & b[89])^(a[37] & b[90])^(a[36] & b[91])^(a[35] & b[92])^(a[34] & b[93])^(a[33] & b[94])^(a[32] & b[95])^(a[31] & b[96])^(a[30] & b[97])^(a[29] & b[98])^(a[28] & b[99])^(a[27] & b[100])^(a[26] & b[101])^(a[25] & b[102])^(a[24] & b[103])^(a[23] & b[104])^(a[22] & b[105])^(a[21] & b[106])^(a[20] & b[107])^(a[19] & b[108])^(a[18] & b[109])^(a[17] & b[110])^(a[16] & b[111])^(a[15] & b[112])^(a[14] & b[113])^(a[13] & b[114])^(a[12] & b[115])^(a[11] & b[116])^(a[10] & b[117])^(a[9] & b[118])^(a[8] & b[119])^(a[7] & b[120])^(a[6] & b[121])^(a[5] & b[122])^(a[4] & b[123])^(a[3] & b[124])^(a[2] & b[125])^(a[1] & b[126])^(a[0] & b[127]);
assign y[128] = (a[128] & b[0])^(a[127] & b[1])^(a[126] & b[2])^(a[125] & b[3])^(a[124] & b[4])^(a[123] & b[5])^(a[122] & b[6])^(a[121] & b[7])^(a[120] & b[8])^(a[119] & b[9])^(a[118] & b[10])^(a[117] & b[11])^(a[116] & b[12])^(a[115] & b[13])^(a[114] & b[14])^(a[113] & b[15])^(a[112] & b[16])^(a[111] & b[17])^(a[110] & b[18])^(a[109] & b[19])^(a[108] & b[20])^(a[107] & b[21])^(a[106] & b[22])^(a[105] & b[23])^(a[104] & b[24])^(a[103] & b[25])^(a[102] & b[26])^(a[101] & b[27])^(a[100] & b[28])^(a[99] & b[29])^(a[98] & b[30])^(a[97] & b[31])^(a[96] & b[32])^(a[95] & b[33])^(a[94] & b[34])^(a[93] & b[35])^(a[92] & b[36])^(a[91] & b[37])^(a[90] & b[38])^(a[89] & b[39])^(a[88] & b[40])^(a[87] & b[41])^(a[86] & b[42])^(a[85] & b[43])^(a[84] & b[44])^(a[83] & b[45])^(a[82] & b[46])^(a[81] & b[47])^(a[80] & b[48])^(a[79] & b[49])^(a[78] & b[50])^(a[77] & b[51])^(a[76] & b[52])^(a[75] & b[53])^(a[74] & b[54])^(a[73] & b[55])^(a[72] & b[56])^(a[71] & b[57])^(a[70] & b[58])^(a[69] & b[59])^(a[68] & b[60])^(a[67] & b[61])^(a[66] & b[62])^(a[65] & b[63])^(a[64] & b[64])^(a[63] & b[65])^(a[62] & b[66])^(a[61] & b[67])^(a[60] & b[68])^(a[59] & b[69])^(a[58] & b[70])^(a[57] & b[71])^(a[56] & b[72])^(a[55] & b[73])^(a[54] & b[74])^(a[53] & b[75])^(a[52] & b[76])^(a[51] & b[77])^(a[50] & b[78])^(a[49] & b[79])^(a[48] & b[80])^(a[47] & b[81])^(a[46] & b[82])^(a[45] & b[83])^(a[44] & b[84])^(a[43] & b[85])^(a[42] & b[86])^(a[41] & b[87])^(a[40] & b[88])^(a[39] & b[89])^(a[38] & b[90])^(a[37] & b[91])^(a[36] & b[92])^(a[35] & b[93])^(a[34] & b[94])^(a[33] & b[95])^(a[32] & b[96])^(a[31] & b[97])^(a[30] & b[98])^(a[29] & b[99])^(a[28] & b[100])^(a[27] & b[101])^(a[26] & b[102])^(a[25] & b[103])^(a[24] & b[104])^(a[23] & b[105])^(a[22] & b[106])^(a[21] & b[107])^(a[20] & b[108])^(a[19] & b[109])^(a[18] & b[110])^(a[17] & b[111])^(a[16] & b[112])^(a[15] & b[113])^(a[14] & b[114])^(a[13] & b[115])^(a[12] & b[116])^(a[11] & b[117])^(a[10] & b[118])^(a[9] & b[119])^(a[8] & b[120])^(a[7] & b[121])^(a[6] & b[122])^(a[5] & b[123])^(a[4] & b[124])^(a[3] & b[125])^(a[2] & b[126])^(a[1] & b[127])^(a[0] & b[128]);
assign y[129] = (a[129] & b[0])^(a[128] & b[1])^(a[127] & b[2])^(a[126] & b[3])^(a[125] & b[4])^(a[124] & b[5])^(a[123] & b[6])^(a[122] & b[7])^(a[121] & b[8])^(a[120] & b[9])^(a[119] & b[10])^(a[118] & b[11])^(a[117] & b[12])^(a[116] & b[13])^(a[115] & b[14])^(a[114] & b[15])^(a[113] & b[16])^(a[112] & b[17])^(a[111] & b[18])^(a[110] & b[19])^(a[109] & b[20])^(a[108] & b[21])^(a[107] & b[22])^(a[106] & b[23])^(a[105] & b[24])^(a[104] & b[25])^(a[103] & b[26])^(a[102] & b[27])^(a[101] & b[28])^(a[100] & b[29])^(a[99] & b[30])^(a[98] & b[31])^(a[97] & b[32])^(a[96] & b[33])^(a[95] & b[34])^(a[94] & b[35])^(a[93] & b[36])^(a[92] & b[37])^(a[91] & b[38])^(a[90] & b[39])^(a[89] & b[40])^(a[88] & b[41])^(a[87] & b[42])^(a[86] & b[43])^(a[85] & b[44])^(a[84] & b[45])^(a[83] & b[46])^(a[82] & b[47])^(a[81] & b[48])^(a[80] & b[49])^(a[79] & b[50])^(a[78] & b[51])^(a[77] & b[52])^(a[76] & b[53])^(a[75] & b[54])^(a[74] & b[55])^(a[73] & b[56])^(a[72] & b[57])^(a[71] & b[58])^(a[70] & b[59])^(a[69] & b[60])^(a[68] & b[61])^(a[67] & b[62])^(a[66] & b[63])^(a[65] & b[64])^(a[64] & b[65])^(a[63] & b[66])^(a[62] & b[67])^(a[61] & b[68])^(a[60] & b[69])^(a[59] & b[70])^(a[58] & b[71])^(a[57] & b[72])^(a[56] & b[73])^(a[55] & b[74])^(a[54] & b[75])^(a[53] & b[76])^(a[52] & b[77])^(a[51] & b[78])^(a[50] & b[79])^(a[49] & b[80])^(a[48] & b[81])^(a[47] & b[82])^(a[46] & b[83])^(a[45] & b[84])^(a[44] & b[85])^(a[43] & b[86])^(a[42] & b[87])^(a[41] & b[88])^(a[40] & b[89])^(a[39] & b[90])^(a[38] & b[91])^(a[37] & b[92])^(a[36] & b[93])^(a[35] & b[94])^(a[34] & b[95])^(a[33] & b[96])^(a[32] & b[97])^(a[31] & b[98])^(a[30] & b[99])^(a[29] & b[100])^(a[28] & b[101])^(a[27] & b[102])^(a[26] & b[103])^(a[25] & b[104])^(a[24] & b[105])^(a[23] & b[106])^(a[22] & b[107])^(a[21] & b[108])^(a[20] & b[109])^(a[19] & b[110])^(a[18] & b[111])^(a[17] & b[112])^(a[16] & b[113])^(a[15] & b[114])^(a[14] & b[115])^(a[13] & b[116])^(a[12] & b[117])^(a[11] & b[118])^(a[10] & b[119])^(a[9] & b[120])^(a[8] & b[121])^(a[7] & b[122])^(a[6] & b[123])^(a[5] & b[124])^(a[4] & b[125])^(a[3] & b[126])^(a[2] & b[127])^(a[1] & b[128])^(a[0] & b[129]);
assign y[130] = (a[130] & b[0])^(a[129] & b[1])^(a[128] & b[2])^(a[127] & b[3])^(a[126] & b[4])^(a[125] & b[5])^(a[124] & b[6])^(a[123] & b[7])^(a[122] & b[8])^(a[121] & b[9])^(a[120] & b[10])^(a[119] & b[11])^(a[118] & b[12])^(a[117] & b[13])^(a[116] & b[14])^(a[115] & b[15])^(a[114] & b[16])^(a[113] & b[17])^(a[112] & b[18])^(a[111] & b[19])^(a[110] & b[20])^(a[109] & b[21])^(a[108] & b[22])^(a[107] & b[23])^(a[106] & b[24])^(a[105] & b[25])^(a[104] & b[26])^(a[103] & b[27])^(a[102] & b[28])^(a[101] & b[29])^(a[100] & b[30])^(a[99] & b[31])^(a[98] & b[32])^(a[97] & b[33])^(a[96] & b[34])^(a[95] & b[35])^(a[94] & b[36])^(a[93] & b[37])^(a[92] & b[38])^(a[91] & b[39])^(a[90] & b[40])^(a[89] & b[41])^(a[88] & b[42])^(a[87] & b[43])^(a[86] & b[44])^(a[85] & b[45])^(a[84] & b[46])^(a[83] & b[47])^(a[82] & b[48])^(a[81] & b[49])^(a[80] & b[50])^(a[79] & b[51])^(a[78] & b[52])^(a[77] & b[53])^(a[76] & b[54])^(a[75] & b[55])^(a[74] & b[56])^(a[73] & b[57])^(a[72] & b[58])^(a[71] & b[59])^(a[70] & b[60])^(a[69] & b[61])^(a[68] & b[62])^(a[67] & b[63])^(a[66] & b[64])^(a[65] & b[65])^(a[64] & b[66])^(a[63] & b[67])^(a[62] & b[68])^(a[61] & b[69])^(a[60] & b[70])^(a[59] & b[71])^(a[58] & b[72])^(a[57] & b[73])^(a[56] & b[74])^(a[55] & b[75])^(a[54] & b[76])^(a[53] & b[77])^(a[52] & b[78])^(a[51] & b[79])^(a[50] & b[80])^(a[49] & b[81])^(a[48] & b[82])^(a[47] & b[83])^(a[46] & b[84])^(a[45] & b[85])^(a[44] & b[86])^(a[43] & b[87])^(a[42] & b[88])^(a[41] & b[89])^(a[40] & b[90])^(a[39] & b[91])^(a[38] & b[92])^(a[37] & b[93])^(a[36] & b[94])^(a[35] & b[95])^(a[34] & b[96])^(a[33] & b[97])^(a[32] & b[98])^(a[31] & b[99])^(a[30] & b[100])^(a[29] & b[101])^(a[28] & b[102])^(a[27] & b[103])^(a[26] & b[104])^(a[25] & b[105])^(a[24] & b[106])^(a[23] & b[107])^(a[22] & b[108])^(a[21] & b[109])^(a[20] & b[110])^(a[19] & b[111])^(a[18] & b[112])^(a[17] & b[113])^(a[16] & b[114])^(a[15] & b[115])^(a[14] & b[116])^(a[13] & b[117])^(a[12] & b[118])^(a[11] & b[119])^(a[10] & b[120])^(a[9] & b[121])^(a[8] & b[122])^(a[7] & b[123])^(a[6] & b[124])^(a[5] & b[125])^(a[4] & b[126])^(a[3] & b[127])^(a[2] & b[128])^(a[1] & b[129])^(a[0] & b[130]);
assign y[131] = (a[131] & b[0])^(a[130] & b[1])^(a[129] & b[2])^(a[128] & b[3])^(a[127] & b[4])^(a[126] & b[5])^(a[125] & b[6])^(a[124] & b[7])^(a[123] & b[8])^(a[122] & b[9])^(a[121] & b[10])^(a[120] & b[11])^(a[119] & b[12])^(a[118] & b[13])^(a[117] & b[14])^(a[116] & b[15])^(a[115] & b[16])^(a[114] & b[17])^(a[113] & b[18])^(a[112] & b[19])^(a[111] & b[20])^(a[110] & b[21])^(a[109] & b[22])^(a[108] & b[23])^(a[107] & b[24])^(a[106] & b[25])^(a[105] & b[26])^(a[104] & b[27])^(a[103] & b[28])^(a[102] & b[29])^(a[101] & b[30])^(a[100] & b[31])^(a[99] & b[32])^(a[98] & b[33])^(a[97] & b[34])^(a[96] & b[35])^(a[95] & b[36])^(a[94] & b[37])^(a[93] & b[38])^(a[92] & b[39])^(a[91] & b[40])^(a[90] & b[41])^(a[89] & b[42])^(a[88] & b[43])^(a[87] & b[44])^(a[86] & b[45])^(a[85] & b[46])^(a[84] & b[47])^(a[83] & b[48])^(a[82] & b[49])^(a[81] & b[50])^(a[80] & b[51])^(a[79] & b[52])^(a[78] & b[53])^(a[77] & b[54])^(a[76] & b[55])^(a[75] & b[56])^(a[74] & b[57])^(a[73] & b[58])^(a[72] & b[59])^(a[71] & b[60])^(a[70] & b[61])^(a[69] & b[62])^(a[68] & b[63])^(a[67] & b[64])^(a[66] & b[65])^(a[65] & b[66])^(a[64] & b[67])^(a[63] & b[68])^(a[62] & b[69])^(a[61] & b[70])^(a[60] & b[71])^(a[59] & b[72])^(a[58] & b[73])^(a[57] & b[74])^(a[56] & b[75])^(a[55] & b[76])^(a[54] & b[77])^(a[53] & b[78])^(a[52] & b[79])^(a[51] & b[80])^(a[50] & b[81])^(a[49] & b[82])^(a[48] & b[83])^(a[47] & b[84])^(a[46] & b[85])^(a[45] & b[86])^(a[44] & b[87])^(a[43] & b[88])^(a[42] & b[89])^(a[41] & b[90])^(a[40] & b[91])^(a[39] & b[92])^(a[38] & b[93])^(a[37] & b[94])^(a[36] & b[95])^(a[35] & b[96])^(a[34] & b[97])^(a[33] & b[98])^(a[32] & b[99])^(a[31] & b[100])^(a[30] & b[101])^(a[29] & b[102])^(a[28] & b[103])^(a[27] & b[104])^(a[26] & b[105])^(a[25] & b[106])^(a[24] & b[107])^(a[23] & b[108])^(a[22] & b[109])^(a[21] & b[110])^(a[20] & b[111])^(a[19] & b[112])^(a[18] & b[113])^(a[17] & b[114])^(a[16] & b[115])^(a[15] & b[116])^(a[14] & b[117])^(a[13] & b[118])^(a[12] & b[119])^(a[11] & b[120])^(a[10] & b[121])^(a[9] & b[122])^(a[8] & b[123])^(a[7] & b[124])^(a[6] & b[125])^(a[5] & b[126])^(a[4] & b[127])^(a[3] & b[128])^(a[2] & b[129])^(a[1] & b[130])^(a[0] & b[131]);
assign y[132] = (a[132] & b[0])^(a[131] & b[1])^(a[130] & b[2])^(a[129] & b[3])^(a[128] & b[4])^(a[127] & b[5])^(a[126] & b[6])^(a[125] & b[7])^(a[124] & b[8])^(a[123] & b[9])^(a[122] & b[10])^(a[121] & b[11])^(a[120] & b[12])^(a[119] & b[13])^(a[118] & b[14])^(a[117] & b[15])^(a[116] & b[16])^(a[115] & b[17])^(a[114] & b[18])^(a[113] & b[19])^(a[112] & b[20])^(a[111] & b[21])^(a[110] & b[22])^(a[109] & b[23])^(a[108] & b[24])^(a[107] & b[25])^(a[106] & b[26])^(a[105] & b[27])^(a[104] & b[28])^(a[103] & b[29])^(a[102] & b[30])^(a[101] & b[31])^(a[100] & b[32])^(a[99] & b[33])^(a[98] & b[34])^(a[97] & b[35])^(a[96] & b[36])^(a[95] & b[37])^(a[94] & b[38])^(a[93] & b[39])^(a[92] & b[40])^(a[91] & b[41])^(a[90] & b[42])^(a[89] & b[43])^(a[88] & b[44])^(a[87] & b[45])^(a[86] & b[46])^(a[85] & b[47])^(a[84] & b[48])^(a[83] & b[49])^(a[82] & b[50])^(a[81] & b[51])^(a[80] & b[52])^(a[79] & b[53])^(a[78] & b[54])^(a[77] & b[55])^(a[76] & b[56])^(a[75] & b[57])^(a[74] & b[58])^(a[73] & b[59])^(a[72] & b[60])^(a[71] & b[61])^(a[70] & b[62])^(a[69] & b[63])^(a[68] & b[64])^(a[67] & b[65])^(a[66] & b[66])^(a[65] & b[67])^(a[64] & b[68])^(a[63] & b[69])^(a[62] & b[70])^(a[61] & b[71])^(a[60] & b[72])^(a[59] & b[73])^(a[58] & b[74])^(a[57] & b[75])^(a[56] & b[76])^(a[55] & b[77])^(a[54] & b[78])^(a[53] & b[79])^(a[52] & b[80])^(a[51] & b[81])^(a[50] & b[82])^(a[49] & b[83])^(a[48] & b[84])^(a[47] & b[85])^(a[46] & b[86])^(a[45] & b[87])^(a[44] & b[88])^(a[43] & b[89])^(a[42] & b[90])^(a[41] & b[91])^(a[40] & b[92])^(a[39] & b[93])^(a[38] & b[94])^(a[37] & b[95])^(a[36] & b[96])^(a[35] & b[97])^(a[34] & b[98])^(a[33] & b[99])^(a[32] & b[100])^(a[31] & b[101])^(a[30] & b[102])^(a[29] & b[103])^(a[28] & b[104])^(a[27] & b[105])^(a[26] & b[106])^(a[25] & b[107])^(a[24] & b[108])^(a[23] & b[109])^(a[22] & b[110])^(a[21] & b[111])^(a[20] & b[112])^(a[19] & b[113])^(a[18] & b[114])^(a[17] & b[115])^(a[16] & b[116])^(a[15] & b[117])^(a[14] & b[118])^(a[13] & b[119])^(a[12] & b[120])^(a[11] & b[121])^(a[10] & b[122])^(a[9] & b[123])^(a[8] & b[124])^(a[7] & b[125])^(a[6] & b[126])^(a[5] & b[127])^(a[4] & b[128])^(a[3] & b[129])^(a[2] & b[130])^(a[1] & b[131])^(a[0] & b[132]);
assign y[133] = (a[133] & b[0])^(a[132] & b[1])^(a[131] & b[2])^(a[130] & b[3])^(a[129] & b[4])^(a[128] & b[5])^(a[127] & b[6])^(a[126] & b[7])^(a[125] & b[8])^(a[124] & b[9])^(a[123] & b[10])^(a[122] & b[11])^(a[121] & b[12])^(a[120] & b[13])^(a[119] & b[14])^(a[118] & b[15])^(a[117] & b[16])^(a[116] & b[17])^(a[115] & b[18])^(a[114] & b[19])^(a[113] & b[20])^(a[112] & b[21])^(a[111] & b[22])^(a[110] & b[23])^(a[109] & b[24])^(a[108] & b[25])^(a[107] & b[26])^(a[106] & b[27])^(a[105] & b[28])^(a[104] & b[29])^(a[103] & b[30])^(a[102] & b[31])^(a[101] & b[32])^(a[100] & b[33])^(a[99] & b[34])^(a[98] & b[35])^(a[97] & b[36])^(a[96] & b[37])^(a[95] & b[38])^(a[94] & b[39])^(a[93] & b[40])^(a[92] & b[41])^(a[91] & b[42])^(a[90] & b[43])^(a[89] & b[44])^(a[88] & b[45])^(a[87] & b[46])^(a[86] & b[47])^(a[85] & b[48])^(a[84] & b[49])^(a[83] & b[50])^(a[82] & b[51])^(a[81] & b[52])^(a[80] & b[53])^(a[79] & b[54])^(a[78] & b[55])^(a[77] & b[56])^(a[76] & b[57])^(a[75] & b[58])^(a[74] & b[59])^(a[73] & b[60])^(a[72] & b[61])^(a[71] & b[62])^(a[70] & b[63])^(a[69] & b[64])^(a[68] & b[65])^(a[67] & b[66])^(a[66] & b[67])^(a[65] & b[68])^(a[64] & b[69])^(a[63] & b[70])^(a[62] & b[71])^(a[61] & b[72])^(a[60] & b[73])^(a[59] & b[74])^(a[58] & b[75])^(a[57] & b[76])^(a[56] & b[77])^(a[55] & b[78])^(a[54] & b[79])^(a[53] & b[80])^(a[52] & b[81])^(a[51] & b[82])^(a[50] & b[83])^(a[49] & b[84])^(a[48] & b[85])^(a[47] & b[86])^(a[46] & b[87])^(a[45] & b[88])^(a[44] & b[89])^(a[43] & b[90])^(a[42] & b[91])^(a[41] & b[92])^(a[40] & b[93])^(a[39] & b[94])^(a[38] & b[95])^(a[37] & b[96])^(a[36] & b[97])^(a[35] & b[98])^(a[34] & b[99])^(a[33] & b[100])^(a[32] & b[101])^(a[31] & b[102])^(a[30] & b[103])^(a[29] & b[104])^(a[28] & b[105])^(a[27] & b[106])^(a[26] & b[107])^(a[25] & b[108])^(a[24] & b[109])^(a[23] & b[110])^(a[22] & b[111])^(a[21] & b[112])^(a[20] & b[113])^(a[19] & b[114])^(a[18] & b[115])^(a[17] & b[116])^(a[16] & b[117])^(a[15] & b[118])^(a[14] & b[119])^(a[13] & b[120])^(a[12] & b[121])^(a[11] & b[122])^(a[10] & b[123])^(a[9] & b[124])^(a[8] & b[125])^(a[7] & b[126])^(a[6] & b[127])^(a[5] & b[128])^(a[4] & b[129])^(a[3] & b[130])^(a[2] & b[131])^(a[1] & b[132])^(a[0] & b[133]);
assign y[134] = (a[134] & b[0])^(a[133] & b[1])^(a[132] & b[2])^(a[131] & b[3])^(a[130] & b[4])^(a[129] & b[5])^(a[128] & b[6])^(a[127] & b[7])^(a[126] & b[8])^(a[125] & b[9])^(a[124] & b[10])^(a[123] & b[11])^(a[122] & b[12])^(a[121] & b[13])^(a[120] & b[14])^(a[119] & b[15])^(a[118] & b[16])^(a[117] & b[17])^(a[116] & b[18])^(a[115] & b[19])^(a[114] & b[20])^(a[113] & b[21])^(a[112] & b[22])^(a[111] & b[23])^(a[110] & b[24])^(a[109] & b[25])^(a[108] & b[26])^(a[107] & b[27])^(a[106] & b[28])^(a[105] & b[29])^(a[104] & b[30])^(a[103] & b[31])^(a[102] & b[32])^(a[101] & b[33])^(a[100] & b[34])^(a[99] & b[35])^(a[98] & b[36])^(a[97] & b[37])^(a[96] & b[38])^(a[95] & b[39])^(a[94] & b[40])^(a[93] & b[41])^(a[92] & b[42])^(a[91] & b[43])^(a[90] & b[44])^(a[89] & b[45])^(a[88] & b[46])^(a[87] & b[47])^(a[86] & b[48])^(a[85] & b[49])^(a[84] & b[50])^(a[83] & b[51])^(a[82] & b[52])^(a[81] & b[53])^(a[80] & b[54])^(a[79] & b[55])^(a[78] & b[56])^(a[77] & b[57])^(a[76] & b[58])^(a[75] & b[59])^(a[74] & b[60])^(a[73] & b[61])^(a[72] & b[62])^(a[71] & b[63])^(a[70] & b[64])^(a[69] & b[65])^(a[68] & b[66])^(a[67] & b[67])^(a[66] & b[68])^(a[65] & b[69])^(a[64] & b[70])^(a[63] & b[71])^(a[62] & b[72])^(a[61] & b[73])^(a[60] & b[74])^(a[59] & b[75])^(a[58] & b[76])^(a[57] & b[77])^(a[56] & b[78])^(a[55] & b[79])^(a[54] & b[80])^(a[53] & b[81])^(a[52] & b[82])^(a[51] & b[83])^(a[50] & b[84])^(a[49] & b[85])^(a[48] & b[86])^(a[47] & b[87])^(a[46] & b[88])^(a[45] & b[89])^(a[44] & b[90])^(a[43] & b[91])^(a[42] & b[92])^(a[41] & b[93])^(a[40] & b[94])^(a[39] & b[95])^(a[38] & b[96])^(a[37] & b[97])^(a[36] & b[98])^(a[35] & b[99])^(a[34] & b[100])^(a[33] & b[101])^(a[32] & b[102])^(a[31] & b[103])^(a[30] & b[104])^(a[29] & b[105])^(a[28] & b[106])^(a[27] & b[107])^(a[26] & b[108])^(a[25] & b[109])^(a[24] & b[110])^(a[23] & b[111])^(a[22] & b[112])^(a[21] & b[113])^(a[20] & b[114])^(a[19] & b[115])^(a[18] & b[116])^(a[17] & b[117])^(a[16] & b[118])^(a[15] & b[119])^(a[14] & b[120])^(a[13] & b[121])^(a[12] & b[122])^(a[11] & b[123])^(a[10] & b[124])^(a[9] & b[125])^(a[8] & b[126])^(a[7] & b[127])^(a[6] & b[128])^(a[5] & b[129])^(a[4] & b[130])^(a[3] & b[131])^(a[2] & b[132])^(a[1] & b[133])^(a[0] & b[134]);
assign y[135] = (a[135] & b[0])^(a[134] & b[1])^(a[133] & b[2])^(a[132] & b[3])^(a[131] & b[4])^(a[130] & b[5])^(a[129] & b[6])^(a[128] & b[7])^(a[127] & b[8])^(a[126] & b[9])^(a[125] & b[10])^(a[124] & b[11])^(a[123] & b[12])^(a[122] & b[13])^(a[121] & b[14])^(a[120] & b[15])^(a[119] & b[16])^(a[118] & b[17])^(a[117] & b[18])^(a[116] & b[19])^(a[115] & b[20])^(a[114] & b[21])^(a[113] & b[22])^(a[112] & b[23])^(a[111] & b[24])^(a[110] & b[25])^(a[109] & b[26])^(a[108] & b[27])^(a[107] & b[28])^(a[106] & b[29])^(a[105] & b[30])^(a[104] & b[31])^(a[103] & b[32])^(a[102] & b[33])^(a[101] & b[34])^(a[100] & b[35])^(a[99] & b[36])^(a[98] & b[37])^(a[97] & b[38])^(a[96] & b[39])^(a[95] & b[40])^(a[94] & b[41])^(a[93] & b[42])^(a[92] & b[43])^(a[91] & b[44])^(a[90] & b[45])^(a[89] & b[46])^(a[88] & b[47])^(a[87] & b[48])^(a[86] & b[49])^(a[85] & b[50])^(a[84] & b[51])^(a[83] & b[52])^(a[82] & b[53])^(a[81] & b[54])^(a[80] & b[55])^(a[79] & b[56])^(a[78] & b[57])^(a[77] & b[58])^(a[76] & b[59])^(a[75] & b[60])^(a[74] & b[61])^(a[73] & b[62])^(a[72] & b[63])^(a[71] & b[64])^(a[70] & b[65])^(a[69] & b[66])^(a[68] & b[67])^(a[67] & b[68])^(a[66] & b[69])^(a[65] & b[70])^(a[64] & b[71])^(a[63] & b[72])^(a[62] & b[73])^(a[61] & b[74])^(a[60] & b[75])^(a[59] & b[76])^(a[58] & b[77])^(a[57] & b[78])^(a[56] & b[79])^(a[55] & b[80])^(a[54] & b[81])^(a[53] & b[82])^(a[52] & b[83])^(a[51] & b[84])^(a[50] & b[85])^(a[49] & b[86])^(a[48] & b[87])^(a[47] & b[88])^(a[46] & b[89])^(a[45] & b[90])^(a[44] & b[91])^(a[43] & b[92])^(a[42] & b[93])^(a[41] & b[94])^(a[40] & b[95])^(a[39] & b[96])^(a[38] & b[97])^(a[37] & b[98])^(a[36] & b[99])^(a[35] & b[100])^(a[34] & b[101])^(a[33] & b[102])^(a[32] & b[103])^(a[31] & b[104])^(a[30] & b[105])^(a[29] & b[106])^(a[28] & b[107])^(a[27] & b[108])^(a[26] & b[109])^(a[25] & b[110])^(a[24] & b[111])^(a[23] & b[112])^(a[22] & b[113])^(a[21] & b[114])^(a[20] & b[115])^(a[19] & b[116])^(a[18] & b[117])^(a[17] & b[118])^(a[16] & b[119])^(a[15] & b[120])^(a[14] & b[121])^(a[13] & b[122])^(a[12] & b[123])^(a[11] & b[124])^(a[10] & b[125])^(a[9] & b[126])^(a[8] & b[127])^(a[7] & b[128])^(a[6] & b[129])^(a[5] & b[130])^(a[4] & b[131])^(a[3] & b[132])^(a[2] & b[133])^(a[1] & b[134])^(a[0] & b[135]);
assign y[136] = (a[136] & b[0])^(a[135] & b[1])^(a[134] & b[2])^(a[133] & b[3])^(a[132] & b[4])^(a[131] & b[5])^(a[130] & b[6])^(a[129] & b[7])^(a[128] & b[8])^(a[127] & b[9])^(a[126] & b[10])^(a[125] & b[11])^(a[124] & b[12])^(a[123] & b[13])^(a[122] & b[14])^(a[121] & b[15])^(a[120] & b[16])^(a[119] & b[17])^(a[118] & b[18])^(a[117] & b[19])^(a[116] & b[20])^(a[115] & b[21])^(a[114] & b[22])^(a[113] & b[23])^(a[112] & b[24])^(a[111] & b[25])^(a[110] & b[26])^(a[109] & b[27])^(a[108] & b[28])^(a[107] & b[29])^(a[106] & b[30])^(a[105] & b[31])^(a[104] & b[32])^(a[103] & b[33])^(a[102] & b[34])^(a[101] & b[35])^(a[100] & b[36])^(a[99] & b[37])^(a[98] & b[38])^(a[97] & b[39])^(a[96] & b[40])^(a[95] & b[41])^(a[94] & b[42])^(a[93] & b[43])^(a[92] & b[44])^(a[91] & b[45])^(a[90] & b[46])^(a[89] & b[47])^(a[88] & b[48])^(a[87] & b[49])^(a[86] & b[50])^(a[85] & b[51])^(a[84] & b[52])^(a[83] & b[53])^(a[82] & b[54])^(a[81] & b[55])^(a[80] & b[56])^(a[79] & b[57])^(a[78] & b[58])^(a[77] & b[59])^(a[76] & b[60])^(a[75] & b[61])^(a[74] & b[62])^(a[73] & b[63])^(a[72] & b[64])^(a[71] & b[65])^(a[70] & b[66])^(a[69] & b[67])^(a[68] & b[68])^(a[67] & b[69])^(a[66] & b[70])^(a[65] & b[71])^(a[64] & b[72])^(a[63] & b[73])^(a[62] & b[74])^(a[61] & b[75])^(a[60] & b[76])^(a[59] & b[77])^(a[58] & b[78])^(a[57] & b[79])^(a[56] & b[80])^(a[55] & b[81])^(a[54] & b[82])^(a[53] & b[83])^(a[52] & b[84])^(a[51] & b[85])^(a[50] & b[86])^(a[49] & b[87])^(a[48] & b[88])^(a[47] & b[89])^(a[46] & b[90])^(a[45] & b[91])^(a[44] & b[92])^(a[43] & b[93])^(a[42] & b[94])^(a[41] & b[95])^(a[40] & b[96])^(a[39] & b[97])^(a[38] & b[98])^(a[37] & b[99])^(a[36] & b[100])^(a[35] & b[101])^(a[34] & b[102])^(a[33] & b[103])^(a[32] & b[104])^(a[31] & b[105])^(a[30] & b[106])^(a[29] & b[107])^(a[28] & b[108])^(a[27] & b[109])^(a[26] & b[110])^(a[25] & b[111])^(a[24] & b[112])^(a[23] & b[113])^(a[22] & b[114])^(a[21] & b[115])^(a[20] & b[116])^(a[19] & b[117])^(a[18] & b[118])^(a[17] & b[119])^(a[16] & b[120])^(a[15] & b[121])^(a[14] & b[122])^(a[13] & b[123])^(a[12] & b[124])^(a[11] & b[125])^(a[10] & b[126])^(a[9] & b[127])^(a[8] & b[128])^(a[7] & b[129])^(a[6] & b[130])^(a[5] & b[131])^(a[4] & b[132])^(a[3] & b[133])^(a[2] & b[134])^(a[1] & b[135])^(a[0] & b[136]);
assign y[137] = (a[137] & b[0])^(a[136] & b[1])^(a[135] & b[2])^(a[134] & b[3])^(a[133] & b[4])^(a[132] & b[5])^(a[131] & b[6])^(a[130] & b[7])^(a[129] & b[8])^(a[128] & b[9])^(a[127] & b[10])^(a[126] & b[11])^(a[125] & b[12])^(a[124] & b[13])^(a[123] & b[14])^(a[122] & b[15])^(a[121] & b[16])^(a[120] & b[17])^(a[119] & b[18])^(a[118] & b[19])^(a[117] & b[20])^(a[116] & b[21])^(a[115] & b[22])^(a[114] & b[23])^(a[113] & b[24])^(a[112] & b[25])^(a[111] & b[26])^(a[110] & b[27])^(a[109] & b[28])^(a[108] & b[29])^(a[107] & b[30])^(a[106] & b[31])^(a[105] & b[32])^(a[104] & b[33])^(a[103] & b[34])^(a[102] & b[35])^(a[101] & b[36])^(a[100] & b[37])^(a[99] & b[38])^(a[98] & b[39])^(a[97] & b[40])^(a[96] & b[41])^(a[95] & b[42])^(a[94] & b[43])^(a[93] & b[44])^(a[92] & b[45])^(a[91] & b[46])^(a[90] & b[47])^(a[89] & b[48])^(a[88] & b[49])^(a[87] & b[50])^(a[86] & b[51])^(a[85] & b[52])^(a[84] & b[53])^(a[83] & b[54])^(a[82] & b[55])^(a[81] & b[56])^(a[80] & b[57])^(a[79] & b[58])^(a[78] & b[59])^(a[77] & b[60])^(a[76] & b[61])^(a[75] & b[62])^(a[74] & b[63])^(a[73] & b[64])^(a[72] & b[65])^(a[71] & b[66])^(a[70] & b[67])^(a[69] & b[68])^(a[68] & b[69])^(a[67] & b[70])^(a[66] & b[71])^(a[65] & b[72])^(a[64] & b[73])^(a[63] & b[74])^(a[62] & b[75])^(a[61] & b[76])^(a[60] & b[77])^(a[59] & b[78])^(a[58] & b[79])^(a[57] & b[80])^(a[56] & b[81])^(a[55] & b[82])^(a[54] & b[83])^(a[53] & b[84])^(a[52] & b[85])^(a[51] & b[86])^(a[50] & b[87])^(a[49] & b[88])^(a[48] & b[89])^(a[47] & b[90])^(a[46] & b[91])^(a[45] & b[92])^(a[44] & b[93])^(a[43] & b[94])^(a[42] & b[95])^(a[41] & b[96])^(a[40] & b[97])^(a[39] & b[98])^(a[38] & b[99])^(a[37] & b[100])^(a[36] & b[101])^(a[35] & b[102])^(a[34] & b[103])^(a[33] & b[104])^(a[32] & b[105])^(a[31] & b[106])^(a[30] & b[107])^(a[29] & b[108])^(a[28] & b[109])^(a[27] & b[110])^(a[26] & b[111])^(a[25] & b[112])^(a[24] & b[113])^(a[23] & b[114])^(a[22] & b[115])^(a[21] & b[116])^(a[20] & b[117])^(a[19] & b[118])^(a[18] & b[119])^(a[17] & b[120])^(a[16] & b[121])^(a[15] & b[122])^(a[14] & b[123])^(a[13] & b[124])^(a[12] & b[125])^(a[11] & b[126])^(a[10] & b[127])^(a[9] & b[128])^(a[8] & b[129])^(a[7] & b[130])^(a[6] & b[131])^(a[5] & b[132])^(a[4] & b[133])^(a[3] & b[134])^(a[2] & b[135])^(a[1] & b[136])^(a[0] & b[137]);
assign y[138] = (a[138] & b[0])^(a[137] & b[1])^(a[136] & b[2])^(a[135] & b[3])^(a[134] & b[4])^(a[133] & b[5])^(a[132] & b[6])^(a[131] & b[7])^(a[130] & b[8])^(a[129] & b[9])^(a[128] & b[10])^(a[127] & b[11])^(a[126] & b[12])^(a[125] & b[13])^(a[124] & b[14])^(a[123] & b[15])^(a[122] & b[16])^(a[121] & b[17])^(a[120] & b[18])^(a[119] & b[19])^(a[118] & b[20])^(a[117] & b[21])^(a[116] & b[22])^(a[115] & b[23])^(a[114] & b[24])^(a[113] & b[25])^(a[112] & b[26])^(a[111] & b[27])^(a[110] & b[28])^(a[109] & b[29])^(a[108] & b[30])^(a[107] & b[31])^(a[106] & b[32])^(a[105] & b[33])^(a[104] & b[34])^(a[103] & b[35])^(a[102] & b[36])^(a[101] & b[37])^(a[100] & b[38])^(a[99] & b[39])^(a[98] & b[40])^(a[97] & b[41])^(a[96] & b[42])^(a[95] & b[43])^(a[94] & b[44])^(a[93] & b[45])^(a[92] & b[46])^(a[91] & b[47])^(a[90] & b[48])^(a[89] & b[49])^(a[88] & b[50])^(a[87] & b[51])^(a[86] & b[52])^(a[85] & b[53])^(a[84] & b[54])^(a[83] & b[55])^(a[82] & b[56])^(a[81] & b[57])^(a[80] & b[58])^(a[79] & b[59])^(a[78] & b[60])^(a[77] & b[61])^(a[76] & b[62])^(a[75] & b[63])^(a[74] & b[64])^(a[73] & b[65])^(a[72] & b[66])^(a[71] & b[67])^(a[70] & b[68])^(a[69] & b[69])^(a[68] & b[70])^(a[67] & b[71])^(a[66] & b[72])^(a[65] & b[73])^(a[64] & b[74])^(a[63] & b[75])^(a[62] & b[76])^(a[61] & b[77])^(a[60] & b[78])^(a[59] & b[79])^(a[58] & b[80])^(a[57] & b[81])^(a[56] & b[82])^(a[55] & b[83])^(a[54] & b[84])^(a[53] & b[85])^(a[52] & b[86])^(a[51] & b[87])^(a[50] & b[88])^(a[49] & b[89])^(a[48] & b[90])^(a[47] & b[91])^(a[46] & b[92])^(a[45] & b[93])^(a[44] & b[94])^(a[43] & b[95])^(a[42] & b[96])^(a[41] & b[97])^(a[40] & b[98])^(a[39] & b[99])^(a[38] & b[100])^(a[37] & b[101])^(a[36] & b[102])^(a[35] & b[103])^(a[34] & b[104])^(a[33] & b[105])^(a[32] & b[106])^(a[31] & b[107])^(a[30] & b[108])^(a[29] & b[109])^(a[28] & b[110])^(a[27] & b[111])^(a[26] & b[112])^(a[25] & b[113])^(a[24] & b[114])^(a[23] & b[115])^(a[22] & b[116])^(a[21] & b[117])^(a[20] & b[118])^(a[19] & b[119])^(a[18] & b[120])^(a[17] & b[121])^(a[16] & b[122])^(a[15] & b[123])^(a[14] & b[124])^(a[13] & b[125])^(a[12] & b[126])^(a[11] & b[127])^(a[10] & b[128])^(a[9] & b[129])^(a[8] & b[130])^(a[7] & b[131])^(a[6] & b[132])^(a[5] & b[133])^(a[4] & b[134])^(a[3] & b[135])^(a[2] & b[136])^(a[1] & b[137])^(a[0] & b[138]);
assign y[139] = (a[139] & b[0])^(a[138] & b[1])^(a[137] & b[2])^(a[136] & b[3])^(a[135] & b[4])^(a[134] & b[5])^(a[133] & b[6])^(a[132] & b[7])^(a[131] & b[8])^(a[130] & b[9])^(a[129] & b[10])^(a[128] & b[11])^(a[127] & b[12])^(a[126] & b[13])^(a[125] & b[14])^(a[124] & b[15])^(a[123] & b[16])^(a[122] & b[17])^(a[121] & b[18])^(a[120] & b[19])^(a[119] & b[20])^(a[118] & b[21])^(a[117] & b[22])^(a[116] & b[23])^(a[115] & b[24])^(a[114] & b[25])^(a[113] & b[26])^(a[112] & b[27])^(a[111] & b[28])^(a[110] & b[29])^(a[109] & b[30])^(a[108] & b[31])^(a[107] & b[32])^(a[106] & b[33])^(a[105] & b[34])^(a[104] & b[35])^(a[103] & b[36])^(a[102] & b[37])^(a[101] & b[38])^(a[100] & b[39])^(a[99] & b[40])^(a[98] & b[41])^(a[97] & b[42])^(a[96] & b[43])^(a[95] & b[44])^(a[94] & b[45])^(a[93] & b[46])^(a[92] & b[47])^(a[91] & b[48])^(a[90] & b[49])^(a[89] & b[50])^(a[88] & b[51])^(a[87] & b[52])^(a[86] & b[53])^(a[85] & b[54])^(a[84] & b[55])^(a[83] & b[56])^(a[82] & b[57])^(a[81] & b[58])^(a[80] & b[59])^(a[79] & b[60])^(a[78] & b[61])^(a[77] & b[62])^(a[76] & b[63])^(a[75] & b[64])^(a[74] & b[65])^(a[73] & b[66])^(a[72] & b[67])^(a[71] & b[68])^(a[70] & b[69])^(a[69] & b[70])^(a[68] & b[71])^(a[67] & b[72])^(a[66] & b[73])^(a[65] & b[74])^(a[64] & b[75])^(a[63] & b[76])^(a[62] & b[77])^(a[61] & b[78])^(a[60] & b[79])^(a[59] & b[80])^(a[58] & b[81])^(a[57] & b[82])^(a[56] & b[83])^(a[55] & b[84])^(a[54] & b[85])^(a[53] & b[86])^(a[52] & b[87])^(a[51] & b[88])^(a[50] & b[89])^(a[49] & b[90])^(a[48] & b[91])^(a[47] & b[92])^(a[46] & b[93])^(a[45] & b[94])^(a[44] & b[95])^(a[43] & b[96])^(a[42] & b[97])^(a[41] & b[98])^(a[40] & b[99])^(a[39] & b[100])^(a[38] & b[101])^(a[37] & b[102])^(a[36] & b[103])^(a[35] & b[104])^(a[34] & b[105])^(a[33] & b[106])^(a[32] & b[107])^(a[31] & b[108])^(a[30] & b[109])^(a[29] & b[110])^(a[28] & b[111])^(a[27] & b[112])^(a[26] & b[113])^(a[25] & b[114])^(a[24] & b[115])^(a[23] & b[116])^(a[22] & b[117])^(a[21] & b[118])^(a[20] & b[119])^(a[19] & b[120])^(a[18] & b[121])^(a[17] & b[122])^(a[16] & b[123])^(a[15] & b[124])^(a[14] & b[125])^(a[13] & b[126])^(a[12] & b[127])^(a[11] & b[128])^(a[10] & b[129])^(a[9] & b[130])^(a[8] & b[131])^(a[7] & b[132])^(a[6] & b[133])^(a[5] & b[134])^(a[4] & b[135])^(a[3] & b[136])^(a[2] & b[137])^(a[1] & b[138])^(a[0] & b[139]);
assign y[140] = (a[140] & b[0])^(a[139] & b[1])^(a[138] & b[2])^(a[137] & b[3])^(a[136] & b[4])^(a[135] & b[5])^(a[134] & b[6])^(a[133] & b[7])^(a[132] & b[8])^(a[131] & b[9])^(a[130] & b[10])^(a[129] & b[11])^(a[128] & b[12])^(a[127] & b[13])^(a[126] & b[14])^(a[125] & b[15])^(a[124] & b[16])^(a[123] & b[17])^(a[122] & b[18])^(a[121] & b[19])^(a[120] & b[20])^(a[119] & b[21])^(a[118] & b[22])^(a[117] & b[23])^(a[116] & b[24])^(a[115] & b[25])^(a[114] & b[26])^(a[113] & b[27])^(a[112] & b[28])^(a[111] & b[29])^(a[110] & b[30])^(a[109] & b[31])^(a[108] & b[32])^(a[107] & b[33])^(a[106] & b[34])^(a[105] & b[35])^(a[104] & b[36])^(a[103] & b[37])^(a[102] & b[38])^(a[101] & b[39])^(a[100] & b[40])^(a[99] & b[41])^(a[98] & b[42])^(a[97] & b[43])^(a[96] & b[44])^(a[95] & b[45])^(a[94] & b[46])^(a[93] & b[47])^(a[92] & b[48])^(a[91] & b[49])^(a[90] & b[50])^(a[89] & b[51])^(a[88] & b[52])^(a[87] & b[53])^(a[86] & b[54])^(a[85] & b[55])^(a[84] & b[56])^(a[83] & b[57])^(a[82] & b[58])^(a[81] & b[59])^(a[80] & b[60])^(a[79] & b[61])^(a[78] & b[62])^(a[77] & b[63])^(a[76] & b[64])^(a[75] & b[65])^(a[74] & b[66])^(a[73] & b[67])^(a[72] & b[68])^(a[71] & b[69])^(a[70] & b[70])^(a[69] & b[71])^(a[68] & b[72])^(a[67] & b[73])^(a[66] & b[74])^(a[65] & b[75])^(a[64] & b[76])^(a[63] & b[77])^(a[62] & b[78])^(a[61] & b[79])^(a[60] & b[80])^(a[59] & b[81])^(a[58] & b[82])^(a[57] & b[83])^(a[56] & b[84])^(a[55] & b[85])^(a[54] & b[86])^(a[53] & b[87])^(a[52] & b[88])^(a[51] & b[89])^(a[50] & b[90])^(a[49] & b[91])^(a[48] & b[92])^(a[47] & b[93])^(a[46] & b[94])^(a[45] & b[95])^(a[44] & b[96])^(a[43] & b[97])^(a[42] & b[98])^(a[41] & b[99])^(a[40] & b[100])^(a[39] & b[101])^(a[38] & b[102])^(a[37] & b[103])^(a[36] & b[104])^(a[35] & b[105])^(a[34] & b[106])^(a[33] & b[107])^(a[32] & b[108])^(a[31] & b[109])^(a[30] & b[110])^(a[29] & b[111])^(a[28] & b[112])^(a[27] & b[113])^(a[26] & b[114])^(a[25] & b[115])^(a[24] & b[116])^(a[23] & b[117])^(a[22] & b[118])^(a[21] & b[119])^(a[20] & b[120])^(a[19] & b[121])^(a[18] & b[122])^(a[17] & b[123])^(a[16] & b[124])^(a[15] & b[125])^(a[14] & b[126])^(a[13] & b[127])^(a[12] & b[128])^(a[11] & b[129])^(a[10] & b[130])^(a[9] & b[131])^(a[8] & b[132])^(a[7] & b[133])^(a[6] & b[134])^(a[5] & b[135])^(a[4] & b[136])^(a[3] & b[137])^(a[2] & b[138])^(a[1] & b[139])^(a[0] & b[140]);
assign y[141] = (a[141] & b[0])^(a[140] & b[1])^(a[139] & b[2])^(a[138] & b[3])^(a[137] & b[4])^(a[136] & b[5])^(a[135] & b[6])^(a[134] & b[7])^(a[133] & b[8])^(a[132] & b[9])^(a[131] & b[10])^(a[130] & b[11])^(a[129] & b[12])^(a[128] & b[13])^(a[127] & b[14])^(a[126] & b[15])^(a[125] & b[16])^(a[124] & b[17])^(a[123] & b[18])^(a[122] & b[19])^(a[121] & b[20])^(a[120] & b[21])^(a[119] & b[22])^(a[118] & b[23])^(a[117] & b[24])^(a[116] & b[25])^(a[115] & b[26])^(a[114] & b[27])^(a[113] & b[28])^(a[112] & b[29])^(a[111] & b[30])^(a[110] & b[31])^(a[109] & b[32])^(a[108] & b[33])^(a[107] & b[34])^(a[106] & b[35])^(a[105] & b[36])^(a[104] & b[37])^(a[103] & b[38])^(a[102] & b[39])^(a[101] & b[40])^(a[100] & b[41])^(a[99] & b[42])^(a[98] & b[43])^(a[97] & b[44])^(a[96] & b[45])^(a[95] & b[46])^(a[94] & b[47])^(a[93] & b[48])^(a[92] & b[49])^(a[91] & b[50])^(a[90] & b[51])^(a[89] & b[52])^(a[88] & b[53])^(a[87] & b[54])^(a[86] & b[55])^(a[85] & b[56])^(a[84] & b[57])^(a[83] & b[58])^(a[82] & b[59])^(a[81] & b[60])^(a[80] & b[61])^(a[79] & b[62])^(a[78] & b[63])^(a[77] & b[64])^(a[76] & b[65])^(a[75] & b[66])^(a[74] & b[67])^(a[73] & b[68])^(a[72] & b[69])^(a[71] & b[70])^(a[70] & b[71])^(a[69] & b[72])^(a[68] & b[73])^(a[67] & b[74])^(a[66] & b[75])^(a[65] & b[76])^(a[64] & b[77])^(a[63] & b[78])^(a[62] & b[79])^(a[61] & b[80])^(a[60] & b[81])^(a[59] & b[82])^(a[58] & b[83])^(a[57] & b[84])^(a[56] & b[85])^(a[55] & b[86])^(a[54] & b[87])^(a[53] & b[88])^(a[52] & b[89])^(a[51] & b[90])^(a[50] & b[91])^(a[49] & b[92])^(a[48] & b[93])^(a[47] & b[94])^(a[46] & b[95])^(a[45] & b[96])^(a[44] & b[97])^(a[43] & b[98])^(a[42] & b[99])^(a[41] & b[100])^(a[40] & b[101])^(a[39] & b[102])^(a[38] & b[103])^(a[37] & b[104])^(a[36] & b[105])^(a[35] & b[106])^(a[34] & b[107])^(a[33] & b[108])^(a[32] & b[109])^(a[31] & b[110])^(a[30] & b[111])^(a[29] & b[112])^(a[28] & b[113])^(a[27] & b[114])^(a[26] & b[115])^(a[25] & b[116])^(a[24] & b[117])^(a[23] & b[118])^(a[22] & b[119])^(a[21] & b[120])^(a[20] & b[121])^(a[19] & b[122])^(a[18] & b[123])^(a[17] & b[124])^(a[16] & b[125])^(a[15] & b[126])^(a[14] & b[127])^(a[13] & b[128])^(a[12] & b[129])^(a[11] & b[130])^(a[10] & b[131])^(a[9] & b[132])^(a[8] & b[133])^(a[7] & b[134])^(a[6] & b[135])^(a[5] & b[136])^(a[4] & b[137])^(a[3] & b[138])^(a[2] & b[139])^(a[1] & b[140])^(a[0] & b[141]);
assign y[142] = (a[142] & b[0])^(a[141] & b[1])^(a[140] & b[2])^(a[139] & b[3])^(a[138] & b[4])^(a[137] & b[5])^(a[136] & b[6])^(a[135] & b[7])^(a[134] & b[8])^(a[133] & b[9])^(a[132] & b[10])^(a[131] & b[11])^(a[130] & b[12])^(a[129] & b[13])^(a[128] & b[14])^(a[127] & b[15])^(a[126] & b[16])^(a[125] & b[17])^(a[124] & b[18])^(a[123] & b[19])^(a[122] & b[20])^(a[121] & b[21])^(a[120] & b[22])^(a[119] & b[23])^(a[118] & b[24])^(a[117] & b[25])^(a[116] & b[26])^(a[115] & b[27])^(a[114] & b[28])^(a[113] & b[29])^(a[112] & b[30])^(a[111] & b[31])^(a[110] & b[32])^(a[109] & b[33])^(a[108] & b[34])^(a[107] & b[35])^(a[106] & b[36])^(a[105] & b[37])^(a[104] & b[38])^(a[103] & b[39])^(a[102] & b[40])^(a[101] & b[41])^(a[100] & b[42])^(a[99] & b[43])^(a[98] & b[44])^(a[97] & b[45])^(a[96] & b[46])^(a[95] & b[47])^(a[94] & b[48])^(a[93] & b[49])^(a[92] & b[50])^(a[91] & b[51])^(a[90] & b[52])^(a[89] & b[53])^(a[88] & b[54])^(a[87] & b[55])^(a[86] & b[56])^(a[85] & b[57])^(a[84] & b[58])^(a[83] & b[59])^(a[82] & b[60])^(a[81] & b[61])^(a[80] & b[62])^(a[79] & b[63])^(a[78] & b[64])^(a[77] & b[65])^(a[76] & b[66])^(a[75] & b[67])^(a[74] & b[68])^(a[73] & b[69])^(a[72] & b[70])^(a[71] & b[71])^(a[70] & b[72])^(a[69] & b[73])^(a[68] & b[74])^(a[67] & b[75])^(a[66] & b[76])^(a[65] & b[77])^(a[64] & b[78])^(a[63] & b[79])^(a[62] & b[80])^(a[61] & b[81])^(a[60] & b[82])^(a[59] & b[83])^(a[58] & b[84])^(a[57] & b[85])^(a[56] & b[86])^(a[55] & b[87])^(a[54] & b[88])^(a[53] & b[89])^(a[52] & b[90])^(a[51] & b[91])^(a[50] & b[92])^(a[49] & b[93])^(a[48] & b[94])^(a[47] & b[95])^(a[46] & b[96])^(a[45] & b[97])^(a[44] & b[98])^(a[43] & b[99])^(a[42] & b[100])^(a[41] & b[101])^(a[40] & b[102])^(a[39] & b[103])^(a[38] & b[104])^(a[37] & b[105])^(a[36] & b[106])^(a[35] & b[107])^(a[34] & b[108])^(a[33] & b[109])^(a[32] & b[110])^(a[31] & b[111])^(a[30] & b[112])^(a[29] & b[113])^(a[28] & b[114])^(a[27] & b[115])^(a[26] & b[116])^(a[25] & b[117])^(a[24] & b[118])^(a[23] & b[119])^(a[22] & b[120])^(a[21] & b[121])^(a[20] & b[122])^(a[19] & b[123])^(a[18] & b[124])^(a[17] & b[125])^(a[16] & b[126])^(a[15] & b[127])^(a[14] & b[128])^(a[13] & b[129])^(a[12] & b[130])^(a[11] & b[131])^(a[10] & b[132])^(a[9] & b[133])^(a[8] & b[134])^(a[7] & b[135])^(a[6] & b[136])^(a[5] & b[137])^(a[4] & b[138])^(a[3] & b[139])^(a[2] & b[140])^(a[1] & b[141])^(a[0] & b[142]);
assign y[143] = (a[143] & b[0])^(a[142] & b[1])^(a[141] & b[2])^(a[140] & b[3])^(a[139] & b[4])^(a[138] & b[5])^(a[137] & b[6])^(a[136] & b[7])^(a[135] & b[8])^(a[134] & b[9])^(a[133] & b[10])^(a[132] & b[11])^(a[131] & b[12])^(a[130] & b[13])^(a[129] & b[14])^(a[128] & b[15])^(a[127] & b[16])^(a[126] & b[17])^(a[125] & b[18])^(a[124] & b[19])^(a[123] & b[20])^(a[122] & b[21])^(a[121] & b[22])^(a[120] & b[23])^(a[119] & b[24])^(a[118] & b[25])^(a[117] & b[26])^(a[116] & b[27])^(a[115] & b[28])^(a[114] & b[29])^(a[113] & b[30])^(a[112] & b[31])^(a[111] & b[32])^(a[110] & b[33])^(a[109] & b[34])^(a[108] & b[35])^(a[107] & b[36])^(a[106] & b[37])^(a[105] & b[38])^(a[104] & b[39])^(a[103] & b[40])^(a[102] & b[41])^(a[101] & b[42])^(a[100] & b[43])^(a[99] & b[44])^(a[98] & b[45])^(a[97] & b[46])^(a[96] & b[47])^(a[95] & b[48])^(a[94] & b[49])^(a[93] & b[50])^(a[92] & b[51])^(a[91] & b[52])^(a[90] & b[53])^(a[89] & b[54])^(a[88] & b[55])^(a[87] & b[56])^(a[86] & b[57])^(a[85] & b[58])^(a[84] & b[59])^(a[83] & b[60])^(a[82] & b[61])^(a[81] & b[62])^(a[80] & b[63])^(a[79] & b[64])^(a[78] & b[65])^(a[77] & b[66])^(a[76] & b[67])^(a[75] & b[68])^(a[74] & b[69])^(a[73] & b[70])^(a[72] & b[71])^(a[71] & b[72])^(a[70] & b[73])^(a[69] & b[74])^(a[68] & b[75])^(a[67] & b[76])^(a[66] & b[77])^(a[65] & b[78])^(a[64] & b[79])^(a[63] & b[80])^(a[62] & b[81])^(a[61] & b[82])^(a[60] & b[83])^(a[59] & b[84])^(a[58] & b[85])^(a[57] & b[86])^(a[56] & b[87])^(a[55] & b[88])^(a[54] & b[89])^(a[53] & b[90])^(a[52] & b[91])^(a[51] & b[92])^(a[50] & b[93])^(a[49] & b[94])^(a[48] & b[95])^(a[47] & b[96])^(a[46] & b[97])^(a[45] & b[98])^(a[44] & b[99])^(a[43] & b[100])^(a[42] & b[101])^(a[41] & b[102])^(a[40] & b[103])^(a[39] & b[104])^(a[38] & b[105])^(a[37] & b[106])^(a[36] & b[107])^(a[35] & b[108])^(a[34] & b[109])^(a[33] & b[110])^(a[32] & b[111])^(a[31] & b[112])^(a[30] & b[113])^(a[29] & b[114])^(a[28] & b[115])^(a[27] & b[116])^(a[26] & b[117])^(a[25] & b[118])^(a[24] & b[119])^(a[23] & b[120])^(a[22] & b[121])^(a[21] & b[122])^(a[20] & b[123])^(a[19] & b[124])^(a[18] & b[125])^(a[17] & b[126])^(a[16] & b[127])^(a[15] & b[128])^(a[14] & b[129])^(a[13] & b[130])^(a[12] & b[131])^(a[11] & b[132])^(a[10] & b[133])^(a[9] & b[134])^(a[8] & b[135])^(a[7] & b[136])^(a[6] & b[137])^(a[5] & b[138])^(a[4] & b[139])^(a[3] & b[140])^(a[2] & b[141])^(a[1] & b[142])^(a[0] & b[143]);
assign y[144] = (a[144] & b[0])^(a[143] & b[1])^(a[142] & b[2])^(a[141] & b[3])^(a[140] & b[4])^(a[139] & b[5])^(a[138] & b[6])^(a[137] & b[7])^(a[136] & b[8])^(a[135] & b[9])^(a[134] & b[10])^(a[133] & b[11])^(a[132] & b[12])^(a[131] & b[13])^(a[130] & b[14])^(a[129] & b[15])^(a[128] & b[16])^(a[127] & b[17])^(a[126] & b[18])^(a[125] & b[19])^(a[124] & b[20])^(a[123] & b[21])^(a[122] & b[22])^(a[121] & b[23])^(a[120] & b[24])^(a[119] & b[25])^(a[118] & b[26])^(a[117] & b[27])^(a[116] & b[28])^(a[115] & b[29])^(a[114] & b[30])^(a[113] & b[31])^(a[112] & b[32])^(a[111] & b[33])^(a[110] & b[34])^(a[109] & b[35])^(a[108] & b[36])^(a[107] & b[37])^(a[106] & b[38])^(a[105] & b[39])^(a[104] & b[40])^(a[103] & b[41])^(a[102] & b[42])^(a[101] & b[43])^(a[100] & b[44])^(a[99] & b[45])^(a[98] & b[46])^(a[97] & b[47])^(a[96] & b[48])^(a[95] & b[49])^(a[94] & b[50])^(a[93] & b[51])^(a[92] & b[52])^(a[91] & b[53])^(a[90] & b[54])^(a[89] & b[55])^(a[88] & b[56])^(a[87] & b[57])^(a[86] & b[58])^(a[85] & b[59])^(a[84] & b[60])^(a[83] & b[61])^(a[82] & b[62])^(a[81] & b[63])^(a[80] & b[64])^(a[79] & b[65])^(a[78] & b[66])^(a[77] & b[67])^(a[76] & b[68])^(a[75] & b[69])^(a[74] & b[70])^(a[73] & b[71])^(a[72] & b[72])^(a[71] & b[73])^(a[70] & b[74])^(a[69] & b[75])^(a[68] & b[76])^(a[67] & b[77])^(a[66] & b[78])^(a[65] & b[79])^(a[64] & b[80])^(a[63] & b[81])^(a[62] & b[82])^(a[61] & b[83])^(a[60] & b[84])^(a[59] & b[85])^(a[58] & b[86])^(a[57] & b[87])^(a[56] & b[88])^(a[55] & b[89])^(a[54] & b[90])^(a[53] & b[91])^(a[52] & b[92])^(a[51] & b[93])^(a[50] & b[94])^(a[49] & b[95])^(a[48] & b[96])^(a[47] & b[97])^(a[46] & b[98])^(a[45] & b[99])^(a[44] & b[100])^(a[43] & b[101])^(a[42] & b[102])^(a[41] & b[103])^(a[40] & b[104])^(a[39] & b[105])^(a[38] & b[106])^(a[37] & b[107])^(a[36] & b[108])^(a[35] & b[109])^(a[34] & b[110])^(a[33] & b[111])^(a[32] & b[112])^(a[31] & b[113])^(a[30] & b[114])^(a[29] & b[115])^(a[28] & b[116])^(a[27] & b[117])^(a[26] & b[118])^(a[25] & b[119])^(a[24] & b[120])^(a[23] & b[121])^(a[22] & b[122])^(a[21] & b[123])^(a[20] & b[124])^(a[19] & b[125])^(a[18] & b[126])^(a[17] & b[127])^(a[16] & b[128])^(a[15] & b[129])^(a[14] & b[130])^(a[13] & b[131])^(a[12] & b[132])^(a[11] & b[133])^(a[10] & b[134])^(a[9] & b[135])^(a[8] & b[136])^(a[7] & b[137])^(a[6] & b[138])^(a[5] & b[139])^(a[4] & b[140])^(a[3] & b[141])^(a[2] & b[142])^(a[1] & b[143])^(a[0] & b[144]);
assign y[145] = (a[145] & b[0])^(a[144] & b[1])^(a[143] & b[2])^(a[142] & b[3])^(a[141] & b[4])^(a[140] & b[5])^(a[139] & b[6])^(a[138] & b[7])^(a[137] & b[8])^(a[136] & b[9])^(a[135] & b[10])^(a[134] & b[11])^(a[133] & b[12])^(a[132] & b[13])^(a[131] & b[14])^(a[130] & b[15])^(a[129] & b[16])^(a[128] & b[17])^(a[127] & b[18])^(a[126] & b[19])^(a[125] & b[20])^(a[124] & b[21])^(a[123] & b[22])^(a[122] & b[23])^(a[121] & b[24])^(a[120] & b[25])^(a[119] & b[26])^(a[118] & b[27])^(a[117] & b[28])^(a[116] & b[29])^(a[115] & b[30])^(a[114] & b[31])^(a[113] & b[32])^(a[112] & b[33])^(a[111] & b[34])^(a[110] & b[35])^(a[109] & b[36])^(a[108] & b[37])^(a[107] & b[38])^(a[106] & b[39])^(a[105] & b[40])^(a[104] & b[41])^(a[103] & b[42])^(a[102] & b[43])^(a[101] & b[44])^(a[100] & b[45])^(a[99] & b[46])^(a[98] & b[47])^(a[97] & b[48])^(a[96] & b[49])^(a[95] & b[50])^(a[94] & b[51])^(a[93] & b[52])^(a[92] & b[53])^(a[91] & b[54])^(a[90] & b[55])^(a[89] & b[56])^(a[88] & b[57])^(a[87] & b[58])^(a[86] & b[59])^(a[85] & b[60])^(a[84] & b[61])^(a[83] & b[62])^(a[82] & b[63])^(a[81] & b[64])^(a[80] & b[65])^(a[79] & b[66])^(a[78] & b[67])^(a[77] & b[68])^(a[76] & b[69])^(a[75] & b[70])^(a[74] & b[71])^(a[73] & b[72])^(a[72] & b[73])^(a[71] & b[74])^(a[70] & b[75])^(a[69] & b[76])^(a[68] & b[77])^(a[67] & b[78])^(a[66] & b[79])^(a[65] & b[80])^(a[64] & b[81])^(a[63] & b[82])^(a[62] & b[83])^(a[61] & b[84])^(a[60] & b[85])^(a[59] & b[86])^(a[58] & b[87])^(a[57] & b[88])^(a[56] & b[89])^(a[55] & b[90])^(a[54] & b[91])^(a[53] & b[92])^(a[52] & b[93])^(a[51] & b[94])^(a[50] & b[95])^(a[49] & b[96])^(a[48] & b[97])^(a[47] & b[98])^(a[46] & b[99])^(a[45] & b[100])^(a[44] & b[101])^(a[43] & b[102])^(a[42] & b[103])^(a[41] & b[104])^(a[40] & b[105])^(a[39] & b[106])^(a[38] & b[107])^(a[37] & b[108])^(a[36] & b[109])^(a[35] & b[110])^(a[34] & b[111])^(a[33] & b[112])^(a[32] & b[113])^(a[31] & b[114])^(a[30] & b[115])^(a[29] & b[116])^(a[28] & b[117])^(a[27] & b[118])^(a[26] & b[119])^(a[25] & b[120])^(a[24] & b[121])^(a[23] & b[122])^(a[22] & b[123])^(a[21] & b[124])^(a[20] & b[125])^(a[19] & b[126])^(a[18] & b[127])^(a[17] & b[128])^(a[16] & b[129])^(a[15] & b[130])^(a[14] & b[131])^(a[13] & b[132])^(a[12] & b[133])^(a[11] & b[134])^(a[10] & b[135])^(a[9] & b[136])^(a[8] & b[137])^(a[7] & b[138])^(a[6] & b[139])^(a[5] & b[140])^(a[4] & b[141])^(a[3] & b[142])^(a[2] & b[143])^(a[1] & b[144])^(a[0] & b[145]);
assign y[146] = (a[146] & b[0])^(a[145] & b[1])^(a[144] & b[2])^(a[143] & b[3])^(a[142] & b[4])^(a[141] & b[5])^(a[140] & b[6])^(a[139] & b[7])^(a[138] & b[8])^(a[137] & b[9])^(a[136] & b[10])^(a[135] & b[11])^(a[134] & b[12])^(a[133] & b[13])^(a[132] & b[14])^(a[131] & b[15])^(a[130] & b[16])^(a[129] & b[17])^(a[128] & b[18])^(a[127] & b[19])^(a[126] & b[20])^(a[125] & b[21])^(a[124] & b[22])^(a[123] & b[23])^(a[122] & b[24])^(a[121] & b[25])^(a[120] & b[26])^(a[119] & b[27])^(a[118] & b[28])^(a[117] & b[29])^(a[116] & b[30])^(a[115] & b[31])^(a[114] & b[32])^(a[113] & b[33])^(a[112] & b[34])^(a[111] & b[35])^(a[110] & b[36])^(a[109] & b[37])^(a[108] & b[38])^(a[107] & b[39])^(a[106] & b[40])^(a[105] & b[41])^(a[104] & b[42])^(a[103] & b[43])^(a[102] & b[44])^(a[101] & b[45])^(a[100] & b[46])^(a[99] & b[47])^(a[98] & b[48])^(a[97] & b[49])^(a[96] & b[50])^(a[95] & b[51])^(a[94] & b[52])^(a[93] & b[53])^(a[92] & b[54])^(a[91] & b[55])^(a[90] & b[56])^(a[89] & b[57])^(a[88] & b[58])^(a[87] & b[59])^(a[86] & b[60])^(a[85] & b[61])^(a[84] & b[62])^(a[83] & b[63])^(a[82] & b[64])^(a[81] & b[65])^(a[80] & b[66])^(a[79] & b[67])^(a[78] & b[68])^(a[77] & b[69])^(a[76] & b[70])^(a[75] & b[71])^(a[74] & b[72])^(a[73] & b[73])^(a[72] & b[74])^(a[71] & b[75])^(a[70] & b[76])^(a[69] & b[77])^(a[68] & b[78])^(a[67] & b[79])^(a[66] & b[80])^(a[65] & b[81])^(a[64] & b[82])^(a[63] & b[83])^(a[62] & b[84])^(a[61] & b[85])^(a[60] & b[86])^(a[59] & b[87])^(a[58] & b[88])^(a[57] & b[89])^(a[56] & b[90])^(a[55] & b[91])^(a[54] & b[92])^(a[53] & b[93])^(a[52] & b[94])^(a[51] & b[95])^(a[50] & b[96])^(a[49] & b[97])^(a[48] & b[98])^(a[47] & b[99])^(a[46] & b[100])^(a[45] & b[101])^(a[44] & b[102])^(a[43] & b[103])^(a[42] & b[104])^(a[41] & b[105])^(a[40] & b[106])^(a[39] & b[107])^(a[38] & b[108])^(a[37] & b[109])^(a[36] & b[110])^(a[35] & b[111])^(a[34] & b[112])^(a[33] & b[113])^(a[32] & b[114])^(a[31] & b[115])^(a[30] & b[116])^(a[29] & b[117])^(a[28] & b[118])^(a[27] & b[119])^(a[26] & b[120])^(a[25] & b[121])^(a[24] & b[122])^(a[23] & b[123])^(a[22] & b[124])^(a[21] & b[125])^(a[20] & b[126])^(a[19] & b[127])^(a[18] & b[128])^(a[17] & b[129])^(a[16] & b[130])^(a[15] & b[131])^(a[14] & b[132])^(a[13] & b[133])^(a[12] & b[134])^(a[11] & b[135])^(a[10] & b[136])^(a[9] & b[137])^(a[8] & b[138])^(a[7] & b[139])^(a[6] & b[140])^(a[5] & b[141])^(a[4] & b[142])^(a[3] & b[143])^(a[2] & b[144])^(a[1] & b[145])^(a[0] & b[146]);
assign y[147] = (a[147] & b[0])^(a[146] & b[1])^(a[145] & b[2])^(a[144] & b[3])^(a[143] & b[4])^(a[142] & b[5])^(a[141] & b[6])^(a[140] & b[7])^(a[139] & b[8])^(a[138] & b[9])^(a[137] & b[10])^(a[136] & b[11])^(a[135] & b[12])^(a[134] & b[13])^(a[133] & b[14])^(a[132] & b[15])^(a[131] & b[16])^(a[130] & b[17])^(a[129] & b[18])^(a[128] & b[19])^(a[127] & b[20])^(a[126] & b[21])^(a[125] & b[22])^(a[124] & b[23])^(a[123] & b[24])^(a[122] & b[25])^(a[121] & b[26])^(a[120] & b[27])^(a[119] & b[28])^(a[118] & b[29])^(a[117] & b[30])^(a[116] & b[31])^(a[115] & b[32])^(a[114] & b[33])^(a[113] & b[34])^(a[112] & b[35])^(a[111] & b[36])^(a[110] & b[37])^(a[109] & b[38])^(a[108] & b[39])^(a[107] & b[40])^(a[106] & b[41])^(a[105] & b[42])^(a[104] & b[43])^(a[103] & b[44])^(a[102] & b[45])^(a[101] & b[46])^(a[100] & b[47])^(a[99] & b[48])^(a[98] & b[49])^(a[97] & b[50])^(a[96] & b[51])^(a[95] & b[52])^(a[94] & b[53])^(a[93] & b[54])^(a[92] & b[55])^(a[91] & b[56])^(a[90] & b[57])^(a[89] & b[58])^(a[88] & b[59])^(a[87] & b[60])^(a[86] & b[61])^(a[85] & b[62])^(a[84] & b[63])^(a[83] & b[64])^(a[82] & b[65])^(a[81] & b[66])^(a[80] & b[67])^(a[79] & b[68])^(a[78] & b[69])^(a[77] & b[70])^(a[76] & b[71])^(a[75] & b[72])^(a[74] & b[73])^(a[73] & b[74])^(a[72] & b[75])^(a[71] & b[76])^(a[70] & b[77])^(a[69] & b[78])^(a[68] & b[79])^(a[67] & b[80])^(a[66] & b[81])^(a[65] & b[82])^(a[64] & b[83])^(a[63] & b[84])^(a[62] & b[85])^(a[61] & b[86])^(a[60] & b[87])^(a[59] & b[88])^(a[58] & b[89])^(a[57] & b[90])^(a[56] & b[91])^(a[55] & b[92])^(a[54] & b[93])^(a[53] & b[94])^(a[52] & b[95])^(a[51] & b[96])^(a[50] & b[97])^(a[49] & b[98])^(a[48] & b[99])^(a[47] & b[100])^(a[46] & b[101])^(a[45] & b[102])^(a[44] & b[103])^(a[43] & b[104])^(a[42] & b[105])^(a[41] & b[106])^(a[40] & b[107])^(a[39] & b[108])^(a[38] & b[109])^(a[37] & b[110])^(a[36] & b[111])^(a[35] & b[112])^(a[34] & b[113])^(a[33] & b[114])^(a[32] & b[115])^(a[31] & b[116])^(a[30] & b[117])^(a[29] & b[118])^(a[28] & b[119])^(a[27] & b[120])^(a[26] & b[121])^(a[25] & b[122])^(a[24] & b[123])^(a[23] & b[124])^(a[22] & b[125])^(a[21] & b[126])^(a[20] & b[127])^(a[19] & b[128])^(a[18] & b[129])^(a[17] & b[130])^(a[16] & b[131])^(a[15] & b[132])^(a[14] & b[133])^(a[13] & b[134])^(a[12] & b[135])^(a[11] & b[136])^(a[10] & b[137])^(a[9] & b[138])^(a[8] & b[139])^(a[7] & b[140])^(a[6] & b[141])^(a[5] & b[142])^(a[4] & b[143])^(a[3] & b[144])^(a[2] & b[145])^(a[1] & b[146])^(a[0] & b[147]);
assign y[148] = (a[148] & b[0])^(a[147] & b[1])^(a[146] & b[2])^(a[145] & b[3])^(a[144] & b[4])^(a[143] & b[5])^(a[142] & b[6])^(a[141] & b[7])^(a[140] & b[8])^(a[139] & b[9])^(a[138] & b[10])^(a[137] & b[11])^(a[136] & b[12])^(a[135] & b[13])^(a[134] & b[14])^(a[133] & b[15])^(a[132] & b[16])^(a[131] & b[17])^(a[130] & b[18])^(a[129] & b[19])^(a[128] & b[20])^(a[127] & b[21])^(a[126] & b[22])^(a[125] & b[23])^(a[124] & b[24])^(a[123] & b[25])^(a[122] & b[26])^(a[121] & b[27])^(a[120] & b[28])^(a[119] & b[29])^(a[118] & b[30])^(a[117] & b[31])^(a[116] & b[32])^(a[115] & b[33])^(a[114] & b[34])^(a[113] & b[35])^(a[112] & b[36])^(a[111] & b[37])^(a[110] & b[38])^(a[109] & b[39])^(a[108] & b[40])^(a[107] & b[41])^(a[106] & b[42])^(a[105] & b[43])^(a[104] & b[44])^(a[103] & b[45])^(a[102] & b[46])^(a[101] & b[47])^(a[100] & b[48])^(a[99] & b[49])^(a[98] & b[50])^(a[97] & b[51])^(a[96] & b[52])^(a[95] & b[53])^(a[94] & b[54])^(a[93] & b[55])^(a[92] & b[56])^(a[91] & b[57])^(a[90] & b[58])^(a[89] & b[59])^(a[88] & b[60])^(a[87] & b[61])^(a[86] & b[62])^(a[85] & b[63])^(a[84] & b[64])^(a[83] & b[65])^(a[82] & b[66])^(a[81] & b[67])^(a[80] & b[68])^(a[79] & b[69])^(a[78] & b[70])^(a[77] & b[71])^(a[76] & b[72])^(a[75] & b[73])^(a[74] & b[74])^(a[73] & b[75])^(a[72] & b[76])^(a[71] & b[77])^(a[70] & b[78])^(a[69] & b[79])^(a[68] & b[80])^(a[67] & b[81])^(a[66] & b[82])^(a[65] & b[83])^(a[64] & b[84])^(a[63] & b[85])^(a[62] & b[86])^(a[61] & b[87])^(a[60] & b[88])^(a[59] & b[89])^(a[58] & b[90])^(a[57] & b[91])^(a[56] & b[92])^(a[55] & b[93])^(a[54] & b[94])^(a[53] & b[95])^(a[52] & b[96])^(a[51] & b[97])^(a[50] & b[98])^(a[49] & b[99])^(a[48] & b[100])^(a[47] & b[101])^(a[46] & b[102])^(a[45] & b[103])^(a[44] & b[104])^(a[43] & b[105])^(a[42] & b[106])^(a[41] & b[107])^(a[40] & b[108])^(a[39] & b[109])^(a[38] & b[110])^(a[37] & b[111])^(a[36] & b[112])^(a[35] & b[113])^(a[34] & b[114])^(a[33] & b[115])^(a[32] & b[116])^(a[31] & b[117])^(a[30] & b[118])^(a[29] & b[119])^(a[28] & b[120])^(a[27] & b[121])^(a[26] & b[122])^(a[25] & b[123])^(a[24] & b[124])^(a[23] & b[125])^(a[22] & b[126])^(a[21] & b[127])^(a[20] & b[128])^(a[19] & b[129])^(a[18] & b[130])^(a[17] & b[131])^(a[16] & b[132])^(a[15] & b[133])^(a[14] & b[134])^(a[13] & b[135])^(a[12] & b[136])^(a[11] & b[137])^(a[10] & b[138])^(a[9] & b[139])^(a[8] & b[140])^(a[7] & b[141])^(a[6] & b[142])^(a[5] & b[143])^(a[4] & b[144])^(a[3] & b[145])^(a[2] & b[146])^(a[1] & b[147])^(a[0] & b[148]);
assign y[149] = (a[149] & b[0])^(a[148] & b[1])^(a[147] & b[2])^(a[146] & b[3])^(a[145] & b[4])^(a[144] & b[5])^(a[143] & b[6])^(a[142] & b[7])^(a[141] & b[8])^(a[140] & b[9])^(a[139] & b[10])^(a[138] & b[11])^(a[137] & b[12])^(a[136] & b[13])^(a[135] & b[14])^(a[134] & b[15])^(a[133] & b[16])^(a[132] & b[17])^(a[131] & b[18])^(a[130] & b[19])^(a[129] & b[20])^(a[128] & b[21])^(a[127] & b[22])^(a[126] & b[23])^(a[125] & b[24])^(a[124] & b[25])^(a[123] & b[26])^(a[122] & b[27])^(a[121] & b[28])^(a[120] & b[29])^(a[119] & b[30])^(a[118] & b[31])^(a[117] & b[32])^(a[116] & b[33])^(a[115] & b[34])^(a[114] & b[35])^(a[113] & b[36])^(a[112] & b[37])^(a[111] & b[38])^(a[110] & b[39])^(a[109] & b[40])^(a[108] & b[41])^(a[107] & b[42])^(a[106] & b[43])^(a[105] & b[44])^(a[104] & b[45])^(a[103] & b[46])^(a[102] & b[47])^(a[101] & b[48])^(a[100] & b[49])^(a[99] & b[50])^(a[98] & b[51])^(a[97] & b[52])^(a[96] & b[53])^(a[95] & b[54])^(a[94] & b[55])^(a[93] & b[56])^(a[92] & b[57])^(a[91] & b[58])^(a[90] & b[59])^(a[89] & b[60])^(a[88] & b[61])^(a[87] & b[62])^(a[86] & b[63])^(a[85] & b[64])^(a[84] & b[65])^(a[83] & b[66])^(a[82] & b[67])^(a[81] & b[68])^(a[80] & b[69])^(a[79] & b[70])^(a[78] & b[71])^(a[77] & b[72])^(a[76] & b[73])^(a[75] & b[74])^(a[74] & b[75])^(a[73] & b[76])^(a[72] & b[77])^(a[71] & b[78])^(a[70] & b[79])^(a[69] & b[80])^(a[68] & b[81])^(a[67] & b[82])^(a[66] & b[83])^(a[65] & b[84])^(a[64] & b[85])^(a[63] & b[86])^(a[62] & b[87])^(a[61] & b[88])^(a[60] & b[89])^(a[59] & b[90])^(a[58] & b[91])^(a[57] & b[92])^(a[56] & b[93])^(a[55] & b[94])^(a[54] & b[95])^(a[53] & b[96])^(a[52] & b[97])^(a[51] & b[98])^(a[50] & b[99])^(a[49] & b[100])^(a[48] & b[101])^(a[47] & b[102])^(a[46] & b[103])^(a[45] & b[104])^(a[44] & b[105])^(a[43] & b[106])^(a[42] & b[107])^(a[41] & b[108])^(a[40] & b[109])^(a[39] & b[110])^(a[38] & b[111])^(a[37] & b[112])^(a[36] & b[113])^(a[35] & b[114])^(a[34] & b[115])^(a[33] & b[116])^(a[32] & b[117])^(a[31] & b[118])^(a[30] & b[119])^(a[29] & b[120])^(a[28] & b[121])^(a[27] & b[122])^(a[26] & b[123])^(a[25] & b[124])^(a[24] & b[125])^(a[23] & b[126])^(a[22] & b[127])^(a[21] & b[128])^(a[20] & b[129])^(a[19] & b[130])^(a[18] & b[131])^(a[17] & b[132])^(a[16] & b[133])^(a[15] & b[134])^(a[14] & b[135])^(a[13] & b[136])^(a[12] & b[137])^(a[11] & b[138])^(a[10] & b[139])^(a[9] & b[140])^(a[8] & b[141])^(a[7] & b[142])^(a[6] & b[143])^(a[5] & b[144])^(a[4] & b[145])^(a[3] & b[146])^(a[2] & b[147])^(a[1] & b[148])^(a[0] & b[149]);
assign y[150] = (a[150] & b[0])^(a[149] & b[1])^(a[148] & b[2])^(a[147] & b[3])^(a[146] & b[4])^(a[145] & b[5])^(a[144] & b[6])^(a[143] & b[7])^(a[142] & b[8])^(a[141] & b[9])^(a[140] & b[10])^(a[139] & b[11])^(a[138] & b[12])^(a[137] & b[13])^(a[136] & b[14])^(a[135] & b[15])^(a[134] & b[16])^(a[133] & b[17])^(a[132] & b[18])^(a[131] & b[19])^(a[130] & b[20])^(a[129] & b[21])^(a[128] & b[22])^(a[127] & b[23])^(a[126] & b[24])^(a[125] & b[25])^(a[124] & b[26])^(a[123] & b[27])^(a[122] & b[28])^(a[121] & b[29])^(a[120] & b[30])^(a[119] & b[31])^(a[118] & b[32])^(a[117] & b[33])^(a[116] & b[34])^(a[115] & b[35])^(a[114] & b[36])^(a[113] & b[37])^(a[112] & b[38])^(a[111] & b[39])^(a[110] & b[40])^(a[109] & b[41])^(a[108] & b[42])^(a[107] & b[43])^(a[106] & b[44])^(a[105] & b[45])^(a[104] & b[46])^(a[103] & b[47])^(a[102] & b[48])^(a[101] & b[49])^(a[100] & b[50])^(a[99] & b[51])^(a[98] & b[52])^(a[97] & b[53])^(a[96] & b[54])^(a[95] & b[55])^(a[94] & b[56])^(a[93] & b[57])^(a[92] & b[58])^(a[91] & b[59])^(a[90] & b[60])^(a[89] & b[61])^(a[88] & b[62])^(a[87] & b[63])^(a[86] & b[64])^(a[85] & b[65])^(a[84] & b[66])^(a[83] & b[67])^(a[82] & b[68])^(a[81] & b[69])^(a[80] & b[70])^(a[79] & b[71])^(a[78] & b[72])^(a[77] & b[73])^(a[76] & b[74])^(a[75] & b[75])^(a[74] & b[76])^(a[73] & b[77])^(a[72] & b[78])^(a[71] & b[79])^(a[70] & b[80])^(a[69] & b[81])^(a[68] & b[82])^(a[67] & b[83])^(a[66] & b[84])^(a[65] & b[85])^(a[64] & b[86])^(a[63] & b[87])^(a[62] & b[88])^(a[61] & b[89])^(a[60] & b[90])^(a[59] & b[91])^(a[58] & b[92])^(a[57] & b[93])^(a[56] & b[94])^(a[55] & b[95])^(a[54] & b[96])^(a[53] & b[97])^(a[52] & b[98])^(a[51] & b[99])^(a[50] & b[100])^(a[49] & b[101])^(a[48] & b[102])^(a[47] & b[103])^(a[46] & b[104])^(a[45] & b[105])^(a[44] & b[106])^(a[43] & b[107])^(a[42] & b[108])^(a[41] & b[109])^(a[40] & b[110])^(a[39] & b[111])^(a[38] & b[112])^(a[37] & b[113])^(a[36] & b[114])^(a[35] & b[115])^(a[34] & b[116])^(a[33] & b[117])^(a[32] & b[118])^(a[31] & b[119])^(a[30] & b[120])^(a[29] & b[121])^(a[28] & b[122])^(a[27] & b[123])^(a[26] & b[124])^(a[25] & b[125])^(a[24] & b[126])^(a[23] & b[127])^(a[22] & b[128])^(a[21] & b[129])^(a[20] & b[130])^(a[19] & b[131])^(a[18] & b[132])^(a[17] & b[133])^(a[16] & b[134])^(a[15] & b[135])^(a[14] & b[136])^(a[13] & b[137])^(a[12] & b[138])^(a[11] & b[139])^(a[10] & b[140])^(a[9] & b[141])^(a[8] & b[142])^(a[7] & b[143])^(a[6] & b[144])^(a[5] & b[145])^(a[4] & b[146])^(a[3] & b[147])^(a[2] & b[148])^(a[1] & b[149])^(a[0] & b[150]);
assign y[151] = (a[151] & b[0])^(a[150] & b[1])^(a[149] & b[2])^(a[148] & b[3])^(a[147] & b[4])^(a[146] & b[5])^(a[145] & b[6])^(a[144] & b[7])^(a[143] & b[8])^(a[142] & b[9])^(a[141] & b[10])^(a[140] & b[11])^(a[139] & b[12])^(a[138] & b[13])^(a[137] & b[14])^(a[136] & b[15])^(a[135] & b[16])^(a[134] & b[17])^(a[133] & b[18])^(a[132] & b[19])^(a[131] & b[20])^(a[130] & b[21])^(a[129] & b[22])^(a[128] & b[23])^(a[127] & b[24])^(a[126] & b[25])^(a[125] & b[26])^(a[124] & b[27])^(a[123] & b[28])^(a[122] & b[29])^(a[121] & b[30])^(a[120] & b[31])^(a[119] & b[32])^(a[118] & b[33])^(a[117] & b[34])^(a[116] & b[35])^(a[115] & b[36])^(a[114] & b[37])^(a[113] & b[38])^(a[112] & b[39])^(a[111] & b[40])^(a[110] & b[41])^(a[109] & b[42])^(a[108] & b[43])^(a[107] & b[44])^(a[106] & b[45])^(a[105] & b[46])^(a[104] & b[47])^(a[103] & b[48])^(a[102] & b[49])^(a[101] & b[50])^(a[100] & b[51])^(a[99] & b[52])^(a[98] & b[53])^(a[97] & b[54])^(a[96] & b[55])^(a[95] & b[56])^(a[94] & b[57])^(a[93] & b[58])^(a[92] & b[59])^(a[91] & b[60])^(a[90] & b[61])^(a[89] & b[62])^(a[88] & b[63])^(a[87] & b[64])^(a[86] & b[65])^(a[85] & b[66])^(a[84] & b[67])^(a[83] & b[68])^(a[82] & b[69])^(a[81] & b[70])^(a[80] & b[71])^(a[79] & b[72])^(a[78] & b[73])^(a[77] & b[74])^(a[76] & b[75])^(a[75] & b[76])^(a[74] & b[77])^(a[73] & b[78])^(a[72] & b[79])^(a[71] & b[80])^(a[70] & b[81])^(a[69] & b[82])^(a[68] & b[83])^(a[67] & b[84])^(a[66] & b[85])^(a[65] & b[86])^(a[64] & b[87])^(a[63] & b[88])^(a[62] & b[89])^(a[61] & b[90])^(a[60] & b[91])^(a[59] & b[92])^(a[58] & b[93])^(a[57] & b[94])^(a[56] & b[95])^(a[55] & b[96])^(a[54] & b[97])^(a[53] & b[98])^(a[52] & b[99])^(a[51] & b[100])^(a[50] & b[101])^(a[49] & b[102])^(a[48] & b[103])^(a[47] & b[104])^(a[46] & b[105])^(a[45] & b[106])^(a[44] & b[107])^(a[43] & b[108])^(a[42] & b[109])^(a[41] & b[110])^(a[40] & b[111])^(a[39] & b[112])^(a[38] & b[113])^(a[37] & b[114])^(a[36] & b[115])^(a[35] & b[116])^(a[34] & b[117])^(a[33] & b[118])^(a[32] & b[119])^(a[31] & b[120])^(a[30] & b[121])^(a[29] & b[122])^(a[28] & b[123])^(a[27] & b[124])^(a[26] & b[125])^(a[25] & b[126])^(a[24] & b[127])^(a[23] & b[128])^(a[22] & b[129])^(a[21] & b[130])^(a[20] & b[131])^(a[19] & b[132])^(a[18] & b[133])^(a[17] & b[134])^(a[16] & b[135])^(a[15] & b[136])^(a[14] & b[137])^(a[13] & b[138])^(a[12] & b[139])^(a[11] & b[140])^(a[10] & b[141])^(a[9] & b[142])^(a[8] & b[143])^(a[7] & b[144])^(a[6] & b[145])^(a[5] & b[146])^(a[4] & b[147])^(a[3] & b[148])^(a[2] & b[149])^(a[1] & b[150])^(a[0] & b[151]);
assign y[152] = (a[152] & b[0])^(a[151] & b[1])^(a[150] & b[2])^(a[149] & b[3])^(a[148] & b[4])^(a[147] & b[5])^(a[146] & b[6])^(a[145] & b[7])^(a[144] & b[8])^(a[143] & b[9])^(a[142] & b[10])^(a[141] & b[11])^(a[140] & b[12])^(a[139] & b[13])^(a[138] & b[14])^(a[137] & b[15])^(a[136] & b[16])^(a[135] & b[17])^(a[134] & b[18])^(a[133] & b[19])^(a[132] & b[20])^(a[131] & b[21])^(a[130] & b[22])^(a[129] & b[23])^(a[128] & b[24])^(a[127] & b[25])^(a[126] & b[26])^(a[125] & b[27])^(a[124] & b[28])^(a[123] & b[29])^(a[122] & b[30])^(a[121] & b[31])^(a[120] & b[32])^(a[119] & b[33])^(a[118] & b[34])^(a[117] & b[35])^(a[116] & b[36])^(a[115] & b[37])^(a[114] & b[38])^(a[113] & b[39])^(a[112] & b[40])^(a[111] & b[41])^(a[110] & b[42])^(a[109] & b[43])^(a[108] & b[44])^(a[107] & b[45])^(a[106] & b[46])^(a[105] & b[47])^(a[104] & b[48])^(a[103] & b[49])^(a[102] & b[50])^(a[101] & b[51])^(a[100] & b[52])^(a[99] & b[53])^(a[98] & b[54])^(a[97] & b[55])^(a[96] & b[56])^(a[95] & b[57])^(a[94] & b[58])^(a[93] & b[59])^(a[92] & b[60])^(a[91] & b[61])^(a[90] & b[62])^(a[89] & b[63])^(a[88] & b[64])^(a[87] & b[65])^(a[86] & b[66])^(a[85] & b[67])^(a[84] & b[68])^(a[83] & b[69])^(a[82] & b[70])^(a[81] & b[71])^(a[80] & b[72])^(a[79] & b[73])^(a[78] & b[74])^(a[77] & b[75])^(a[76] & b[76])^(a[75] & b[77])^(a[74] & b[78])^(a[73] & b[79])^(a[72] & b[80])^(a[71] & b[81])^(a[70] & b[82])^(a[69] & b[83])^(a[68] & b[84])^(a[67] & b[85])^(a[66] & b[86])^(a[65] & b[87])^(a[64] & b[88])^(a[63] & b[89])^(a[62] & b[90])^(a[61] & b[91])^(a[60] & b[92])^(a[59] & b[93])^(a[58] & b[94])^(a[57] & b[95])^(a[56] & b[96])^(a[55] & b[97])^(a[54] & b[98])^(a[53] & b[99])^(a[52] & b[100])^(a[51] & b[101])^(a[50] & b[102])^(a[49] & b[103])^(a[48] & b[104])^(a[47] & b[105])^(a[46] & b[106])^(a[45] & b[107])^(a[44] & b[108])^(a[43] & b[109])^(a[42] & b[110])^(a[41] & b[111])^(a[40] & b[112])^(a[39] & b[113])^(a[38] & b[114])^(a[37] & b[115])^(a[36] & b[116])^(a[35] & b[117])^(a[34] & b[118])^(a[33] & b[119])^(a[32] & b[120])^(a[31] & b[121])^(a[30] & b[122])^(a[29] & b[123])^(a[28] & b[124])^(a[27] & b[125])^(a[26] & b[126])^(a[25] & b[127])^(a[24] & b[128])^(a[23] & b[129])^(a[22] & b[130])^(a[21] & b[131])^(a[20] & b[132])^(a[19] & b[133])^(a[18] & b[134])^(a[17] & b[135])^(a[16] & b[136])^(a[15] & b[137])^(a[14] & b[138])^(a[13] & b[139])^(a[12] & b[140])^(a[11] & b[141])^(a[10] & b[142])^(a[9] & b[143])^(a[8] & b[144])^(a[7] & b[145])^(a[6] & b[146])^(a[5] & b[147])^(a[4] & b[148])^(a[3] & b[149])^(a[2] & b[150])^(a[1] & b[151])^(a[0] & b[152]);
assign y[153] = (a[153] & b[0])^(a[152] & b[1])^(a[151] & b[2])^(a[150] & b[3])^(a[149] & b[4])^(a[148] & b[5])^(a[147] & b[6])^(a[146] & b[7])^(a[145] & b[8])^(a[144] & b[9])^(a[143] & b[10])^(a[142] & b[11])^(a[141] & b[12])^(a[140] & b[13])^(a[139] & b[14])^(a[138] & b[15])^(a[137] & b[16])^(a[136] & b[17])^(a[135] & b[18])^(a[134] & b[19])^(a[133] & b[20])^(a[132] & b[21])^(a[131] & b[22])^(a[130] & b[23])^(a[129] & b[24])^(a[128] & b[25])^(a[127] & b[26])^(a[126] & b[27])^(a[125] & b[28])^(a[124] & b[29])^(a[123] & b[30])^(a[122] & b[31])^(a[121] & b[32])^(a[120] & b[33])^(a[119] & b[34])^(a[118] & b[35])^(a[117] & b[36])^(a[116] & b[37])^(a[115] & b[38])^(a[114] & b[39])^(a[113] & b[40])^(a[112] & b[41])^(a[111] & b[42])^(a[110] & b[43])^(a[109] & b[44])^(a[108] & b[45])^(a[107] & b[46])^(a[106] & b[47])^(a[105] & b[48])^(a[104] & b[49])^(a[103] & b[50])^(a[102] & b[51])^(a[101] & b[52])^(a[100] & b[53])^(a[99] & b[54])^(a[98] & b[55])^(a[97] & b[56])^(a[96] & b[57])^(a[95] & b[58])^(a[94] & b[59])^(a[93] & b[60])^(a[92] & b[61])^(a[91] & b[62])^(a[90] & b[63])^(a[89] & b[64])^(a[88] & b[65])^(a[87] & b[66])^(a[86] & b[67])^(a[85] & b[68])^(a[84] & b[69])^(a[83] & b[70])^(a[82] & b[71])^(a[81] & b[72])^(a[80] & b[73])^(a[79] & b[74])^(a[78] & b[75])^(a[77] & b[76])^(a[76] & b[77])^(a[75] & b[78])^(a[74] & b[79])^(a[73] & b[80])^(a[72] & b[81])^(a[71] & b[82])^(a[70] & b[83])^(a[69] & b[84])^(a[68] & b[85])^(a[67] & b[86])^(a[66] & b[87])^(a[65] & b[88])^(a[64] & b[89])^(a[63] & b[90])^(a[62] & b[91])^(a[61] & b[92])^(a[60] & b[93])^(a[59] & b[94])^(a[58] & b[95])^(a[57] & b[96])^(a[56] & b[97])^(a[55] & b[98])^(a[54] & b[99])^(a[53] & b[100])^(a[52] & b[101])^(a[51] & b[102])^(a[50] & b[103])^(a[49] & b[104])^(a[48] & b[105])^(a[47] & b[106])^(a[46] & b[107])^(a[45] & b[108])^(a[44] & b[109])^(a[43] & b[110])^(a[42] & b[111])^(a[41] & b[112])^(a[40] & b[113])^(a[39] & b[114])^(a[38] & b[115])^(a[37] & b[116])^(a[36] & b[117])^(a[35] & b[118])^(a[34] & b[119])^(a[33] & b[120])^(a[32] & b[121])^(a[31] & b[122])^(a[30] & b[123])^(a[29] & b[124])^(a[28] & b[125])^(a[27] & b[126])^(a[26] & b[127])^(a[25] & b[128])^(a[24] & b[129])^(a[23] & b[130])^(a[22] & b[131])^(a[21] & b[132])^(a[20] & b[133])^(a[19] & b[134])^(a[18] & b[135])^(a[17] & b[136])^(a[16] & b[137])^(a[15] & b[138])^(a[14] & b[139])^(a[13] & b[140])^(a[12] & b[141])^(a[11] & b[142])^(a[10] & b[143])^(a[9] & b[144])^(a[8] & b[145])^(a[7] & b[146])^(a[6] & b[147])^(a[5] & b[148])^(a[4] & b[149])^(a[3] & b[150])^(a[2] & b[151])^(a[1] & b[152])^(a[0] & b[153]);
assign y[154] = (a[154] & b[0])^(a[153] & b[1])^(a[152] & b[2])^(a[151] & b[3])^(a[150] & b[4])^(a[149] & b[5])^(a[148] & b[6])^(a[147] & b[7])^(a[146] & b[8])^(a[145] & b[9])^(a[144] & b[10])^(a[143] & b[11])^(a[142] & b[12])^(a[141] & b[13])^(a[140] & b[14])^(a[139] & b[15])^(a[138] & b[16])^(a[137] & b[17])^(a[136] & b[18])^(a[135] & b[19])^(a[134] & b[20])^(a[133] & b[21])^(a[132] & b[22])^(a[131] & b[23])^(a[130] & b[24])^(a[129] & b[25])^(a[128] & b[26])^(a[127] & b[27])^(a[126] & b[28])^(a[125] & b[29])^(a[124] & b[30])^(a[123] & b[31])^(a[122] & b[32])^(a[121] & b[33])^(a[120] & b[34])^(a[119] & b[35])^(a[118] & b[36])^(a[117] & b[37])^(a[116] & b[38])^(a[115] & b[39])^(a[114] & b[40])^(a[113] & b[41])^(a[112] & b[42])^(a[111] & b[43])^(a[110] & b[44])^(a[109] & b[45])^(a[108] & b[46])^(a[107] & b[47])^(a[106] & b[48])^(a[105] & b[49])^(a[104] & b[50])^(a[103] & b[51])^(a[102] & b[52])^(a[101] & b[53])^(a[100] & b[54])^(a[99] & b[55])^(a[98] & b[56])^(a[97] & b[57])^(a[96] & b[58])^(a[95] & b[59])^(a[94] & b[60])^(a[93] & b[61])^(a[92] & b[62])^(a[91] & b[63])^(a[90] & b[64])^(a[89] & b[65])^(a[88] & b[66])^(a[87] & b[67])^(a[86] & b[68])^(a[85] & b[69])^(a[84] & b[70])^(a[83] & b[71])^(a[82] & b[72])^(a[81] & b[73])^(a[80] & b[74])^(a[79] & b[75])^(a[78] & b[76])^(a[77] & b[77])^(a[76] & b[78])^(a[75] & b[79])^(a[74] & b[80])^(a[73] & b[81])^(a[72] & b[82])^(a[71] & b[83])^(a[70] & b[84])^(a[69] & b[85])^(a[68] & b[86])^(a[67] & b[87])^(a[66] & b[88])^(a[65] & b[89])^(a[64] & b[90])^(a[63] & b[91])^(a[62] & b[92])^(a[61] & b[93])^(a[60] & b[94])^(a[59] & b[95])^(a[58] & b[96])^(a[57] & b[97])^(a[56] & b[98])^(a[55] & b[99])^(a[54] & b[100])^(a[53] & b[101])^(a[52] & b[102])^(a[51] & b[103])^(a[50] & b[104])^(a[49] & b[105])^(a[48] & b[106])^(a[47] & b[107])^(a[46] & b[108])^(a[45] & b[109])^(a[44] & b[110])^(a[43] & b[111])^(a[42] & b[112])^(a[41] & b[113])^(a[40] & b[114])^(a[39] & b[115])^(a[38] & b[116])^(a[37] & b[117])^(a[36] & b[118])^(a[35] & b[119])^(a[34] & b[120])^(a[33] & b[121])^(a[32] & b[122])^(a[31] & b[123])^(a[30] & b[124])^(a[29] & b[125])^(a[28] & b[126])^(a[27] & b[127])^(a[26] & b[128])^(a[25] & b[129])^(a[24] & b[130])^(a[23] & b[131])^(a[22] & b[132])^(a[21] & b[133])^(a[20] & b[134])^(a[19] & b[135])^(a[18] & b[136])^(a[17] & b[137])^(a[16] & b[138])^(a[15] & b[139])^(a[14] & b[140])^(a[13] & b[141])^(a[12] & b[142])^(a[11] & b[143])^(a[10] & b[144])^(a[9] & b[145])^(a[8] & b[146])^(a[7] & b[147])^(a[6] & b[148])^(a[5] & b[149])^(a[4] & b[150])^(a[3] & b[151])^(a[2] & b[152])^(a[1] & b[153])^(a[0] & b[154]);
assign y[155] = (a[155] & b[0])^(a[154] & b[1])^(a[153] & b[2])^(a[152] & b[3])^(a[151] & b[4])^(a[150] & b[5])^(a[149] & b[6])^(a[148] & b[7])^(a[147] & b[8])^(a[146] & b[9])^(a[145] & b[10])^(a[144] & b[11])^(a[143] & b[12])^(a[142] & b[13])^(a[141] & b[14])^(a[140] & b[15])^(a[139] & b[16])^(a[138] & b[17])^(a[137] & b[18])^(a[136] & b[19])^(a[135] & b[20])^(a[134] & b[21])^(a[133] & b[22])^(a[132] & b[23])^(a[131] & b[24])^(a[130] & b[25])^(a[129] & b[26])^(a[128] & b[27])^(a[127] & b[28])^(a[126] & b[29])^(a[125] & b[30])^(a[124] & b[31])^(a[123] & b[32])^(a[122] & b[33])^(a[121] & b[34])^(a[120] & b[35])^(a[119] & b[36])^(a[118] & b[37])^(a[117] & b[38])^(a[116] & b[39])^(a[115] & b[40])^(a[114] & b[41])^(a[113] & b[42])^(a[112] & b[43])^(a[111] & b[44])^(a[110] & b[45])^(a[109] & b[46])^(a[108] & b[47])^(a[107] & b[48])^(a[106] & b[49])^(a[105] & b[50])^(a[104] & b[51])^(a[103] & b[52])^(a[102] & b[53])^(a[101] & b[54])^(a[100] & b[55])^(a[99] & b[56])^(a[98] & b[57])^(a[97] & b[58])^(a[96] & b[59])^(a[95] & b[60])^(a[94] & b[61])^(a[93] & b[62])^(a[92] & b[63])^(a[91] & b[64])^(a[90] & b[65])^(a[89] & b[66])^(a[88] & b[67])^(a[87] & b[68])^(a[86] & b[69])^(a[85] & b[70])^(a[84] & b[71])^(a[83] & b[72])^(a[82] & b[73])^(a[81] & b[74])^(a[80] & b[75])^(a[79] & b[76])^(a[78] & b[77])^(a[77] & b[78])^(a[76] & b[79])^(a[75] & b[80])^(a[74] & b[81])^(a[73] & b[82])^(a[72] & b[83])^(a[71] & b[84])^(a[70] & b[85])^(a[69] & b[86])^(a[68] & b[87])^(a[67] & b[88])^(a[66] & b[89])^(a[65] & b[90])^(a[64] & b[91])^(a[63] & b[92])^(a[62] & b[93])^(a[61] & b[94])^(a[60] & b[95])^(a[59] & b[96])^(a[58] & b[97])^(a[57] & b[98])^(a[56] & b[99])^(a[55] & b[100])^(a[54] & b[101])^(a[53] & b[102])^(a[52] & b[103])^(a[51] & b[104])^(a[50] & b[105])^(a[49] & b[106])^(a[48] & b[107])^(a[47] & b[108])^(a[46] & b[109])^(a[45] & b[110])^(a[44] & b[111])^(a[43] & b[112])^(a[42] & b[113])^(a[41] & b[114])^(a[40] & b[115])^(a[39] & b[116])^(a[38] & b[117])^(a[37] & b[118])^(a[36] & b[119])^(a[35] & b[120])^(a[34] & b[121])^(a[33] & b[122])^(a[32] & b[123])^(a[31] & b[124])^(a[30] & b[125])^(a[29] & b[126])^(a[28] & b[127])^(a[27] & b[128])^(a[26] & b[129])^(a[25] & b[130])^(a[24] & b[131])^(a[23] & b[132])^(a[22] & b[133])^(a[21] & b[134])^(a[20] & b[135])^(a[19] & b[136])^(a[18] & b[137])^(a[17] & b[138])^(a[16] & b[139])^(a[15] & b[140])^(a[14] & b[141])^(a[13] & b[142])^(a[12] & b[143])^(a[11] & b[144])^(a[10] & b[145])^(a[9] & b[146])^(a[8] & b[147])^(a[7] & b[148])^(a[6] & b[149])^(a[5] & b[150])^(a[4] & b[151])^(a[3] & b[152])^(a[2] & b[153])^(a[1] & b[154])^(a[0] & b[155]);
assign y[156] = (a[156] & b[0])^(a[155] & b[1])^(a[154] & b[2])^(a[153] & b[3])^(a[152] & b[4])^(a[151] & b[5])^(a[150] & b[6])^(a[149] & b[7])^(a[148] & b[8])^(a[147] & b[9])^(a[146] & b[10])^(a[145] & b[11])^(a[144] & b[12])^(a[143] & b[13])^(a[142] & b[14])^(a[141] & b[15])^(a[140] & b[16])^(a[139] & b[17])^(a[138] & b[18])^(a[137] & b[19])^(a[136] & b[20])^(a[135] & b[21])^(a[134] & b[22])^(a[133] & b[23])^(a[132] & b[24])^(a[131] & b[25])^(a[130] & b[26])^(a[129] & b[27])^(a[128] & b[28])^(a[127] & b[29])^(a[126] & b[30])^(a[125] & b[31])^(a[124] & b[32])^(a[123] & b[33])^(a[122] & b[34])^(a[121] & b[35])^(a[120] & b[36])^(a[119] & b[37])^(a[118] & b[38])^(a[117] & b[39])^(a[116] & b[40])^(a[115] & b[41])^(a[114] & b[42])^(a[113] & b[43])^(a[112] & b[44])^(a[111] & b[45])^(a[110] & b[46])^(a[109] & b[47])^(a[108] & b[48])^(a[107] & b[49])^(a[106] & b[50])^(a[105] & b[51])^(a[104] & b[52])^(a[103] & b[53])^(a[102] & b[54])^(a[101] & b[55])^(a[100] & b[56])^(a[99] & b[57])^(a[98] & b[58])^(a[97] & b[59])^(a[96] & b[60])^(a[95] & b[61])^(a[94] & b[62])^(a[93] & b[63])^(a[92] & b[64])^(a[91] & b[65])^(a[90] & b[66])^(a[89] & b[67])^(a[88] & b[68])^(a[87] & b[69])^(a[86] & b[70])^(a[85] & b[71])^(a[84] & b[72])^(a[83] & b[73])^(a[82] & b[74])^(a[81] & b[75])^(a[80] & b[76])^(a[79] & b[77])^(a[78] & b[78])^(a[77] & b[79])^(a[76] & b[80])^(a[75] & b[81])^(a[74] & b[82])^(a[73] & b[83])^(a[72] & b[84])^(a[71] & b[85])^(a[70] & b[86])^(a[69] & b[87])^(a[68] & b[88])^(a[67] & b[89])^(a[66] & b[90])^(a[65] & b[91])^(a[64] & b[92])^(a[63] & b[93])^(a[62] & b[94])^(a[61] & b[95])^(a[60] & b[96])^(a[59] & b[97])^(a[58] & b[98])^(a[57] & b[99])^(a[56] & b[100])^(a[55] & b[101])^(a[54] & b[102])^(a[53] & b[103])^(a[52] & b[104])^(a[51] & b[105])^(a[50] & b[106])^(a[49] & b[107])^(a[48] & b[108])^(a[47] & b[109])^(a[46] & b[110])^(a[45] & b[111])^(a[44] & b[112])^(a[43] & b[113])^(a[42] & b[114])^(a[41] & b[115])^(a[40] & b[116])^(a[39] & b[117])^(a[38] & b[118])^(a[37] & b[119])^(a[36] & b[120])^(a[35] & b[121])^(a[34] & b[122])^(a[33] & b[123])^(a[32] & b[124])^(a[31] & b[125])^(a[30] & b[126])^(a[29] & b[127])^(a[28] & b[128])^(a[27] & b[129])^(a[26] & b[130])^(a[25] & b[131])^(a[24] & b[132])^(a[23] & b[133])^(a[22] & b[134])^(a[21] & b[135])^(a[20] & b[136])^(a[19] & b[137])^(a[18] & b[138])^(a[17] & b[139])^(a[16] & b[140])^(a[15] & b[141])^(a[14] & b[142])^(a[13] & b[143])^(a[12] & b[144])^(a[11] & b[145])^(a[10] & b[146])^(a[9] & b[147])^(a[8] & b[148])^(a[7] & b[149])^(a[6] & b[150])^(a[5] & b[151])^(a[4] & b[152])^(a[3] & b[153])^(a[2] & b[154])^(a[1] & b[155])^(a[0] & b[156]);
assign y[157] = (a[157] & b[0])^(a[156] & b[1])^(a[155] & b[2])^(a[154] & b[3])^(a[153] & b[4])^(a[152] & b[5])^(a[151] & b[6])^(a[150] & b[7])^(a[149] & b[8])^(a[148] & b[9])^(a[147] & b[10])^(a[146] & b[11])^(a[145] & b[12])^(a[144] & b[13])^(a[143] & b[14])^(a[142] & b[15])^(a[141] & b[16])^(a[140] & b[17])^(a[139] & b[18])^(a[138] & b[19])^(a[137] & b[20])^(a[136] & b[21])^(a[135] & b[22])^(a[134] & b[23])^(a[133] & b[24])^(a[132] & b[25])^(a[131] & b[26])^(a[130] & b[27])^(a[129] & b[28])^(a[128] & b[29])^(a[127] & b[30])^(a[126] & b[31])^(a[125] & b[32])^(a[124] & b[33])^(a[123] & b[34])^(a[122] & b[35])^(a[121] & b[36])^(a[120] & b[37])^(a[119] & b[38])^(a[118] & b[39])^(a[117] & b[40])^(a[116] & b[41])^(a[115] & b[42])^(a[114] & b[43])^(a[113] & b[44])^(a[112] & b[45])^(a[111] & b[46])^(a[110] & b[47])^(a[109] & b[48])^(a[108] & b[49])^(a[107] & b[50])^(a[106] & b[51])^(a[105] & b[52])^(a[104] & b[53])^(a[103] & b[54])^(a[102] & b[55])^(a[101] & b[56])^(a[100] & b[57])^(a[99] & b[58])^(a[98] & b[59])^(a[97] & b[60])^(a[96] & b[61])^(a[95] & b[62])^(a[94] & b[63])^(a[93] & b[64])^(a[92] & b[65])^(a[91] & b[66])^(a[90] & b[67])^(a[89] & b[68])^(a[88] & b[69])^(a[87] & b[70])^(a[86] & b[71])^(a[85] & b[72])^(a[84] & b[73])^(a[83] & b[74])^(a[82] & b[75])^(a[81] & b[76])^(a[80] & b[77])^(a[79] & b[78])^(a[78] & b[79])^(a[77] & b[80])^(a[76] & b[81])^(a[75] & b[82])^(a[74] & b[83])^(a[73] & b[84])^(a[72] & b[85])^(a[71] & b[86])^(a[70] & b[87])^(a[69] & b[88])^(a[68] & b[89])^(a[67] & b[90])^(a[66] & b[91])^(a[65] & b[92])^(a[64] & b[93])^(a[63] & b[94])^(a[62] & b[95])^(a[61] & b[96])^(a[60] & b[97])^(a[59] & b[98])^(a[58] & b[99])^(a[57] & b[100])^(a[56] & b[101])^(a[55] & b[102])^(a[54] & b[103])^(a[53] & b[104])^(a[52] & b[105])^(a[51] & b[106])^(a[50] & b[107])^(a[49] & b[108])^(a[48] & b[109])^(a[47] & b[110])^(a[46] & b[111])^(a[45] & b[112])^(a[44] & b[113])^(a[43] & b[114])^(a[42] & b[115])^(a[41] & b[116])^(a[40] & b[117])^(a[39] & b[118])^(a[38] & b[119])^(a[37] & b[120])^(a[36] & b[121])^(a[35] & b[122])^(a[34] & b[123])^(a[33] & b[124])^(a[32] & b[125])^(a[31] & b[126])^(a[30] & b[127])^(a[29] & b[128])^(a[28] & b[129])^(a[27] & b[130])^(a[26] & b[131])^(a[25] & b[132])^(a[24] & b[133])^(a[23] & b[134])^(a[22] & b[135])^(a[21] & b[136])^(a[20] & b[137])^(a[19] & b[138])^(a[18] & b[139])^(a[17] & b[140])^(a[16] & b[141])^(a[15] & b[142])^(a[14] & b[143])^(a[13] & b[144])^(a[12] & b[145])^(a[11] & b[146])^(a[10] & b[147])^(a[9] & b[148])^(a[8] & b[149])^(a[7] & b[150])^(a[6] & b[151])^(a[5] & b[152])^(a[4] & b[153])^(a[3] & b[154])^(a[2] & b[155])^(a[1] & b[156])^(a[0] & b[157]);
assign y[158] = (a[158] & b[0])^(a[157] & b[1])^(a[156] & b[2])^(a[155] & b[3])^(a[154] & b[4])^(a[153] & b[5])^(a[152] & b[6])^(a[151] & b[7])^(a[150] & b[8])^(a[149] & b[9])^(a[148] & b[10])^(a[147] & b[11])^(a[146] & b[12])^(a[145] & b[13])^(a[144] & b[14])^(a[143] & b[15])^(a[142] & b[16])^(a[141] & b[17])^(a[140] & b[18])^(a[139] & b[19])^(a[138] & b[20])^(a[137] & b[21])^(a[136] & b[22])^(a[135] & b[23])^(a[134] & b[24])^(a[133] & b[25])^(a[132] & b[26])^(a[131] & b[27])^(a[130] & b[28])^(a[129] & b[29])^(a[128] & b[30])^(a[127] & b[31])^(a[126] & b[32])^(a[125] & b[33])^(a[124] & b[34])^(a[123] & b[35])^(a[122] & b[36])^(a[121] & b[37])^(a[120] & b[38])^(a[119] & b[39])^(a[118] & b[40])^(a[117] & b[41])^(a[116] & b[42])^(a[115] & b[43])^(a[114] & b[44])^(a[113] & b[45])^(a[112] & b[46])^(a[111] & b[47])^(a[110] & b[48])^(a[109] & b[49])^(a[108] & b[50])^(a[107] & b[51])^(a[106] & b[52])^(a[105] & b[53])^(a[104] & b[54])^(a[103] & b[55])^(a[102] & b[56])^(a[101] & b[57])^(a[100] & b[58])^(a[99] & b[59])^(a[98] & b[60])^(a[97] & b[61])^(a[96] & b[62])^(a[95] & b[63])^(a[94] & b[64])^(a[93] & b[65])^(a[92] & b[66])^(a[91] & b[67])^(a[90] & b[68])^(a[89] & b[69])^(a[88] & b[70])^(a[87] & b[71])^(a[86] & b[72])^(a[85] & b[73])^(a[84] & b[74])^(a[83] & b[75])^(a[82] & b[76])^(a[81] & b[77])^(a[80] & b[78])^(a[79] & b[79])^(a[78] & b[80])^(a[77] & b[81])^(a[76] & b[82])^(a[75] & b[83])^(a[74] & b[84])^(a[73] & b[85])^(a[72] & b[86])^(a[71] & b[87])^(a[70] & b[88])^(a[69] & b[89])^(a[68] & b[90])^(a[67] & b[91])^(a[66] & b[92])^(a[65] & b[93])^(a[64] & b[94])^(a[63] & b[95])^(a[62] & b[96])^(a[61] & b[97])^(a[60] & b[98])^(a[59] & b[99])^(a[58] & b[100])^(a[57] & b[101])^(a[56] & b[102])^(a[55] & b[103])^(a[54] & b[104])^(a[53] & b[105])^(a[52] & b[106])^(a[51] & b[107])^(a[50] & b[108])^(a[49] & b[109])^(a[48] & b[110])^(a[47] & b[111])^(a[46] & b[112])^(a[45] & b[113])^(a[44] & b[114])^(a[43] & b[115])^(a[42] & b[116])^(a[41] & b[117])^(a[40] & b[118])^(a[39] & b[119])^(a[38] & b[120])^(a[37] & b[121])^(a[36] & b[122])^(a[35] & b[123])^(a[34] & b[124])^(a[33] & b[125])^(a[32] & b[126])^(a[31] & b[127])^(a[30] & b[128])^(a[29] & b[129])^(a[28] & b[130])^(a[27] & b[131])^(a[26] & b[132])^(a[25] & b[133])^(a[24] & b[134])^(a[23] & b[135])^(a[22] & b[136])^(a[21] & b[137])^(a[20] & b[138])^(a[19] & b[139])^(a[18] & b[140])^(a[17] & b[141])^(a[16] & b[142])^(a[15] & b[143])^(a[14] & b[144])^(a[13] & b[145])^(a[12] & b[146])^(a[11] & b[147])^(a[10] & b[148])^(a[9] & b[149])^(a[8] & b[150])^(a[7] & b[151])^(a[6] & b[152])^(a[5] & b[153])^(a[4] & b[154])^(a[3] & b[155])^(a[2] & b[156])^(a[1] & b[157])^(a[0] & b[158]);
assign y[159] = (a[159] & b[0])^(a[158] & b[1])^(a[157] & b[2])^(a[156] & b[3])^(a[155] & b[4])^(a[154] & b[5])^(a[153] & b[6])^(a[152] & b[7])^(a[151] & b[8])^(a[150] & b[9])^(a[149] & b[10])^(a[148] & b[11])^(a[147] & b[12])^(a[146] & b[13])^(a[145] & b[14])^(a[144] & b[15])^(a[143] & b[16])^(a[142] & b[17])^(a[141] & b[18])^(a[140] & b[19])^(a[139] & b[20])^(a[138] & b[21])^(a[137] & b[22])^(a[136] & b[23])^(a[135] & b[24])^(a[134] & b[25])^(a[133] & b[26])^(a[132] & b[27])^(a[131] & b[28])^(a[130] & b[29])^(a[129] & b[30])^(a[128] & b[31])^(a[127] & b[32])^(a[126] & b[33])^(a[125] & b[34])^(a[124] & b[35])^(a[123] & b[36])^(a[122] & b[37])^(a[121] & b[38])^(a[120] & b[39])^(a[119] & b[40])^(a[118] & b[41])^(a[117] & b[42])^(a[116] & b[43])^(a[115] & b[44])^(a[114] & b[45])^(a[113] & b[46])^(a[112] & b[47])^(a[111] & b[48])^(a[110] & b[49])^(a[109] & b[50])^(a[108] & b[51])^(a[107] & b[52])^(a[106] & b[53])^(a[105] & b[54])^(a[104] & b[55])^(a[103] & b[56])^(a[102] & b[57])^(a[101] & b[58])^(a[100] & b[59])^(a[99] & b[60])^(a[98] & b[61])^(a[97] & b[62])^(a[96] & b[63])^(a[95] & b[64])^(a[94] & b[65])^(a[93] & b[66])^(a[92] & b[67])^(a[91] & b[68])^(a[90] & b[69])^(a[89] & b[70])^(a[88] & b[71])^(a[87] & b[72])^(a[86] & b[73])^(a[85] & b[74])^(a[84] & b[75])^(a[83] & b[76])^(a[82] & b[77])^(a[81] & b[78])^(a[80] & b[79])^(a[79] & b[80])^(a[78] & b[81])^(a[77] & b[82])^(a[76] & b[83])^(a[75] & b[84])^(a[74] & b[85])^(a[73] & b[86])^(a[72] & b[87])^(a[71] & b[88])^(a[70] & b[89])^(a[69] & b[90])^(a[68] & b[91])^(a[67] & b[92])^(a[66] & b[93])^(a[65] & b[94])^(a[64] & b[95])^(a[63] & b[96])^(a[62] & b[97])^(a[61] & b[98])^(a[60] & b[99])^(a[59] & b[100])^(a[58] & b[101])^(a[57] & b[102])^(a[56] & b[103])^(a[55] & b[104])^(a[54] & b[105])^(a[53] & b[106])^(a[52] & b[107])^(a[51] & b[108])^(a[50] & b[109])^(a[49] & b[110])^(a[48] & b[111])^(a[47] & b[112])^(a[46] & b[113])^(a[45] & b[114])^(a[44] & b[115])^(a[43] & b[116])^(a[42] & b[117])^(a[41] & b[118])^(a[40] & b[119])^(a[39] & b[120])^(a[38] & b[121])^(a[37] & b[122])^(a[36] & b[123])^(a[35] & b[124])^(a[34] & b[125])^(a[33] & b[126])^(a[32] & b[127])^(a[31] & b[128])^(a[30] & b[129])^(a[29] & b[130])^(a[28] & b[131])^(a[27] & b[132])^(a[26] & b[133])^(a[25] & b[134])^(a[24] & b[135])^(a[23] & b[136])^(a[22] & b[137])^(a[21] & b[138])^(a[20] & b[139])^(a[19] & b[140])^(a[18] & b[141])^(a[17] & b[142])^(a[16] & b[143])^(a[15] & b[144])^(a[14] & b[145])^(a[13] & b[146])^(a[12] & b[147])^(a[11] & b[148])^(a[10] & b[149])^(a[9] & b[150])^(a[8] & b[151])^(a[7] & b[152])^(a[6] & b[153])^(a[5] & b[154])^(a[4] & b[155])^(a[3] & b[156])^(a[2] & b[157])^(a[1] & b[158])^(a[0] & b[159]);
assign y[160] = (a[160] & b[0])^(a[159] & b[1])^(a[158] & b[2])^(a[157] & b[3])^(a[156] & b[4])^(a[155] & b[5])^(a[154] & b[6])^(a[153] & b[7])^(a[152] & b[8])^(a[151] & b[9])^(a[150] & b[10])^(a[149] & b[11])^(a[148] & b[12])^(a[147] & b[13])^(a[146] & b[14])^(a[145] & b[15])^(a[144] & b[16])^(a[143] & b[17])^(a[142] & b[18])^(a[141] & b[19])^(a[140] & b[20])^(a[139] & b[21])^(a[138] & b[22])^(a[137] & b[23])^(a[136] & b[24])^(a[135] & b[25])^(a[134] & b[26])^(a[133] & b[27])^(a[132] & b[28])^(a[131] & b[29])^(a[130] & b[30])^(a[129] & b[31])^(a[128] & b[32])^(a[127] & b[33])^(a[126] & b[34])^(a[125] & b[35])^(a[124] & b[36])^(a[123] & b[37])^(a[122] & b[38])^(a[121] & b[39])^(a[120] & b[40])^(a[119] & b[41])^(a[118] & b[42])^(a[117] & b[43])^(a[116] & b[44])^(a[115] & b[45])^(a[114] & b[46])^(a[113] & b[47])^(a[112] & b[48])^(a[111] & b[49])^(a[110] & b[50])^(a[109] & b[51])^(a[108] & b[52])^(a[107] & b[53])^(a[106] & b[54])^(a[105] & b[55])^(a[104] & b[56])^(a[103] & b[57])^(a[102] & b[58])^(a[101] & b[59])^(a[100] & b[60])^(a[99] & b[61])^(a[98] & b[62])^(a[97] & b[63])^(a[96] & b[64])^(a[95] & b[65])^(a[94] & b[66])^(a[93] & b[67])^(a[92] & b[68])^(a[91] & b[69])^(a[90] & b[70])^(a[89] & b[71])^(a[88] & b[72])^(a[87] & b[73])^(a[86] & b[74])^(a[85] & b[75])^(a[84] & b[76])^(a[83] & b[77])^(a[82] & b[78])^(a[81] & b[79])^(a[80] & b[80])^(a[79] & b[81])^(a[78] & b[82])^(a[77] & b[83])^(a[76] & b[84])^(a[75] & b[85])^(a[74] & b[86])^(a[73] & b[87])^(a[72] & b[88])^(a[71] & b[89])^(a[70] & b[90])^(a[69] & b[91])^(a[68] & b[92])^(a[67] & b[93])^(a[66] & b[94])^(a[65] & b[95])^(a[64] & b[96])^(a[63] & b[97])^(a[62] & b[98])^(a[61] & b[99])^(a[60] & b[100])^(a[59] & b[101])^(a[58] & b[102])^(a[57] & b[103])^(a[56] & b[104])^(a[55] & b[105])^(a[54] & b[106])^(a[53] & b[107])^(a[52] & b[108])^(a[51] & b[109])^(a[50] & b[110])^(a[49] & b[111])^(a[48] & b[112])^(a[47] & b[113])^(a[46] & b[114])^(a[45] & b[115])^(a[44] & b[116])^(a[43] & b[117])^(a[42] & b[118])^(a[41] & b[119])^(a[40] & b[120])^(a[39] & b[121])^(a[38] & b[122])^(a[37] & b[123])^(a[36] & b[124])^(a[35] & b[125])^(a[34] & b[126])^(a[33] & b[127])^(a[32] & b[128])^(a[31] & b[129])^(a[30] & b[130])^(a[29] & b[131])^(a[28] & b[132])^(a[27] & b[133])^(a[26] & b[134])^(a[25] & b[135])^(a[24] & b[136])^(a[23] & b[137])^(a[22] & b[138])^(a[21] & b[139])^(a[20] & b[140])^(a[19] & b[141])^(a[18] & b[142])^(a[17] & b[143])^(a[16] & b[144])^(a[15] & b[145])^(a[14] & b[146])^(a[13] & b[147])^(a[12] & b[148])^(a[11] & b[149])^(a[10] & b[150])^(a[9] & b[151])^(a[8] & b[152])^(a[7] & b[153])^(a[6] & b[154])^(a[5] & b[155])^(a[4] & b[156])^(a[3] & b[157])^(a[2] & b[158])^(a[1] & b[159])^(a[0] & b[160]);
assign y[161] = (a[161] & b[0])^(a[160] & b[1])^(a[159] & b[2])^(a[158] & b[3])^(a[157] & b[4])^(a[156] & b[5])^(a[155] & b[6])^(a[154] & b[7])^(a[153] & b[8])^(a[152] & b[9])^(a[151] & b[10])^(a[150] & b[11])^(a[149] & b[12])^(a[148] & b[13])^(a[147] & b[14])^(a[146] & b[15])^(a[145] & b[16])^(a[144] & b[17])^(a[143] & b[18])^(a[142] & b[19])^(a[141] & b[20])^(a[140] & b[21])^(a[139] & b[22])^(a[138] & b[23])^(a[137] & b[24])^(a[136] & b[25])^(a[135] & b[26])^(a[134] & b[27])^(a[133] & b[28])^(a[132] & b[29])^(a[131] & b[30])^(a[130] & b[31])^(a[129] & b[32])^(a[128] & b[33])^(a[127] & b[34])^(a[126] & b[35])^(a[125] & b[36])^(a[124] & b[37])^(a[123] & b[38])^(a[122] & b[39])^(a[121] & b[40])^(a[120] & b[41])^(a[119] & b[42])^(a[118] & b[43])^(a[117] & b[44])^(a[116] & b[45])^(a[115] & b[46])^(a[114] & b[47])^(a[113] & b[48])^(a[112] & b[49])^(a[111] & b[50])^(a[110] & b[51])^(a[109] & b[52])^(a[108] & b[53])^(a[107] & b[54])^(a[106] & b[55])^(a[105] & b[56])^(a[104] & b[57])^(a[103] & b[58])^(a[102] & b[59])^(a[101] & b[60])^(a[100] & b[61])^(a[99] & b[62])^(a[98] & b[63])^(a[97] & b[64])^(a[96] & b[65])^(a[95] & b[66])^(a[94] & b[67])^(a[93] & b[68])^(a[92] & b[69])^(a[91] & b[70])^(a[90] & b[71])^(a[89] & b[72])^(a[88] & b[73])^(a[87] & b[74])^(a[86] & b[75])^(a[85] & b[76])^(a[84] & b[77])^(a[83] & b[78])^(a[82] & b[79])^(a[81] & b[80])^(a[80] & b[81])^(a[79] & b[82])^(a[78] & b[83])^(a[77] & b[84])^(a[76] & b[85])^(a[75] & b[86])^(a[74] & b[87])^(a[73] & b[88])^(a[72] & b[89])^(a[71] & b[90])^(a[70] & b[91])^(a[69] & b[92])^(a[68] & b[93])^(a[67] & b[94])^(a[66] & b[95])^(a[65] & b[96])^(a[64] & b[97])^(a[63] & b[98])^(a[62] & b[99])^(a[61] & b[100])^(a[60] & b[101])^(a[59] & b[102])^(a[58] & b[103])^(a[57] & b[104])^(a[56] & b[105])^(a[55] & b[106])^(a[54] & b[107])^(a[53] & b[108])^(a[52] & b[109])^(a[51] & b[110])^(a[50] & b[111])^(a[49] & b[112])^(a[48] & b[113])^(a[47] & b[114])^(a[46] & b[115])^(a[45] & b[116])^(a[44] & b[117])^(a[43] & b[118])^(a[42] & b[119])^(a[41] & b[120])^(a[40] & b[121])^(a[39] & b[122])^(a[38] & b[123])^(a[37] & b[124])^(a[36] & b[125])^(a[35] & b[126])^(a[34] & b[127])^(a[33] & b[128])^(a[32] & b[129])^(a[31] & b[130])^(a[30] & b[131])^(a[29] & b[132])^(a[28] & b[133])^(a[27] & b[134])^(a[26] & b[135])^(a[25] & b[136])^(a[24] & b[137])^(a[23] & b[138])^(a[22] & b[139])^(a[21] & b[140])^(a[20] & b[141])^(a[19] & b[142])^(a[18] & b[143])^(a[17] & b[144])^(a[16] & b[145])^(a[15] & b[146])^(a[14] & b[147])^(a[13] & b[148])^(a[12] & b[149])^(a[11] & b[150])^(a[10] & b[151])^(a[9] & b[152])^(a[8] & b[153])^(a[7] & b[154])^(a[6] & b[155])^(a[5] & b[156])^(a[4] & b[157])^(a[3] & b[158])^(a[2] & b[159])^(a[1] & b[160])^(a[0] & b[161]);
assign y[162] = (a[162] & b[0])^(a[161] & b[1])^(a[160] & b[2])^(a[159] & b[3])^(a[158] & b[4])^(a[157] & b[5])^(a[156] & b[6])^(a[155] & b[7])^(a[154] & b[8])^(a[153] & b[9])^(a[152] & b[10])^(a[151] & b[11])^(a[150] & b[12])^(a[149] & b[13])^(a[148] & b[14])^(a[147] & b[15])^(a[146] & b[16])^(a[145] & b[17])^(a[144] & b[18])^(a[143] & b[19])^(a[142] & b[20])^(a[141] & b[21])^(a[140] & b[22])^(a[139] & b[23])^(a[138] & b[24])^(a[137] & b[25])^(a[136] & b[26])^(a[135] & b[27])^(a[134] & b[28])^(a[133] & b[29])^(a[132] & b[30])^(a[131] & b[31])^(a[130] & b[32])^(a[129] & b[33])^(a[128] & b[34])^(a[127] & b[35])^(a[126] & b[36])^(a[125] & b[37])^(a[124] & b[38])^(a[123] & b[39])^(a[122] & b[40])^(a[121] & b[41])^(a[120] & b[42])^(a[119] & b[43])^(a[118] & b[44])^(a[117] & b[45])^(a[116] & b[46])^(a[115] & b[47])^(a[114] & b[48])^(a[113] & b[49])^(a[112] & b[50])^(a[111] & b[51])^(a[110] & b[52])^(a[109] & b[53])^(a[108] & b[54])^(a[107] & b[55])^(a[106] & b[56])^(a[105] & b[57])^(a[104] & b[58])^(a[103] & b[59])^(a[102] & b[60])^(a[101] & b[61])^(a[100] & b[62])^(a[99] & b[63])^(a[98] & b[64])^(a[97] & b[65])^(a[96] & b[66])^(a[95] & b[67])^(a[94] & b[68])^(a[93] & b[69])^(a[92] & b[70])^(a[91] & b[71])^(a[90] & b[72])^(a[89] & b[73])^(a[88] & b[74])^(a[87] & b[75])^(a[86] & b[76])^(a[85] & b[77])^(a[84] & b[78])^(a[83] & b[79])^(a[82] & b[80])^(a[81] & b[81])^(a[80] & b[82])^(a[79] & b[83])^(a[78] & b[84])^(a[77] & b[85])^(a[76] & b[86])^(a[75] & b[87])^(a[74] & b[88])^(a[73] & b[89])^(a[72] & b[90])^(a[71] & b[91])^(a[70] & b[92])^(a[69] & b[93])^(a[68] & b[94])^(a[67] & b[95])^(a[66] & b[96])^(a[65] & b[97])^(a[64] & b[98])^(a[63] & b[99])^(a[62] & b[100])^(a[61] & b[101])^(a[60] & b[102])^(a[59] & b[103])^(a[58] & b[104])^(a[57] & b[105])^(a[56] & b[106])^(a[55] & b[107])^(a[54] & b[108])^(a[53] & b[109])^(a[52] & b[110])^(a[51] & b[111])^(a[50] & b[112])^(a[49] & b[113])^(a[48] & b[114])^(a[47] & b[115])^(a[46] & b[116])^(a[45] & b[117])^(a[44] & b[118])^(a[43] & b[119])^(a[42] & b[120])^(a[41] & b[121])^(a[40] & b[122])^(a[39] & b[123])^(a[38] & b[124])^(a[37] & b[125])^(a[36] & b[126])^(a[35] & b[127])^(a[34] & b[128])^(a[33] & b[129])^(a[32] & b[130])^(a[31] & b[131])^(a[30] & b[132])^(a[29] & b[133])^(a[28] & b[134])^(a[27] & b[135])^(a[26] & b[136])^(a[25] & b[137])^(a[24] & b[138])^(a[23] & b[139])^(a[22] & b[140])^(a[21] & b[141])^(a[20] & b[142])^(a[19] & b[143])^(a[18] & b[144])^(a[17] & b[145])^(a[16] & b[146])^(a[15] & b[147])^(a[14] & b[148])^(a[13] & b[149])^(a[12] & b[150])^(a[11] & b[151])^(a[10] & b[152])^(a[9] & b[153])^(a[8] & b[154])^(a[7] & b[155])^(a[6] & b[156])^(a[5] & b[157])^(a[4] & b[158])^(a[3] & b[159])^(a[2] & b[160])^(a[1] & b[161])^(a[0] & b[162]);
assign y[163] = (a[163] & b[0])^(a[162] & b[1])^(a[161] & b[2])^(a[160] & b[3])^(a[159] & b[4])^(a[158] & b[5])^(a[157] & b[6])^(a[156] & b[7])^(a[155] & b[8])^(a[154] & b[9])^(a[153] & b[10])^(a[152] & b[11])^(a[151] & b[12])^(a[150] & b[13])^(a[149] & b[14])^(a[148] & b[15])^(a[147] & b[16])^(a[146] & b[17])^(a[145] & b[18])^(a[144] & b[19])^(a[143] & b[20])^(a[142] & b[21])^(a[141] & b[22])^(a[140] & b[23])^(a[139] & b[24])^(a[138] & b[25])^(a[137] & b[26])^(a[136] & b[27])^(a[135] & b[28])^(a[134] & b[29])^(a[133] & b[30])^(a[132] & b[31])^(a[131] & b[32])^(a[130] & b[33])^(a[129] & b[34])^(a[128] & b[35])^(a[127] & b[36])^(a[126] & b[37])^(a[125] & b[38])^(a[124] & b[39])^(a[123] & b[40])^(a[122] & b[41])^(a[121] & b[42])^(a[120] & b[43])^(a[119] & b[44])^(a[118] & b[45])^(a[117] & b[46])^(a[116] & b[47])^(a[115] & b[48])^(a[114] & b[49])^(a[113] & b[50])^(a[112] & b[51])^(a[111] & b[52])^(a[110] & b[53])^(a[109] & b[54])^(a[108] & b[55])^(a[107] & b[56])^(a[106] & b[57])^(a[105] & b[58])^(a[104] & b[59])^(a[103] & b[60])^(a[102] & b[61])^(a[101] & b[62])^(a[100] & b[63])^(a[99] & b[64])^(a[98] & b[65])^(a[97] & b[66])^(a[96] & b[67])^(a[95] & b[68])^(a[94] & b[69])^(a[93] & b[70])^(a[92] & b[71])^(a[91] & b[72])^(a[90] & b[73])^(a[89] & b[74])^(a[88] & b[75])^(a[87] & b[76])^(a[86] & b[77])^(a[85] & b[78])^(a[84] & b[79])^(a[83] & b[80])^(a[82] & b[81])^(a[81] & b[82])^(a[80] & b[83])^(a[79] & b[84])^(a[78] & b[85])^(a[77] & b[86])^(a[76] & b[87])^(a[75] & b[88])^(a[74] & b[89])^(a[73] & b[90])^(a[72] & b[91])^(a[71] & b[92])^(a[70] & b[93])^(a[69] & b[94])^(a[68] & b[95])^(a[67] & b[96])^(a[66] & b[97])^(a[65] & b[98])^(a[64] & b[99])^(a[63] & b[100])^(a[62] & b[101])^(a[61] & b[102])^(a[60] & b[103])^(a[59] & b[104])^(a[58] & b[105])^(a[57] & b[106])^(a[56] & b[107])^(a[55] & b[108])^(a[54] & b[109])^(a[53] & b[110])^(a[52] & b[111])^(a[51] & b[112])^(a[50] & b[113])^(a[49] & b[114])^(a[48] & b[115])^(a[47] & b[116])^(a[46] & b[117])^(a[45] & b[118])^(a[44] & b[119])^(a[43] & b[120])^(a[42] & b[121])^(a[41] & b[122])^(a[40] & b[123])^(a[39] & b[124])^(a[38] & b[125])^(a[37] & b[126])^(a[36] & b[127])^(a[35] & b[128])^(a[34] & b[129])^(a[33] & b[130])^(a[32] & b[131])^(a[31] & b[132])^(a[30] & b[133])^(a[29] & b[134])^(a[28] & b[135])^(a[27] & b[136])^(a[26] & b[137])^(a[25] & b[138])^(a[24] & b[139])^(a[23] & b[140])^(a[22] & b[141])^(a[21] & b[142])^(a[20] & b[143])^(a[19] & b[144])^(a[18] & b[145])^(a[17] & b[146])^(a[16] & b[147])^(a[15] & b[148])^(a[14] & b[149])^(a[13] & b[150])^(a[12] & b[151])^(a[11] & b[152])^(a[10] & b[153])^(a[9] & b[154])^(a[8] & b[155])^(a[7] & b[156])^(a[6] & b[157])^(a[5] & b[158])^(a[4] & b[159])^(a[3] & b[160])^(a[2] & b[161])^(a[1] & b[162])^(a[0] & b[163]);
assign y[164] = (a[164] & b[0])^(a[163] & b[1])^(a[162] & b[2])^(a[161] & b[3])^(a[160] & b[4])^(a[159] & b[5])^(a[158] & b[6])^(a[157] & b[7])^(a[156] & b[8])^(a[155] & b[9])^(a[154] & b[10])^(a[153] & b[11])^(a[152] & b[12])^(a[151] & b[13])^(a[150] & b[14])^(a[149] & b[15])^(a[148] & b[16])^(a[147] & b[17])^(a[146] & b[18])^(a[145] & b[19])^(a[144] & b[20])^(a[143] & b[21])^(a[142] & b[22])^(a[141] & b[23])^(a[140] & b[24])^(a[139] & b[25])^(a[138] & b[26])^(a[137] & b[27])^(a[136] & b[28])^(a[135] & b[29])^(a[134] & b[30])^(a[133] & b[31])^(a[132] & b[32])^(a[131] & b[33])^(a[130] & b[34])^(a[129] & b[35])^(a[128] & b[36])^(a[127] & b[37])^(a[126] & b[38])^(a[125] & b[39])^(a[124] & b[40])^(a[123] & b[41])^(a[122] & b[42])^(a[121] & b[43])^(a[120] & b[44])^(a[119] & b[45])^(a[118] & b[46])^(a[117] & b[47])^(a[116] & b[48])^(a[115] & b[49])^(a[114] & b[50])^(a[113] & b[51])^(a[112] & b[52])^(a[111] & b[53])^(a[110] & b[54])^(a[109] & b[55])^(a[108] & b[56])^(a[107] & b[57])^(a[106] & b[58])^(a[105] & b[59])^(a[104] & b[60])^(a[103] & b[61])^(a[102] & b[62])^(a[101] & b[63])^(a[100] & b[64])^(a[99] & b[65])^(a[98] & b[66])^(a[97] & b[67])^(a[96] & b[68])^(a[95] & b[69])^(a[94] & b[70])^(a[93] & b[71])^(a[92] & b[72])^(a[91] & b[73])^(a[90] & b[74])^(a[89] & b[75])^(a[88] & b[76])^(a[87] & b[77])^(a[86] & b[78])^(a[85] & b[79])^(a[84] & b[80])^(a[83] & b[81])^(a[82] & b[82])^(a[81] & b[83])^(a[80] & b[84])^(a[79] & b[85])^(a[78] & b[86])^(a[77] & b[87])^(a[76] & b[88])^(a[75] & b[89])^(a[74] & b[90])^(a[73] & b[91])^(a[72] & b[92])^(a[71] & b[93])^(a[70] & b[94])^(a[69] & b[95])^(a[68] & b[96])^(a[67] & b[97])^(a[66] & b[98])^(a[65] & b[99])^(a[64] & b[100])^(a[63] & b[101])^(a[62] & b[102])^(a[61] & b[103])^(a[60] & b[104])^(a[59] & b[105])^(a[58] & b[106])^(a[57] & b[107])^(a[56] & b[108])^(a[55] & b[109])^(a[54] & b[110])^(a[53] & b[111])^(a[52] & b[112])^(a[51] & b[113])^(a[50] & b[114])^(a[49] & b[115])^(a[48] & b[116])^(a[47] & b[117])^(a[46] & b[118])^(a[45] & b[119])^(a[44] & b[120])^(a[43] & b[121])^(a[42] & b[122])^(a[41] & b[123])^(a[40] & b[124])^(a[39] & b[125])^(a[38] & b[126])^(a[37] & b[127])^(a[36] & b[128])^(a[35] & b[129])^(a[34] & b[130])^(a[33] & b[131])^(a[32] & b[132])^(a[31] & b[133])^(a[30] & b[134])^(a[29] & b[135])^(a[28] & b[136])^(a[27] & b[137])^(a[26] & b[138])^(a[25] & b[139])^(a[24] & b[140])^(a[23] & b[141])^(a[22] & b[142])^(a[21] & b[143])^(a[20] & b[144])^(a[19] & b[145])^(a[18] & b[146])^(a[17] & b[147])^(a[16] & b[148])^(a[15] & b[149])^(a[14] & b[150])^(a[13] & b[151])^(a[12] & b[152])^(a[11] & b[153])^(a[10] & b[154])^(a[9] & b[155])^(a[8] & b[156])^(a[7] & b[157])^(a[6] & b[158])^(a[5] & b[159])^(a[4] & b[160])^(a[3] & b[161])^(a[2] & b[162])^(a[1] & b[163])^(a[0] & b[164]);
assign y[165] = (a[165] & b[0])^(a[164] & b[1])^(a[163] & b[2])^(a[162] & b[3])^(a[161] & b[4])^(a[160] & b[5])^(a[159] & b[6])^(a[158] & b[7])^(a[157] & b[8])^(a[156] & b[9])^(a[155] & b[10])^(a[154] & b[11])^(a[153] & b[12])^(a[152] & b[13])^(a[151] & b[14])^(a[150] & b[15])^(a[149] & b[16])^(a[148] & b[17])^(a[147] & b[18])^(a[146] & b[19])^(a[145] & b[20])^(a[144] & b[21])^(a[143] & b[22])^(a[142] & b[23])^(a[141] & b[24])^(a[140] & b[25])^(a[139] & b[26])^(a[138] & b[27])^(a[137] & b[28])^(a[136] & b[29])^(a[135] & b[30])^(a[134] & b[31])^(a[133] & b[32])^(a[132] & b[33])^(a[131] & b[34])^(a[130] & b[35])^(a[129] & b[36])^(a[128] & b[37])^(a[127] & b[38])^(a[126] & b[39])^(a[125] & b[40])^(a[124] & b[41])^(a[123] & b[42])^(a[122] & b[43])^(a[121] & b[44])^(a[120] & b[45])^(a[119] & b[46])^(a[118] & b[47])^(a[117] & b[48])^(a[116] & b[49])^(a[115] & b[50])^(a[114] & b[51])^(a[113] & b[52])^(a[112] & b[53])^(a[111] & b[54])^(a[110] & b[55])^(a[109] & b[56])^(a[108] & b[57])^(a[107] & b[58])^(a[106] & b[59])^(a[105] & b[60])^(a[104] & b[61])^(a[103] & b[62])^(a[102] & b[63])^(a[101] & b[64])^(a[100] & b[65])^(a[99] & b[66])^(a[98] & b[67])^(a[97] & b[68])^(a[96] & b[69])^(a[95] & b[70])^(a[94] & b[71])^(a[93] & b[72])^(a[92] & b[73])^(a[91] & b[74])^(a[90] & b[75])^(a[89] & b[76])^(a[88] & b[77])^(a[87] & b[78])^(a[86] & b[79])^(a[85] & b[80])^(a[84] & b[81])^(a[83] & b[82])^(a[82] & b[83])^(a[81] & b[84])^(a[80] & b[85])^(a[79] & b[86])^(a[78] & b[87])^(a[77] & b[88])^(a[76] & b[89])^(a[75] & b[90])^(a[74] & b[91])^(a[73] & b[92])^(a[72] & b[93])^(a[71] & b[94])^(a[70] & b[95])^(a[69] & b[96])^(a[68] & b[97])^(a[67] & b[98])^(a[66] & b[99])^(a[65] & b[100])^(a[64] & b[101])^(a[63] & b[102])^(a[62] & b[103])^(a[61] & b[104])^(a[60] & b[105])^(a[59] & b[106])^(a[58] & b[107])^(a[57] & b[108])^(a[56] & b[109])^(a[55] & b[110])^(a[54] & b[111])^(a[53] & b[112])^(a[52] & b[113])^(a[51] & b[114])^(a[50] & b[115])^(a[49] & b[116])^(a[48] & b[117])^(a[47] & b[118])^(a[46] & b[119])^(a[45] & b[120])^(a[44] & b[121])^(a[43] & b[122])^(a[42] & b[123])^(a[41] & b[124])^(a[40] & b[125])^(a[39] & b[126])^(a[38] & b[127])^(a[37] & b[128])^(a[36] & b[129])^(a[35] & b[130])^(a[34] & b[131])^(a[33] & b[132])^(a[32] & b[133])^(a[31] & b[134])^(a[30] & b[135])^(a[29] & b[136])^(a[28] & b[137])^(a[27] & b[138])^(a[26] & b[139])^(a[25] & b[140])^(a[24] & b[141])^(a[23] & b[142])^(a[22] & b[143])^(a[21] & b[144])^(a[20] & b[145])^(a[19] & b[146])^(a[18] & b[147])^(a[17] & b[148])^(a[16] & b[149])^(a[15] & b[150])^(a[14] & b[151])^(a[13] & b[152])^(a[12] & b[153])^(a[11] & b[154])^(a[10] & b[155])^(a[9] & b[156])^(a[8] & b[157])^(a[7] & b[158])^(a[6] & b[159])^(a[5] & b[160])^(a[4] & b[161])^(a[3] & b[162])^(a[2] & b[163])^(a[1] & b[164])^(a[0] & b[165]);
assign y[166] = (a[166] & b[0])^(a[165] & b[1])^(a[164] & b[2])^(a[163] & b[3])^(a[162] & b[4])^(a[161] & b[5])^(a[160] & b[6])^(a[159] & b[7])^(a[158] & b[8])^(a[157] & b[9])^(a[156] & b[10])^(a[155] & b[11])^(a[154] & b[12])^(a[153] & b[13])^(a[152] & b[14])^(a[151] & b[15])^(a[150] & b[16])^(a[149] & b[17])^(a[148] & b[18])^(a[147] & b[19])^(a[146] & b[20])^(a[145] & b[21])^(a[144] & b[22])^(a[143] & b[23])^(a[142] & b[24])^(a[141] & b[25])^(a[140] & b[26])^(a[139] & b[27])^(a[138] & b[28])^(a[137] & b[29])^(a[136] & b[30])^(a[135] & b[31])^(a[134] & b[32])^(a[133] & b[33])^(a[132] & b[34])^(a[131] & b[35])^(a[130] & b[36])^(a[129] & b[37])^(a[128] & b[38])^(a[127] & b[39])^(a[126] & b[40])^(a[125] & b[41])^(a[124] & b[42])^(a[123] & b[43])^(a[122] & b[44])^(a[121] & b[45])^(a[120] & b[46])^(a[119] & b[47])^(a[118] & b[48])^(a[117] & b[49])^(a[116] & b[50])^(a[115] & b[51])^(a[114] & b[52])^(a[113] & b[53])^(a[112] & b[54])^(a[111] & b[55])^(a[110] & b[56])^(a[109] & b[57])^(a[108] & b[58])^(a[107] & b[59])^(a[106] & b[60])^(a[105] & b[61])^(a[104] & b[62])^(a[103] & b[63])^(a[102] & b[64])^(a[101] & b[65])^(a[100] & b[66])^(a[99] & b[67])^(a[98] & b[68])^(a[97] & b[69])^(a[96] & b[70])^(a[95] & b[71])^(a[94] & b[72])^(a[93] & b[73])^(a[92] & b[74])^(a[91] & b[75])^(a[90] & b[76])^(a[89] & b[77])^(a[88] & b[78])^(a[87] & b[79])^(a[86] & b[80])^(a[85] & b[81])^(a[84] & b[82])^(a[83] & b[83])^(a[82] & b[84])^(a[81] & b[85])^(a[80] & b[86])^(a[79] & b[87])^(a[78] & b[88])^(a[77] & b[89])^(a[76] & b[90])^(a[75] & b[91])^(a[74] & b[92])^(a[73] & b[93])^(a[72] & b[94])^(a[71] & b[95])^(a[70] & b[96])^(a[69] & b[97])^(a[68] & b[98])^(a[67] & b[99])^(a[66] & b[100])^(a[65] & b[101])^(a[64] & b[102])^(a[63] & b[103])^(a[62] & b[104])^(a[61] & b[105])^(a[60] & b[106])^(a[59] & b[107])^(a[58] & b[108])^(a[57] & b[109])^(a[56] & b[110])^(a[55] & b[111])^(a[54] & b[112])^(a[53] & b[113])^(a[52] & b[114])^(a[51] & b[115])^(a[50] & b[116])^(a[49] & b[117])^(a[48] & b[118])^(a[47] & b[119])^(a[46] & b[120])^(a[45] & b[121])^(a[44] & b[122])^(a[43] & b[123])^(a[42] & b[124])^(a[41] & b[125])^(a[40] & b[126])^(a[39] & b[127])^(a[38] & b[128])^(a[37] & b[129])^(a[36] & b[130])^(a[35] & b[131])^(a[34] & b[132])^(a[33] & b[133])^(a[32] & b[134])^(a[31] & b[135])^(a[30] & b[136])^(a[29] & b[137])^(a[28] & b[138])^(a[27] & b[139])^(a[26] & b[140])^(a[25] & b[141])^(a[24] & b[142])^(a[23] & b[143])^(a[22] & b[144])^(a[21] & b[145])^(a[20] & b[146])^(a[19] & b[147])^(a[18] & b[148])^(a[17] & b[149])^(a[16] & b[150])^(a[15] & b[151])^(a[14] & b[152])^(a[13] & b[153])^(a[12] & b[154])^(a[11] & b[155])^(a[10] & b[156])^(a[9] & b[157])^(a[8] & b[158])^(a[7] & b[159])^(a[6] & b[160])^(a[5] & b[161])^(a[4] & b[162])^(a[3] & b[163])^(a[2] & b[164])^(a[1] & b[165])^(a[0] & b[166]);
assign y[167] = (a[167] & b[0])^(a[166] & b[1])^(a[165] & b[2])^(a[164] & b[3])^(a[163] & b[4])^(a[162] & b[5])^(a[161] & b[6])^(a[160] & b[7])^(a[159] & b[8])^(a[158] & b[9])^(a[157] & b[10])^(a[156] & b[11])^(a[155] & b[12])^(a[154] & b[13])^(a[153] & b[14])^(a[152] & b[15])^(a[151] & b[16])^(a[150] & b[17])^(a[149] & b[18])^(a[148] & b[19])^(a[147] & b[20])^(a[146] & b[21])^(a[145] & b[22])^(a[144] & b[23])^(a[143] & b[24])^(a[142] & b[25])^(a[141] & b[26])^(a[140] & b[27])^(a[139] & b[28])^(a[138] & b[29])^(a[137] & b[30])^(a[136] & b[31])^(a[135] & b[32])^(a[134] & b[33])^(a[133] & b[34])^(a[132] & b[35])^(a[131] & b[36])^(a[130] & b[37])^(a[129] & b[38])^(a[128] & b[39])^(a[127] & b[40])^(a[126] & b[41])^(a[125] & b[42])^(a[124] & b[43])^(a[123] & b[44])^(a[122] & b[45])^(a[121] & b[46])^(a[120] & b[47])^(a[119] & b[48])^(a[118] & b[49])^(a[117] & b[50])^(a[116] & b[51])^(a[115] & b[52])^(a[114] & b[53])^(a[113] & b[54])^(a[112] & b[55])^(a[111] & b[56])^(a[110] & b[57])^(a[109] & b[58])^(a[108] & b[59])^(a[107] & b[60])^(a[106] & b[61])^(a[105] & b[62])^(a[104] & b[63])^(a[103] & b[64])^(a[102] & b[65])^(a[101] & b[66])^(a[100] & b[67])^(a[99] & b[68])^(a[98] & b[69])^(a[97] & b[70])^(a[96] & b[71])^(a[95] & b[72])^(a[94] & b[73])^(a[93] & b[74])^(a[92] & b[75])^(a[91] & b[76])^(a[90] & b[77])^(a[89] & b[78])^(a[88] & b[79])^(a[87] & b[80])^(a[86] & b[81])^(a[85] & b[82])^(a[84] & b[83])^(a[83] & b[84])^(a[82] & b[85])^(a[81] & b[86])^(a[80] & b[87])^(a[79] & b[88])^(a[78] & b[89])^(a[77] & b[90])^(a[76] & b[91])^(a[75] & b[92])^(a[74] & b[93])^(a[73] & b[94])^(a[72] & b[95])^(a[71] & b[96])^(a[70] & b[97])^(a[69] & b[98])^(a[68] & b[99])^(a[67] & b[100])^(a[66] & b[101])^(a[65] & b[102])^(a[64] & b[103])^(a[63] & b[104])^(a[62] & b[105])^(a[61] & b[106])^(a[60] & b[107])^(a[59] & b[108])^(a[58] & b[109])^(a[57] & b[110])^(a[56] & b[111])^(a[55] & b[112])^(a[54] & b[113])^(a[53] & b[114])^(a[52] & b[115])^(a[51] & b[116])^(a[50] & b[117])^(a[49] & b[118])^(a[48] & b[119])^(a[47] & b[120])^(a[46] & b[121])^(a[45] & b[122])^(a[44] & b[123])^(a[43] & b[124])^(a[42] & b[125])^(a[41] & b[126])^(a[40] & b[127])^(a[39] & b[128])^(a[38] & b[129])^(a[37] & b[130])^(a[36] & b[131])^(a[35] & b[132])^(a[34] & b[133])^(a[33] & b[134])^(a[32] & b[135])^(a[31] & b[136])^(a[30] & b[137])^(a[29] & b[138])^(a[28] & b[139])^(a[27] & b[140])^(a[26] & b[141])^(a[25] & b[142])^(a[24] & b[143])^(a[23] & b[144])^(a[22] & b[145])^(a[21] & b[146])^(a[20] & b[147])^(a[19] & b[148])^(a[18] & b[149])^(a[17] & b[150])^(a[16] & b[151])^(a[15] & b[152])^(a[14] & b[153])^(a[13] & b[154])^(a[12] & b[155])^(a[11] & b[156])^(a[10] & b[157])^(a[9] & b[158])^(a[8] & b[159])^(a[7] & b[160])^(a[6] & b[161])^(a[5] & b[162])^(a[4] & b[163])^(a[3] & b[164])^(a[2] & b[165])^(a[1] & b[166])^(a[0] & b[167]);
assign y[168] = (a[168] & b[0])^(a[167] & b[1])^(a[166] & b[2])^(a[165] & b[3])^(a[164] & b[4])^(a[163] & b[5])^(a[162] & b[6])^(a[161] & b[7])^(a[160] & b[8])^(a[159] & b[9])^(a[158] & b[10])^(a[157] & b[11])^(a[156] & b[12])^(a[155] & b[13])^(a[154] & b[14])^(a[153] & b[15])^(a[152] & b[16])^(a[151] & b[17])^(a[150] & b[18])^(a[149] & b[19])^(a[148] & b[20])^(a[147] & b[21])^(a[146] & b[22])^(a[145] & b[23])^(a[144] & b[24])^(a[143] & b[25])^(a[142] & b[26])^(a[141] & b[27])^(a[140] & b[28])^(a[139] & b[29])^(a[138] & b[30])^(a[137] & b[31])^(a[136] & b[32])^(a[135] & b[33])^(a[134] & b[34])^(a[133] & b[35])^(a[132] & b[36])^(a[131] & b[37])^(a[130] & b[38])^(a[129] & b[39])^(a[128] & b[40])^(a[127] & b[41])^(a[126] & b[42])^(a[125] & b[43])^(a[124] & b[44])^(a[123] & b[45])^(a[122] & b[46])^(a[121] & b[47])^(a[120] & b[48])^(a[119] & b[49])^(a[118] & b[50])^(a[117] & b[51])^(a[116] & b[52])^(a[115] & b[53])^(a[114] & b[54])^(a[113] & b[55])^(a[112] & b[56])^(a[111] & b[57])^(a[110] & b[58])^(a[109] & b[59])^(a[108] & b[60])^(a[107] & b[61])^(a[106] & b[62])^(a[105] & b[63])^(a[104] & b[64])^(a[103] & b[65])^(a[102] & b[66])^(a[101] & b[67])^(a[100] & b[68])^(a[99] & b[69])^(a[98] & b[70])^(a[97] & b[71])^(a[96] & b[72])^(a[95] & b[73])^(a[94] & b[74])^(a[93] & b[75])^(a[92] & b[76])^(a[91] & b[77])^(a[90] & b[78])^(a[89] & b[79])^(a[88] & b[80])^(a[87] & b[81])^(a[86] & b[82])^(a[85] & b[83])^(a[84] & b[84])^(a[83] & b[85])^(a[82] & b[86])^(a[81] & b[87])^(a[80] & b[88])^(a[79] & b[89])^(a[78] & b[90])^(a[77] & b[91])^(a[76] & b[92])^(a[75] & b[93])^(a[74] & b[94])^(a[73] & b[95])^(a[72] & b[96])^(a[71] & b[97])^(a[70] & b[98])^(a[69] & b[99])^(a[68] & b[100])^(a[67] & b[101])^(a[66] & b[102])^(a[65] & b[103])^(a[64] & b[104])^(a[63] & b[105])^(a[62] & b[106])^(a[61] & b[107])^(a[60] & b[108])^(a[59] & b[109])^(a[58] & b[110])^(a[57] & b[111])^(a[56] & b[112])^(a[55] & b[113])^(a[54] & b[114])^(a[53] & b[115])^(a[52] & b[116])^(a[51] & b[117])^(a[50] & b[118])^(a[49] & b[119])^(a[48] & b[120])^(a[47] & b[121])^(a[46] & b[122])^(a[45] & b[123])^(a[44] & b[124])^(a[43] & b[125])^(a[42] & b[126])^(a[41] & b[127])^(a[40] & b[128])^(a[39] & b[129])^(a[38] & b[130])^(a[37] & b[131])^(a[36] & b[132])^(a[35] & b[133])^(a[34] & b[134])^(a[33] & b[135])^(a[32] & b[136])^(a[31] & b[137])^(a[30] & b[138])^(a[29] & b[139])^(a[28] & b[140])^(a[27] & b[141])^(a[26] & b[142])^(a[25] & b[143])^(a[24] & b[144])^(a[23] & b[145])^(a[22] & b[146])^(a[21] & b[147])^(a[20] & b[148])^(a[19] & b[149])^(a[18] & b[150])^(a[17] & b[151])^(a[16] & b[152])^(a[15] & b[153])^(a[14] & b[154])^(a[13] & b[155])^(a[12] & b[156])^(a[11] & b[157])^(a[10] & b[158])^(a[9] & b[159])^(a[8] & b[160])^(a[7] & b[161])^(a[6] & b[162])^(a[5] & b[163])^(a[4] & b[164])^(a[3] & b[165])^(a[2] & b[166])^(a[1] & b[167])^(a[0] & b[168]);
assign y[169] = (a[169] & b[0])^(a[168] & b[1])^(a[167] & b[2])^(a[166] & b[3])^(a[165] & b[4])^(a[164] & b[5])^(a[163] & b[6])^(a[162] & b[7])^(a[161] & b[8])^(a[160] & b[9])^(a[159] & b[10])^(a[158] & b[11])^(a[157] & b[12])^(a[156] & b[13])^(a[155] & b[14])^(a[154] & b[15])^(a[153] & b[16])^(a[152] & b[17])^(a[151] & b[18])^(a[150] & b[19])^(a[149] & b[20])^(a[148] & b[21])^(a[147] & b[22])^(a[146] & b[23])^(a[145] & b[24])^(a[144] & b[25])^(a[143] & b[26])^(a[142] & b[27])^(a[141] & b[28])^(a[140] & b[29])^(a[139] & b[30])^(a[138] & b[31])^(a[137] & b[32])^(a[136] & b[33])^(a[135] & b[34])^(a[134] & b[35])^(a[133] & b[36])^(a[132] & b[37])^(a[131] & b[38])^(a[130] & b[39])^(a[129] & b[40])^(a[128] & b[41])^(a[127] & b[42])^(a[126] & b[43])^(a[125] & b[44])^(a[124] & b[45])^(a[123] & b[46])^(a[122] & b[47])^(a[121] & b[48])^(a[120] & b[49])^(a[119] & b[50])^(a[118] & b[51])^(a[117] & b[52])^(a[116] & b[53])^(a[115] & b[54])^(a[114] & b[55])^(a[113] & b[56])^(a[112] & b[57])^(a[111] & b[58])^(a[110] & b[59])^(a[109] & b[60])^(a[108] & b[61])^(a[107] & b[62])^(a[106] & b[63])^(a[105] & b[64])^(a[104] & b[65])^(a[103] & b[66])^(a[102] & b[67])^(a[101] & b[68])^(a[100] & b[69])^(a[99] & b[70])^(a[98] & b[71])^(a[97] & b[72])^(a[96] & b[73])^(a[95] & b[74])^(a[94] & b[75])^(a[93] & b[76])^(a[92] & b[77])^(a[91] & b[78])^(a[90] & b[79])^(a[89] & b[80])^(a[88] & b[81])^(a[87] & b[82])^(a[86] & b[83])^(a[85] & b[84])^(a[84] & b[85])^(a[83] & b[86])^(a[82] & b[87])^(a[81] & b[88])^(a[80] & b[89])^(a[79] & b[90])^(a[78] & b[91])^(a[77] & b[92])^(a[76] & b[93])^(a[75] & b[94])^(a[74] & b[95])^(a[73] & b[96])^(a[72] & b[97])^(a[71] & b[98])^(a[70] & b[99])^(a[69] & b[100])^(a[68] & b[101])^(a[67] & b[102])^(a[66] & b[103])^(a[65] & b[104])^(a[64] & b[105])^(a[63] & b[106])^(a[62] & b[107])^(a[61] & b[108])^(a[60] & b[109])^(a[59] & b[110])^(a[58] & b[111])^(a[57] & b[112])^(a[56] & b[113])^(a[55] & b[114])^(a[54] & b[115])^(a[53] & b[116])^(a[52] & b[117])^(a[51] & b[118])^(a[50] & b[119])^(a[49] & b[120])^(a[48] & b[121])^(a[47] & b[122])^(a[46] & b[123])^(a[45] & b[124])^(a[44] & b[125])^(a[43] & b[126])^(a[42] & b[127])^(a[41] & b[128])^(a[40] & b[129])^(a[39] & b[130])^(a[38] & b[131])^(a[37] & b[132])^(a[36] & b[133])^(a[35] & b[134])^(a[34] & b[135])^(a[33] & b[136])^(a[32] & b[137])^(a[31] & b[138])^(a[30] & b[139])^(a[29] & b[140])^(a[28] & b[141])^(a[27] & b[142])^(a[26] & b[143])^(a[25] & b[144])^(a[24] & b[145])^(a[23] & b[146])^(a[22] & b[147])^(a[21] & b[148])^(a[20] & b[149])^(a[19] & b[150])^(a[18] & b[151])^(a[17] & b[152])^(a[16] & b[153])^(a[15] & b[154])^(a[14] & b[155])^(a[13] & b[156])^(a[12] & b[157])^(a[11] & b[158])^(a[10] & b[159])^(a[9] & b[160])^(a[8] & b[161])^(a[7] & b[162])^(a[6] & b[163])^(a[5] & b[164])^(a[4] & b[165])^(a[3] & b[166])^(a[2] & b[167])^(a[1] & b[168])^(a[0] & b[169]);
assign y[170] = (a[170] & b[0])^(a[169] & b[1])^(a[168] & b[2])^(a[167] & b[3])^(a[166] & b[4])^(a[165] & b[5])^(a[164] & b[6])^(a[163] & b[7])^(a[162] & b[8])^(a[161] & b[9])^(a[160] & b[10])^(a[159] & b[11])^(a[158] & b[12])^(a[157] & b[13])^(a[156] & b[14])^(a[155] & b[15])^(a[154] & b[16])^(a[153] & b[17])^(a[152] & b[18])^(a[151] & b[19])^(a[150] & b[20])^(a[149] & b[21])^(a[148] & b[22])^(a[147] & b[23])^(a[146] & b[24])^(a[145] & b[25])^(a[144] & b[26])^(a[143] & b[27])^(a[142] & b[28])^(a[141] & b[29])^(a[140] & b[30])^(a[139] & b[31])^(a[138] & b[32])^(a[137] & b[33])^(a[136] & b[34])^(a[135] & b[35])^(a[134] & b[36])^(a[133] & b[37])^(a[132] & b[38])^(a[131] & b[39])^(a[130] & b[40])^(a[129] & b[41])^(a[128] & b[42])^(a[127] & b[43])^(a[126] & b[44])^(a[125] & b[45])^(a[124] & b[46])^(a[123] & b[47])^(a[122] & b[48])^(a[121] & b[49])^(a[120] & b[50])^(a[119] & b[51])^(a[118] & b[52])^(a[117] & b[53])^(a[116] & b[54])^(a[115] & b[55])^(a[114] & b[56])^(a[113] & b[57])^(a[112] & b[58])^(a[111] & b[59])^(a[110] & b[60])^(a[109] & b[61])^(a[108] & b[62])^(a[107] & b[63])^(a[106] & b[64])^(a[105] & b[65])^(a[104] & b[66])^(a[103] & b[67])^(a[102] & b[68])^(a[101] & b[69])^(a[100] & b[70])^(a[99] & b[71])^(a[98] & b[72])^(a[97] & b[73])^(a[96] & b[74])^(a[95] & b[75])^(a[94] & b[76])^(a[93] & b[77])^(a[92] & b[78])^(a[91] & b[79])^(a[90] & b[80])^(a[89] & b[81])^(a[88] & b[82])^(a[87] & b[83])^(a[86] & b[84])^(a[85] & b[85])^(a[84] & b[86])^(a[83] & b[87])^(a[82] & b[88])^(a[81] & b[89])^(a[80] & b[90])^(a[79] & b[91])^(a[78] & b[92])^(a[77] & b[93])^(a[76] & b[94])^(a[75] & b[95])^(a[74] & b[96])^(a[73] & b[97])^(a[72] & b[98])^(a[71] & b[99])^(a[70] & b[100])^(a[69] & b[101])^(a[68] & b[102])^(a[67] & b[103])^(a[66] & b[104])^(a[65] & b[105])^(a[64] & b[106])^(a[63] & b[107])^(a[62] & b[108])^(a[61] & b[109])^(a[60] & b[110])^(a[59] & b[111])^(a[58] & b[112])^(a[57] & b[113])^(a[56] & b[114])^(a[55] & b[115])^(a[54] & b[116])^(a[53] & b[117])^(a[52] & b[118])^(a[51] & b[119])^(a[50] & b[120])^(a[49] & b[121])^(a[48] & b[122])^(a[47] & b[123])^(a[46] & b[124])^(a[45] & b[125])^(a[44] & b[126])^(a[43] & b[127])^(a[42] & b[128])^(a[41] & b[129])^(a[40] & b[130])^(a[39] & b[131])^(a[38] & b[132])^(a[37] & b[133])^(a[36] & b[134])^(a[35] & b[135])^(a[34] & b[136])^(a[33] & b[137])^(a[32] & b[138])^(a[31] & b[139])^(a[30] & b[140])^(a[29] & b[141])^(a[28] & b[142])^(a[27] & b[143])^(a[26] & b[144])^(a[25] & b[145])^(a[24] & b[146])^(a[23] & b[147])^(a[22] & b[148])^(a[21] & b[149])^(a[20] & b[150])^(a[19] & b[151])^(a[18] & b[152])^(a[17] & b[153])^(a[16] & b[154])^(a[15] & b[155])^(a[14] & b[156])^(a[13] & b[157])^(a[12] & b[158])^(a[11] & b[159])^(a[10] & b[160])^(a[9] & b[161])^(a[8] & b[162])^(a[7] & b[163])^(a[6] & b[164])^(a[5] & b[165])^(a[4] & b[166])^(a[3] & b[167])^(a[2] & b[168])^(a[1] & b[169])^(a[0] & b[170]);
assign y[171] = (a[171] & b[0])^(a[170] & b[1])^(a[169] & b[2])^(a[168] & b[3])^(a[167] & b[4])^(a[166] & b[5])^(a[165] & b[6])^(a[164] & b[7])^(a[163] & b[8])^(a[162] & b[9])^(a[161] & b[10])^(a[160] & b[11])^(a[159] & b[12])^(a[158] & b[13])^(a[157] & b[14])^(a[156] & b[15])^(a[155] & b[16])^(a[154] & b[17])^(a[153] & b[18])^(a[152] & b[19])^(a[151] & b[20])^(a[150] & b[21])^(a[149] & b[22])^(a[148] & b[23])^(a[147] & b[24])^(a[146] & b[25])^(a[145] & b[26])^(a[144] & b[27])^(a[143] & b[28])^(a[142] & b[29])^(a[141] & b[30])^(a[140] & b[31])^(a[139] & b[32])^(a[138] & b[33])^(a[137] & b[34])^(a[136] & b[35])^(a[135] & b[36])^(a[134] & b[37])^(a[133] & b[38])^(a[132] & b[39])^(a[131] & b[40])^(a[130] & b[41])^(a[129] & b[42])^(a[128] & b[43])^(a[127] & b[44])^(a[126] & b[45])^(a[125] & b[46])^(a[124] & b[47])^(a[123] & b[48])^(a[122] & b[49])^(a[121] & b[50])^(a[120] & b[51])^(a[119] & b[52])^(a[118] & b[53])^(a[117] & b[54])^(a[116] & b[55])^(a[115] & b[56])^(a[114] & b[57])^(a[113] & b[58])^(a[112] & b[59])^(a[111] & b[60])^(a[110] & b[61])^(a[109] & b[62])^(a[108] & b[63])^(a[107] & b[64])^(a[106] & b[65])^(a[105] & b[66])^(a[104] & b[67])^(a[103] & b[68])^(a[102] & b[69])^(a[101] & b[70])^(a[100] & b[71])^(a[99] & b[72])^(a[98] & b[73])^(a[97] & b[74])^(a[96] & b[75])^(a[95] & b[76])^(a[94] & b[77])^(a[93] & b[78])^(a[92] & b[79])^(a[91] & b[80])^(a[90] & b[81])^(a[89] & b[82])^(a[88] & b[83])^(a[87] & b[84])^(a[86] & b[85])^(a[85] & b[86])^(a[84] & b[87])^(a[83] & b[88])^(a[82] & b[89])^(a[81] & b[90])^(a[80] & b[91])^(a[79] & b[92])^(a[78] & b[93])^(a[77] & b[94])^(a[76] & b[95])^(a[75] & b[96])^(a[74] & b[97])^(a[73] & b[98])^(a[72] & b[99])^(a[71] & b[100])^(a[70] & b[101])^(a[69] & b[102])^(a[68] & b[103])^(a[67] & b[104])^(a[66] & b[105])^(a[65] & b[106])^(a[64] & b[107])^(a[63] & b[108])^(a[62] & b[109])^(a[61] & b[110])^(a[60] & b[111])^(a[59] & b[112])^(a[58] & b[113])^(a[57] & b[114])^(a[56] & b[115])^(a[55] & b[116])^(a[54] & b[117])^(a[53] & b[118])^(a[52] & b[119])^(a[51] & b[120])^(a[50] & b[121])^(a[49] & b[122])^(a[48] & b[123])^(a[47] & b[124])^(a[46] & b[125])^(a[45] & b[126])^(a[44] & b[127])^(a[43] & b[128])^(a[42] & b[129])^(a[41] & b[130])^(a[40] & b[131])^(a[39] & b[132])^(a[38] & b[133])^(a[37] & b[134])^(a[36] & b[135])^(a[35] & b[136])^(a[34] & b[137])^(a[33] & b[138])^(a[32] & b[139])^(a[31] & b[140])^(a[30] & b[141])^(a[29] & b[142])^(a[28] & b[143])^(a[27] & b[144])^(a[26] & b[145])^(a[25] & b[146])^(a[24] & b[147])^(a[23] & b[148])^(a[22] & b[149])^(a[21] & b[150])^(a[20] & b[151])^(a[19] & b[152])^(a[18] & b[153])^(a[17] & b[154])^(a[16] & b[155])^(a[15] & b[156])^(a[14] & b[157])^(a[13] & b[158])^(a[12] & b[159])^(a[11] & b[160])^(a[10] & b[161])^(a[9] & b[162])^(a[8] & b[163])^(a[7] & b[164])^(a[6] & b[165])^(a[5] & b[166])^(a[4] & b[167])^(a[3] & b[168])^(a[2] & b[169])^(a[1] & b[170])^(a[0] & b[171]);
assign y[172] = (a[172] & b[0])^(a[171] & b[1])^(a[170] & b[2])^(a[169] & b[3])^(a[168] & b[4])^(a[167] & b[5])^(a[166] & b[6])^(a[165] & b[7])^(a[164] & b[8])^(a[163] & b[9])^(a[162] & b[10])^(a[161] & b[11])^(a[160] & b[12])^(a[159] & b[13])^(a[158] & b[14])^(a[157] & b[15])^(a[156] & b[16])^(a[155] & b[17])^(a[154] & b[18])^(a[153] & b[19])^(a[152] & b[20])^(a[151] & b[21])^(a[150] & b[22])^(a[149] & b[23])^(a[148] & b[24])^(a[147] & b[25])^(a[146] & b[26])^(a[145] & b[27])^(a[144] & b[28])^(a[143] & b[29])^(a[142] & b[30])^(a[141] & b[31])^(a[140] & b[32])^(a[139] & b[33])^(a[138] & b[34])^(a[137] & b[35])^(a[136] & b[36])^(a[135] & b[37])^(a[134] & b[38])^(a[133] & b[39])^(a[132] & b[40])^(a[131] & b[41])^(a[130] & b[42])^(a[129] & b[43])^(a[128] & b[44])^(a[127] & b[45])^(a[126] & b[46])^(a[125] & b[47])^(a[124] & b[48])^(a[123] & b[49])^(a[122] & b[50])^(a[121] & b[51])^(a[120] & b[52])^(a[119] & b[53])^(a[118] & b[54])^(a[117] & b[55])^(a[116] & b[56])^(a[115] & b[57])^(a[114] & b[58])^(a[113] & b[59])^(a[112] & b[60])^(a[111] & b[61])^(a[110] & b[62])^(a[109] & b[63])^(a[108] & b[64])^(a[107] & b[65])^(a[106] & b[66])^(a[105] & b[67])^(a[104] & b[68])^(a[103] & b[69])^(a[102] & b[70])^(a[101] & b[71])^(a[100] & b[72])^(a[99] & b[73])^(a[98] & b[74])^(a[97] & b[75])^(a[96] & b[76])^(a[95] & b[77])^(a[94] & b[78])^(a[93] & b[79])^(a[92] & b[80])^(a[91] & b[81])^(a[90] & b[82])^(a[89] & b[83])^(a[88] & b[84])^(a[87] & b[85])^(a[86] & b[86])^(a[85] & b[87])^(a[84] & b[88])^(a[83] & b[89])^(a[82] & b[90])^(a[81] & b[91])^(a[80] & b[92])^(a[79] & b[93])^(a[78] & b[94])^(a[77] & b[95])^(a[76] & b[96])^(a[75] & b[97])^(a[74] & b[98])^(a[73] & b[99])^(a[72] & b[100])^(a[71] & b[101])^(a[70] & b[102])^(a[69] & b[103])^(a[68] & b[104])^(a[67] & b[105])^(a[66] & b[106])^(a[65] & b[107])^(a[64] & b[108])^(a[63] & b[109])^(a[62] & b[110])^(a[61] & b[111])^(a[60] & b[112])^(a[59] & b[113])^(a[58] & b[114])^(a[57] & b[115])^(a[56] & b[116])^(a[55] & b[117])^(a[54] & b[118])^(a[53] & b[119])^(a[52] & b[120])^(a[51] & b[121])^(a[50] & b[122])^(a[49] & b[123])^(a[48] & b[124])^(a[47] & b[125])^(a[46] & b[126])^(a[45] & b[127])^(a[44] & b[128])^(a[43] & b[129])^(a[42] & b[130])^(a[41] & b[131])^(a[40] & b[132])^(a[39] & b[133])^(a[38] & b[134])^(a[37] & b[135])^(a[36] & b[136])^(a[35] & b[137])^(a[34] & b[138])^(a[33] & b[139])^(a[32] & b[140])^(a[31] & b[141])^(a[30] & b[142])^(a[29] & b[143])^(a[28] & b[144])^(a[27] & b[145])^(a[26] & b[146])^(a[25] & b[147])^(a[24] & b[148])^(a[23] & b[149])^(a[22] & b[150])^(a[21] & b[151])^(a[20] & b[152])^(a[19] & b[153])^(a[18] & b[154])^(a[17] & b[155])^(a[16] & b[156])^(a[15] & b[157])^(a[14] & b[158])^(a[13] & b[159])^(a[12] & b[160])^(a[11] & b[161])^(a[10] & b[162])^(a[9] & b[163])^(a[8] & b[164])^(a[7] & b[165])^(a[6] & b[166])^(a[5] & b[167])^(a[4] & b[168])^(a[3] & b[169])^(a[2] & b[170])^(a[1] & b[171])^(a[0] & b[172]);
assign y[173] = (a[173] & b[0])^(a[172] & b[1])^(a[171] & b[2])^(a[170] & b[3])^(a[169] & b[4])^(a[168] & b[5])^(a[167] & b[6])^(a[166] & b[7])^(a[165] & b[8])^(a[164] & b[9])^(a[163] & b[10])^(a[162] & b[11])^(a[161] & b[12])^(a[160] & b[13])^(a[159] & b[14])^(a[158] & b[15])^(a[157] & b[16])^(a[156] & b[17])^(a[155] & b[18])^(a[154] & b[19])^(a[153] & b[20])^(a[152] & b[21])^(a[151] & b[22])^(a[150] & b[23])^(a[149] & b[24])^(a[148] & b[25])^(a[147] & b[26])^(a[146] & b[27])^(a[145] & b[28])^(a[144] & b[29])^(a[143] & b[30])^(a[142] & b[31])^(a[141] & b[32])^(a[140] & b[33])^(a[139] & b[34])^(a[138] & b[35])^(a[137] & b[36])^(a[136] & b[37])^(a[135] & b[38])^(a[134] & b[39])^(a[133] & b[40])^(a[132] & b[41])^(a[131] & b[42])^(a[130] & b[43])^(a[129] & b[44])^(a[128] & b[45])^(a[127] & b[46])^(a[126] & b[47])^(a[125] & b[48])^(a[124] & b[49])^(a[123] & b[50])^(a[122] & b[51])^(a[121] & b[52])^(a[120] & b[53])^(a[119] & b[54])^(a[118] & b[55])^(a[117] & b[56])^(a[116] & b[57])^(a[115] & b[58])^(a[114] & b[59])^(a[113] & b[60])^(a[112] & b[61])^(a[111] & b[62])^(a[110] & b[63])^(a[109] & b[64])^(a[108] & b[65])^(a[107] & b[66])^(a[106] & b[67])^(a[105] & b[68])^(a[104] & b[69])^(a[103] & b[70])^(a[102] & b[71])^(a[101] & b[72])^(a[100] & b[73])^(a[99] & b[74])^(a[98] & b[75])^(a[97] & b[76])^(a[96] & b[77])^(a[95] & b[78])^(a[94] & b[79])^(a[93] & b[80])^(a[92] & b[81])^(a[91] & b[82])^(a[90] & b[83])^(a[89] & b[84])^(a[88] & b[85])^(a[87] & b[86])^(a[86] & b[87])^(a[85] & b[88])^(a[84] & b[89])^(a[83] & b[90])^(a[82] & b[91])^(a[81] & b[92])^(a[80] & b[93])^(a[79] & b[94])^(a[78] & b[95])^(a[77] & b[96])^(a[76] & b[97])^(a[75] & b[98])^(a[74] & b[99])^(a[73] & b[100])^(a[72] & b[101])^(a[71] & b[102])^(a[70] & b[103])^(a[69] & b[104])^(a[68] & b[105])^(a[67] & b[106])^(a[66] & b[107])^(a[65] & b[108])^(a[64] & b[109])^(a[63] & b[110])^(a[62] & b[111])^(a[61] & b[112])^(a[60] & b[113])^(a[59] & b[114])^(a[58] & b[115])^(a[57] & b[116])^(a[56] & b[117])^(a[55] & b[118])^(a[54] & b[119])^(a[53] & b[120])^(a[52] & b[121])^(a[51] & b[122])^(a[50] & b[123])^(a[49] & b[124])^(a[48] & b[125])^(a[47] & b[126])^(a[46] & b[127])^(a[45] & b[128])^(a[44] & b[129])^(a[43] & b[130])^(a[42] & b[131])^(a[41] & b[132])^(a[40] & b[133])^(a[39] & b[134])^(a[38] & b[135])^(a[37] & b[136])^(a[36] & b[137])^(a[35] & b[138])^(a[34] & b[139])^(a[33] & b[140])^(a[32] & b[141])^(a[31] & b[142])^(a[30] & b[143])^(a[29] & b[144])^(a[28] & b[145])^(a[27] & b[146])^(a[26] & b[147])^(a[25] & b[148])^(a[24] & b[149])^(a[23] & b[150])^(a[22] & b[151])^(a[21] & b[152])^(a[20] & b[153])^(a[19] & b[154])^(a[18] & b[155])^(a[17] & b[156])^(a[16] & b[157])^(a[15] & b[158])^(a[14] & b[159])^(a[13] & b[160])^(a[12] & b[161])^(a[11] & b[162])^(a[10] & b[163])^(a[9] & b[164])^(a[8] & b[165])^(a[7] & b[166])^(a[6] & b[167])^(a[5] & b[168])^(a[4] & b[169])^(a[3] & b[170])^(a[2] & b[171])^(a[1] & b[172])^(a[0] & b[173]);
assign y[174] = (a[174] & b[0])^(a[173] & b[1])^(a[172] & b[2])^(a[171] & b[3])^(a[170] & b[4])^(a[169] & b[5])^(a[168] & b[6])^(a[167] & b[7])^(a[166] & b[8])^(a[165] & b[9])^(a[164] & b[10])^(a[163] & b[11])^(a[162] & b[12])^(a[161] & b[13])^(a[160] & b[14])^(a[159] & b[15])^(a[158] & b[16])^(a[157] & b[17])^(a[156] & b[18])^(a[155] & b[19])^(a[154] & b[20])^(a[153] & b[21])^(a[152] & b[22])^(a[151] & b[23])^(a[150] & b[24])^(a[149] & b[25])^(a[148] & b[26])^(a[147] & b[27])^(a[146] & b[28])^(a[145] & b[29])^(a[144] & b[30])^(a[143] & b[31])^(a[142] & b[32])^(a[141] & b[33])^(a[140] & b[34])^(a[139] & b[35])^(a[138] & b[36])^(a[137] & b[37])^(a[136] & b[38])^(a[135] & b[39])^(a[134] & b[40])^(a[133] & b[41])^(a[132] & b[42])^(a[131] & b[43])^(a[130] & b[44])^(a[129] & b[45])^(a[128] & b[46])^(a[127] & b[47])^(a[126] & b[48])^(a[125] & b[49])^(a[124] & b[50])^(a[123] & b[51])^(a[122] & b[52])^(a[121] & b[53])^(a[120] & b[54])^(a[119] & b[55])^(a[118] & b[56])^(a[117] & b[57])^(a[116] & b[58])^(a[115] & b[59])^(a[114] & b[60])^(a[113] & b[61])^(a[112] & b[62])^(a[111] & b[63])^(a[110] & b[64])^(a[109] & b[65])^(a[108] & b[66])^(a[107] & b[67])^(a[106] & b[68])^(a[105] & b[69])^(a[104] & b[70])^(a[103] & b[71])^(a[102] & b[72])^(a[101] & b[73])^(a[100] & b[74])^(a[99] & b[75])^(a[98] & b[76])^(a[97] & b[77])^(a[96] & b[78])^(a[95] & b[79])^(a[94] & b[80])^(a[93] & b[81])^(a[92] & b[82])^(a[91] & b[83])^(a[90] & b[84])^(a[89] & b[85])^(a[88] & b[86])^(a[87] & b[87])^(a[86] & b[88])^(a[85] & b[89])^(a[84] & b[90])^(a[83] & b[91])^(a[82] & b[92])^(a[81] & b[93])^(a[80] & b[94])^(a[79] & b[95])^(a[78] & b[96])^(a[77] & b[97])^(a[76] & b[98])^(a[75] & b[99])^(a[74] & b[100])^(a[73] & b[101])^(a[72] & b[102])^(a[71] & b[103])^(a[70] & b[104])^(a[69] & b[105])^(a[68] & b[106])^(a[67] & b[107])^(a[66] & b[108])^(a[65] & b[109])^(a[64] & b[110])^(a[63] & b[111])^(a[62] & b[112])^(a[61] & b[113])^(a[60] & b[114])^(a[59] & b[115])^(a[58] & b[116])^(a[57] & b[117])^(a[56] & b[118])^(a[55] & b[119])^(a[54] & b[120])^(a[53] & b[121])^(a[52] & b[122])^(a[51] & b[123])^(a[50] & b[124])^(a[49] & b[125])^(a[48] & b[126])^(a[47] & b[127])^(a[46] & b[128])^(a[45] & b[129])^(a[44] & b[130])^(a[43] & b[131])^(a[42] & b[132])^(a[41] & b[133])^(a[40] & b[134])^(a[39] & b[135])^(a[38] & b[136])^(a[37] & b[137])^(a[36] & b[138])^(a[35] & b[139])^(a[34] & b[140])^(a[33] & b[141])^(a[32] & b[142])^(a[31] & b[143])^(a[30] & b[144])^(a[29] & b[145])^(a[28] & b[146])^(a[27] & b[147])^(a[26] & b[148])^(a[25] & b[149])^(a[24] & b[150])^(a[23] & b[151])^(a[22] & b[152])^(a[21] & b[153])^(a[20] & b[154])^(a[19] & b[155])^(a[18] & b[156])^(a[17] & b[157])^(a[16] & b[158])^(a[15] & b[159])^(a[14] & b[160])^(a[13] & b[161])^(a[12] & b[162])^(a[11] & b[163])^(a[10] & b[164])^(a[9] & b[165])^(a[8] & b[166])^(a[7] & b[167])^(a[6] & b[168])^(a[5] & b[169])^(a[4] & b[170])^(a[3] & b[171])^(a[2] & b[172])^(a[1] & b[173])^(a[0] & b[174]);
assign y[175] = (a[175] & b[0])^(a[174] & b[1])^(a[173] & b[2])^(a[172] & b[3])^(a[171] & b[4])^(a[170] & b[5])^(a[169] & b[6])^(a[168] & b[7])^(a[167] & b[8])^(a[166] & b[9])^(a[165] & b[10])^(a[164] & b[11])^(a[163] & b[12])^(a[162] & b[13])^(a[161] & b[14])^(a[160] & b[15])^(a[159] & b[16])^(a[158] & b[17])^(a[157] & b[18])^(a[156] & b[19])^(a[155] & b[20])^(a[154] & b[21])^(a[153] & b[22])^(a[152] & b[23])^(a[151] & b[24])^(a[150] & b[25])^(a[149] & b[26])^(a[148] & b[27])^(a[147] & b[28])^(a[146] & b[29])^(a[145] & b[30])^(a[144] & b[31])^(a[143] & b[32])^(a[142] & b[33])^(a[141] & b[34])^(a[140] & b[35])^(a[139] & b[36])^(a[138] & b[37])^(a[137] & b[38])^(a[136] & b[39])^(a[135] & b[40])^(a[134] & b[41])^(a[133] & b[42])^(a[132] & b[43])^(a[131] & b[44])^(a[130] & b[45])^(a[129] & b[46])^(a[128] & b[47])^(a[127] & b[48])^(a[126] & b[49])^(a[125] & b[50])^(a[124] & b[51])^(a[123] & b[52])^(a[122] & b[53])^(a[121] & b[54])^(a[120] & b[55])^(a[119] & b[56])^(a[118] & b[57])^(a[117] & b[58])^(a[116] & b[59])^(a[115] & b[60])^(a[114] & b[61])^(a[113] & b[62])^(a[112] & b[63])^(a[111] & b[64])^(a[110] & b[65])^(a[109] & b[66])^(a[108] & b[67])^(a[107] & b[68])^(a[106] & b[69])^(a[105] & b[70])^(a[104] & b[71])^(a[103] & b[72])^(a[102] & b[73])^(a[101] & b[74])^(a[100] & b[75])^(a[99] & b[76])^(a[98] & b[77])^(a[97] & b[78])^(a[96] & b[79])^(a[95] & b[80])^(a[94] & b[81])^(a[93] & b[82])^(a[92] & b[83])^(a[91] & b[84])^(a[90] & b[85])^(a[89] & b[86])^(a[88] & b[87])^(a[87] & b[88])^(a[86] & b[89])^(a[85] & b[90])^(a[84] & b[91])^(a[83] & b[92])^(a[82] & b[93])^(a[81] & b[94])^(a[80] & b[95])^(a[79] & b[96])^(a[78] & b[97])^(a[77] & b[98])^(a[76] & b[99])^(a[75] & b[100])^(a[74] & b[101])^(a[73] & b[102])^(a[72] & b[103])^(a[71] & b[104])^(a[70] & b[105])^(a[69] & b[106])^(a[68] & b[107])^(a[67] & b[108])^(a[66] & b[109])^(a[65] & b[110])^(a[64] & b[111])^(a[63] & b[112])^(a[62] & b[113])^(a[61] & b[114])^(a[60] & b[115])^(a[59] & b[116])^(a[58] & b[117])^(a[57] & b[118])^(a[56] & b[119])^(a[55] & b[120])^(a[54] & b[121])^(a[53] & b[122])^(a[52] & b[123])^(a[51] & b[124])^(a[50] & b[125])^(a[49] & b[126])^(a[48] & b[127])^(a[47] & b[128])^(a[46] & b[129])^(a[45] & b[130])^(a[44] & b[131])^(a[43] & b[132])^(a[42] & b[133])^(a[41] & b[134])^(a[40] & b[135])^(a[39] & b[136])^(a[38] & b[137])^(a[37] & b[138])^(a[36] & b[139])^(a[35] & b[140])^(a[34] & b[141])^(a[33] & b[142])^(a[32] & b[143])^(a[31] & b[144])^(a[30] & b[145])^(a[29] & b[146])^(a[28] & b[147])^(a[27] & b[148])^(a[26] & b[149])^(a[25] & b[150])^(a[24] & b[151])^(a[23] & b[152])^(a[22] & b[153])^(a[21] & b[154])^(a[20] & b[155])^(a[19] & b[156])^(a[18] & b[157])^(a[17] & b[158])^(a[16] & b[159])^(a[15] & b[160])^(a[14] & b[161])^(a[13] & b[162])^(a[12] & b[163])^(a[11] & b[164])^(a[10] & b[165])^(a[9] & b[166])^(a[8] & b[167])^(a[7] & b[168])^(a[6] & b[169])^(a[5] & b[170])^(a[4] & b[171])^(a[3] & b[172])^(a[2] & b[173])^(a[1] & b[174])^(a[0] & b[175]);
assign y[176] = (a[176] & b[0])^(a[175] & b[1])^(a[174] & b[2])^(a[173] & b[3])^(a[172] & b[4])^(a[171] & b[5])^(a[170] & b[6])^(a[169] & b[7])^(a[168] & b[8])^(a[167] & b[9])^(a[166] & b[10])^(a[165] & b[11])^(a[164] & b[12])^(a[163] & b[13])^(a[162] & b[14])^(a[161] & b[15])^(a[160] & b[16])^(a[159] & b[17])^(a[158] & b[18])^(a[157] & b[19])^(a[156] & b[20])^(a[155] & b[21])^(a[154] & b[22])^(a[153] & b[23])^(a[152] & b[24])^(a[151] & b[25])^(a[150] & b[26])^(a[149] & b[27])^(a[148] & b[28])^(a[147] & b[29])^(a[146] & b[30])^(a[145] & b[31])^(a[144] & b[32])^(a[143] & b[33])^(a[142] & b[34])^(a[141] & b[35])^(a[140] & b[36])^(a[139] & b[37])^(a[138] & b[38])^(a[137] & b[39])^(a[136] & b[40])^(a[135] & b[41])^(a[134] & b[42])^(a[133] & b[43])^(a[132] & b[44])^(a[131] & b[45])^(a[130] & b[46])^(a[129] & b[47])^(a[128] & b[48])^(a[127] & b[49])^(a[126] & b[50])^(a[125] & b[51])^(a[124] & b[52])^(a[123] & b[53])^(a[122] & b[54])^(a[121] & b[55])^(a[120] & b[56])^(a[119] & b[57])^(a[118] & b[58])^(a[117] & b[59])^(a[116] & b[60])^(a[115] & b[61])^(a[114] & b[62])^(a[113] & b[63])^(a[112] & b[64])^(a[111] & b[65])^(a[110] & b[66])^(a[109] & b[67])^(a[108] & b[68])^(a[107] & b[69])^(a[106] & b[70])^(a[105] & b[71])^(a[104] & b[72])^(a[103] & b[73])^(a[102] & b[74])^(a[101] & b[75])^(a[100] & b[76])^(a[99] & b[77])^(a[98] & b[78])^(a[97] & b[79])^(a[96] & b[80])^(a[95] & b[81])^(a[94] & b[82])^(a[93] & b[83])^(a[92] & b[84])^(a[91] & b[85])^(a[90] & b[86])^(a[89] & b[87])^(a[88] & b[88])^(a[87] & b[89])^(a[86] & b[90])^(a[85] & b[91])^(a[84] & b[92])^(a[83] & b[93])^(a[82] & b[94])^(a[81] & b[95])^(a[80] & b[96])^(a[79] & b[97])^(a[78] & b[98])^(a[77] & b[99])^(a[76] & b[100])^(a[75] & b[101])^(a[74] & b[102])^(a[73] & b[103])^(a[72] & b[104])^(a[71] & b[105])^(a[70] & b[106])^(a[69] & b[107])^(a[68] & b[108])^(a[67] & b[109])^(a[66] & b[110])^(a[65] & b[111])^(a[64] & b[112])^(a[63] & b[113])^(a[62] & b[114])^(a[61] & b[115])^(a[60] & b[116])^(a[59] & b[117])^(a[58] & b[118])^(a[57] & b[119])^(a[56] & b[120])^(a[55] & b[121])^(a[54] & b[122])^(a[53] & b[123])^(a[52] & b[124])^(a[51] & b[125])^(a[50] & b[126])^(a[49] & b[127])^(a[48] & b[128])^(a[47] & b[129])^(a[46] & b[130])^(a[45] & b[131])^(a[44] & b[132])^(a[43] & b[133])^(a[42] & b[134])^(a[41] & b[135])^(a[40] & b[136])^(a[39] & b[137])^(a[38] & b[138])^(a[37] & b[139])^(a[36] & b[140])^(a[35] & b[141])^(a[34] & b[142])^(a[33] & b[143])^(a[32] & b[144])^(a[31] & b[145])^(a[30] & b[146])^(a[29] & b[147])^(a[28] & b[148])^(a[27] & b[149])^(a[26] & b[150])^(a[25] & b[151])^(a[24] & b[152])^(a[23] & b[153])^(a[22] & b[154])^(a[21] & b[155])^(a[20] & b[156])^(a[19] & b[157])^(a[18] & b[158])^(a[17] & b[159])^(a[16] & b[160])^(a[15] & b[161])^(a[14] & b[162])^(a[13] & b[163])^(a[12] & b[164])^(a[11] & b[165])^(a[10] & b[166])^(a[9] & b[167])^(a[8] & b[168])^(a[7] & b[169])^(a[6] & b[170])^(a[5] & b[171])^(a[4] & b[172])^(a[3] & b[173])^(a[2] & b[174])^(a[1] & b[175])^(a[0] & b[176]);
assign y[177] = (a[177] & b[0])^(a[176] & b[1])^(a[175] & b[2])^(a[174] & b[3])^(a[173] & b[4])^(a[172] & b[5])^(a[171] & b[6])^(a[170] & b[7])^(a[169] & b[8])^(a[168] & b[9])^(a[167] & b[10])^(a[166] & b[11])^(a[165] & b[12])^(a[164] & b[13])^(a[163] & b[14])^(a[162] & b[15])^(a[161] & b[16])^(a[160] & b[17])^(a[159] & b[18])^(a[158] & b[19])^(a[157] & b[20])^(a[156] & b[21])^(a[155] & b[22])^(a[154] & b[23])^(a[153] & b[24])^(a[152] & b[25])^(a[151] & b[26])^(a[150] & b[27])^(a[149] & b[28])^(a[148] & b[29])^(a[147] & b[30])^(a[146] & b[31])^(a[145] & b[32])^(a[144] & b[33])^(a[143] & b[34])^(a[142] & b[35])^(a[141] & b[36])^(a[140] & b[37])^(a[139] & b[38])^(a[138] & b[39])^(a[137] & b[40])^(a[136] & b[41])^(a[135] & b[42])^(a[134] & b[43])^(a[133] & b[44])^(a[132] & b[45])^(a[131] & b[46])^(a[130] & b[47])^(a[129] & b[48])^(a[128] & b[49])^(a[127] & b[50])^(a[126] & b[51])^(a[125] & b[52])^(a[124] & b[53])^(a[123] & b[54])^(a[122] & b[55])^(a[121] & b[56])^(a[120] & b[57])^(a[119] & b[58])^(a[118] & b[59])^(a[117] & b[60])^(a[116] & b[61])^(a[115] & b[62])^(a[114] & b[63])^(a[113] & b[64])^(a[112] & b[65])^(a[111] & b[66])^(a[110] & b[67])^(a[109] & b[68])^(a[108] & b[69])^(a[107] & b[70])^(a[106] & b[71])^(a[105] & b[72])^(a[104] & b[73])^(a[103] & b[74])^(a[102] & b[75])^(a[101] & b[76])^(a[100] & b[77])^(a[99] & b[78])^(a[98] & b[79])^(a[97] & b[80])^(a[96] & b[81])^(a[95] & b[82])^(a[94] & b[83])^(a[93] & b[84])^(a[92] & b[85])^(a[91] & b[86])^(a[90] & b[87])^(a[89] & b[88])^(a[88] & b[89])^(a[87] & b[90])^(a[86] & b[91])^(a[85] & b[92])^(a[84] & b[93])^(a[83] & b[94])^(a[82] & b[95])^(a[81] & b[96])^(a[80] & b[97])^(a[79] & b[98])^(a[78] & b[99])^(a[77] & b[100])^(a[76] & b[101])^(a[75] & b[102])^(a[74] & b[103])^(a[73] & b[104])^(a[72] & b[105])^(a[71] & b[106])^(a[70] & b[107])^(a[69] & b[108])^(a[68] & b[109])^(a[67] & b[110])^(a[66] & b[111])^(a[65] & b[112])^(a[64] & b[113])^(a[63] & b[114])^(a[62] & b[115])^(a[61] & b[116])^(a[60] & b[117])^(a[59] & b[118])^(a[58] & b[119])^(a[57] & b[120])^(a[56] & b[121])^(a[55] & b[122])^(a[54] & b[123])^(a[53] & b[124])^(a[52] & b[125])^(a[51] & b[126])^(a[50] & b[127])^(a[49] & b[128])^(a[48] & b[129])^(a[47] & b[130])^(a[46] & b[131])^(a[45] & b[132])^(a[44] & b[133])^(a[43] & b[134])^(a[42] & b[135])^(a[41] & b[136])^(a[40] & b[137])^(a[39] & b[138])^(a[38] & b[139])^(a[37] & b[140])^(a[36] & b[141])^(a[35] & b[142])^(a[34] & b[143])^(a[33] & b[144])^(a[32] & b[145])^(a[31] & b[146])^(a[30] & b[147])^(a[29] & b[148])^(a[28] & b[149])^(a[27] & b[150])^(a[26] & b[151])^(a[25] & b[152])^(a[24] & b[153])^(a[23] & b[154])^(a[22] & b[155])^(a[21] & b[156])^(a[20] & b[157])^(a[19] & b[158])^(a[18] & b[159])^(a[17] & b[160])^(a[16] & b[161])^(a[15] & b[162])^(a[14] & b[163])^(a[13] & b[164])^(a[12] & b[165])^(a[11] & b[166])^(a[10] & b[167])^(a[9] & b[168])^(a[8] & b[169])^(a[7] & b[170])^(a[6] & b[171])^(a[5] & b[172])^(a[4] & b[173])^(a[3] & b[174])^(a[2] & b[175])^(a[1] & b[176])^(a[0] & b[177]);
assign y[178] = (a[178] & b[0])^(a[177] & b[1])^(a[176] & b[2])^(a[175] & b[3])^(a[174] & b[4])^(a[173] & b[5])^(a[172] & b[6])^(a[171] & b[7])^(a[170] & b[8])^(a[169] & b[9])^(a[168] & b[10])^(a[167] & b[11])^(a[166] & b[12])^(a[165] & b[13])^(a[164] & b[14])^(a[163] & b[15])^(a[162] & b[16])^(a[161] & b[17])^(a[160] & b[18])^(a[159] & b[19])^(a[158] & b[20])^(a[157] & b[21])^(a[156] & b[22])^(a[155] & b[23])^(a[154] & b[24])^(a[153] & b[25])^(a[152] & b[26])^(a[151] & b[27])^(a[150] & b[28])^(a[149] & b[29])^(a[148] & b[30])^(a[147] & b[31])^(a[146] & b[32])^(a[145] & b[33])^(a[144] & b[34])^(a[143] & b[35])^(a[142] & b[36])^(a[141] & b[37])^(a[140] & b[38])^(a[139] & b[39])^(a[138] & b[40])^(a[137] & b[41])^(a[136] & b[42])^(a[135] & b[43])^(a[134] & b[44])^(a[133] & b[45])^(a[132] & b[46])^(a[131] & b[47])^(a[130] & b[48])^(a[129] & b[49])^(a[128] & b[50])^(a[127] & b[51])^(a[126] & b[52])^(a[125] & b[53])^(a[124] & b[54])^(a[123] & b[55])^(a[122] & b[56])^(a[121] & b[57])^(a[120] & b[58])^(a[119] & b[59])^(a[118] & b[60])^(a[117] & b[61])^(a[116] & b[62])^(a[115] & b[63])^(a[114] & b[64])^(a[113] & b[65])^(a[112] & b[66])^(a[111] & b[67])^(a[110] & b[68])^(a[109] & b[69])^(a[108] & b[70])^(a[107] & b[71])^(a[106] & b[72])^(a[105] & b[73])^(a[104] & b[74])^(a[103] & b[75])^(a[102] & b[76])^(a[101] & b[77])^(a[100] & b[78])^(a[99] & b[79])^(a[98] & b[80])^(a[97] & b[81])^(a[96] & b[82])^(a[95] & b[83])^(a[94] & b[84])^(a[93] & b[85])^(a[92] & b[86])^(a[91] & b[87])^(a[90] & b[88])^(a[89] & b[89])^(a[88] & b[90])^(a[87] & b[91])^(a[86] & b[92])^(a[85] & b[93])^(a[84] & b[94])^(a[83] & b[95])^(a[82] & b[96])^(a[81] & b[97])^(a[80] & b[98])^(a[79] & b[99])^(a[78] & b[100])^(a[77] & b[101])^(a[76] & b[102])^(a[75] & b[103])^(a[74] & b[104])^(a[73] & b[105])^(a[72] & b[106])^(a[71] & b[107])^(a[70] & b[108])^(a[69] & b[109])^(a[68] & b[110])^(a[67] & b[111])^(a[66] & b[112])^(a[65] & b[113])^(a[64] & b[114])^(a[63] & b[115])^(a[62] & b[116])^(a[61] & b[117])^(a[60] & b[118])^(a[59] & b[119])^(a[58] & b[120])^(a[57] & b[121])^(a[56] & b[122])^(a[55] & b[123])^(a[54] & b[124])^(a[53] & b[125])^(a[52] & b[126])^(a[51] & b[127])^(a[50] & b[128])^(a[49] & b[129])^(a[48] & b[130])^(a[47] & b[131])^(a[46] & b[132])^(a[45] & b[133])^(a[44] & b[134])^(a[43] & b[135])^(a[42] & b[136])^(a[41] & b[137])^(a[40] & b[138])^(a[39] & b[139])^(a[38] & b[140])^(a[37] & b[141])^(a[36] & b[142])^(a[35] & b[143])^(a[34] & b[144])^(a[33] & b[145])^(a[32] & b[146])^(a[31] & b[147])^(a[30] & b[148])^(a[29] & b[149])^(a[28] & b[150])^(a[27] & b[151])^(a[26] & b[152])^(a[25] & b[153])^(a[24] & b[154])^(a[23] & b[155])^(a[22] & b[156])^(a[21] & b[157])^(a[20] & b[158])^(a[19] & b[159])^(a[18] & b[160])^(a[17] & b[161])^(a[16] & b[162])^(a[15] & b[163])^(a[14] & b[164])^(a[13] & b[165])^(a[12] & b[166])^(a[11] & b[167])^(a[10] & b[168])^(a[9] & b[169])^(a[8] & b[170])^(a[7] & b[171])^(a[6] & b[172])^(a[5] & b[173])^(a[4] & b[174])^(a[3] & b[175])^(a[2] & b[176])^(a[1] & b[177])^(a[0] & b[178]);
assign y[179] = (a[179] & b[0])^(a[178] & b[1])^(a[177] & b[2])^(a[176] & b[3])^(a[175] & b[4])^(a[174] & b[5])^(a[173] & b[6])^(a[172] & b[7])^(a[171] & b[8])^(a[170] & b[9])^(a[169] & b[10])^(a[168] & b[11])^(a[167] & b[12])^(a[166] & b[13])^(a[165] & b[14])^(a[164] & b[15])^(a[163] & b[16])^(a[162] & b[17])^(a[161] & b[18])^(a[160] & b[19])^(a[159] & b[20])^(a[158] & b[21])^(a[157] & b[22])^(a[156] & b[23])^(a[155] & b[24])^(a[154] & b[25])^(a[153] & b[26])^(a[152] & b[27])^(a[151] & b[28])^(a[150] & b[29])^(a[149] & b[30])^(a[148] & b[31])^(a[147] & b[32])^(a[146] & b[33])^(a[145] & b[34])^(a[144] & b[35])^(a[143] & b[36])^(a[142] & b[37])^(a[141] & b[38])^(a[140] & b[39])^(a[139] & b[40])^(a[138] & b[41])^(a[137] & b[42])^(a[136] & b[43])^(a[135] & b[44])^(a[134] & b[45])^(a[133] & b[46])^(a[132] & b[47])^(a[131] & b[48])^(a[130] & b[49])^(a[129] & b[50])^(a[128] & b[51])^(a[127] & b[52])^(a[126] & b[53])^(a[125] & b[54])^(a[124] & b[55])^(a[123] & b[56])^(a[122] & b[57])^(a[121] & b[58])^(a[120] & b[59])^(a[119] & b[60])^(a[118] & b[61])^(a[117] & b[62])^(a[116] & b[63])^(a[115] & b[64])^(a[114] & b[65])^(a[113] & b[66])^(a[112] & b[67])^(a[111] & b[68])^(a[110] & b[69])^(a[109] & b[70])^(a[108] & b[71])^(a[107] & b[72])^(a[106] & b[73])^(a[105] & b[74])^(a[104] & b[75])^(a[103] & b[76])^(a[102] & b[77])^(a[101] & b[78])^(a[100] & b[79])^(a[99] & b[80])^(a[98] & b[81])^(a[97] & b[82])^(a[96] & b[83])^(a[95] & b[84])^(a[94] & b[85])^(a[93] & b[86])^(a[92] & b[87])^(a[91] & b[88])^(a[90] & b[89])^(a[89] & b[90])^(a[88] & b[91])^(a[87] & b[92])^(a[86] & b[93])^(a[85] & b[94])^(a[84] & b[95])^(a[83] & b[96])^(a[82] & b[97])^(a[81] & b[98])^(a[80] & b[99])^(a[79] & b[100])^(a[78] & b[101])^(a[77] & b[102])^(a[76] & b[103])^(a[75] & b[104])^(a[74] & b[105])^(a[73] & b[106])^(a[72] & b[107])^(a[71] & b[108])^(a[70] & b[109])^(a[69] & b[110])^(a[68] & b[111])^(a[67] & b[112])^(a[66] & b[113])^(a[65] & b[114])^(a[64] & b[115])^(a[63] & b[116])^(a[62] & b[117])^(a[61] & b[118])^(a[60] & b[119])^(a[59] & b[120])^(a[58] & b[121])^(a[57] & b[122])^(a[56] & b[123])^(a[55] & b[124])^(a[54] & b[125])^(a[53] & b[126])^(a[52] & b[127])^(a[51] & b[128])^(a[50] & b[129])^(a[49] & b[130])^(a[48] & b[131])^(a[47] & b[132])^(a[46] & b[133])^(a[45] & b[134])^(a[44] & b[135])^(a[43] & b[136])^(a[42] & b[137])^(a[41] & b[138])^(a[40] & b[139])^(a[39] & b[140])^(a[38] & b[141])^(a[37] & b[142])^(a[36] & b[143])^(a[35] & b[144])^(a[34] & b[145])^(a[33] & b[146])^(a[32] & b[147])^(a[31] & b[148])^(a[30] & b[149])^(a[29] & b[150])^(a[28] & b[151])^(a[27] & b[152])^(a[26] & b[153])^(a[25] & b[154])^(a[24] & b[155])^(a[23] & b[156])^(a[22] & b[157])^(a[21] & b[158])^(a[20] & b[159])^(a[19] & b[160])^(a[18] & b[161])^(a[17] & b[162])^(a[16] & b[163])^(a[15] & b[164])^(a[14] & b[165])^(a[13] & b[166])^(a[12] & b[167])^(a[11] & b[168])^(a[10] & b[169])^(a[9] & b[170])^(a[8] & b[171])^(a[7] & b[172])^(a[6] & b[173])^(a[5] & b[174])^(a[4] & b[175])^(a[3] & b[176])^(a[2] & b[177])^(a[1] & b[178])^(a[0] & b[179]);
assign y[180] = (a[180] & b[0])^(a[179] & b[1])^(a[178] & b[2])^(a[177] & b[3])^(a[176] & b[4])^(a[175] & b[5])^(a[174] & b[6])^(a[173] & b[7])^(a[172] & b[8])^(a[171] & b[9])^(a[170] & b[10])^(a[169] & b[11])^(a[168] & b[12])^(a[167] & b[13])^(a[166] & b[14])^(a[165] & b[15])^(a[164] & b[16])^(a[163] & b[17])^(a[162] & b[18])^(a[161] & b[19])^(a[160] & b[20])^(a[159] & b[21])^(a[158] & b[22])^(a[157] & b[23])^(a[156] & b[24])^(a[155] & b[25])^(a[154] & b[26])^(a[153] & b[27])^(a[152] & b[28])^(a[151] & b[29])^(a[150] & b[30])^(a[149] & b[31])^(a[148] & b[32])^(a[147] & b[33])^(a[146] & b[34])^(a[145] & b[35])^(a[144] & b[36])^(a[143] & b[37])^(a[142] & b[38])^(a[141] & b[39])^(a[140] & b[40])^(a[139] & b[41])^(a[138] & b[42])^(a[137] & b[43])^(a[136] & b[44])^(a[135] & b[45])^(a[134] & b[46])^(a[133] & b[47])^(a[132] & b[48])^(a[131] & b[49])^(a[130] & b[50])^(a[129] & b[51])^(a[128] & b[52])^(a[127] & b[53])^(a[126] & b[54])^(a[125] & b[55])^(a[124] & b[56])^(a[123] & b[57])^(a[122] & b[58])^(a[121] & b[59])^(a[120] & b[60])^(a[119] & b[61])^(a[118] & b[62])^(a[117] & b[63])^(a[116] & b[64])^(a[115] & b[65])^(a[114] & b[66])^(a[113] & b[67])^(a[112] & b[68])^(a[111] & b[69])^(a[110] & b[70])^(a[109] & b[71])^(a[108] & b[72])^(a[107] & b[73])^(a[106] & b[74])^(a[105] & b[75])^(a[104] & b[76])^(a[103] & b[77])^(a[102] & b[78])^(a[101] & b[79])^(a[100] & b[80])^(a[99] & b[81])^(a[98] & b[82])^(a[97] & b[83])^(a[96] & b[84])^(a[95] & b[85])^(a[94] & b[86])^(a[93] & b[87])^(a[92] & b[88])^(a[91] & b[89])^(a[90] & b[90])^(a[89] & b[91])^(a[88] & b[92])^(a[87] & b[93])^(a[86] & b[94])^(a[85] & b[95])^(a[84] & b[96])^(a[83] & b[97])^(a[82] & b[98])^(a[81] & b[99])^(a[80] & b[100])^(a[79] & b[101])^(a[78] & b[102])^(a[77] & b[103])^(a[76] & b[104])^(a[75] & b[105])^(a[74] & b[106])^(a[73] & b[107])^(a[72] & b[108])^(a[71] & b[109])^(a[70] & b[110])^(a[69] & b[111])^(a[68] & b[112])^(a[67] & b[113])^(a[66] & b[114])^(a[65] & b[115])^(a[64] & b[116])^(a[63] & b[117])^(a[62] & b[118])^(a[61] & b[119])^(a[60] & b[120])^(a[59] & b[121])^(a[58] & b[122])^(a[57] & b[123])^(a[56] & b[124])^(a[55] & b[125])^(a[54] & b[126])^(a[53] & b[127])^(a[52] & b[128])^(a[51] & b[129])^(a[50] & b[130])^(a[49] & b[131])^(a[48] & b[132])^(a[47] & b[133])^(a[46] & b[134])^(a[45] & b[135])^(a[44] & b[136])^(a[43] & b[137])^(a[42] & b[138])^(a[41] & b[139])^(a[40] & b[140])^(a[39] & b[141])^(a[38] & b[142])^(a[37] & b[143])^(a[36] & b[144])^(a[35] & b[145])^(a[34] & b[146])^(a[33] & b[147])^(a[32] & b[148])^(a[31] & b[149])^(a[30] & b[150])^(a[29] & b[151])^(a[28] & b[152])^(a[27] & b[153])^(a[26] & b[154])^(a[25] & b[155])^(a[24] & b[156])^(a[23] & b[157])^(a[22] & b[158])^(a[21] & b[159])^(a[20] & b[160])^(a[19] & b[161])^(a[18] & b[162])^(a[17] & b[163])^(a[16] & b[164])^(a[15] & b[165])^(a[14] & b[166])^(a[13] & b[167])^(a[12] & b[168])^(a[11] & b[169])^(a[10] & b[170])^(a[9] & b[171])^(a[8] & b[172])^(a[7] & b[173])^(a[6] & b[174])^(a[5] & b[175])^(a[4] & b[176])^(a[3] & b[177])^(a[2] & b[178])^(a[1] & b[179])^(a[0] & b[180]);
assign y[181] = (a[181] & b[0])^(a[180] & b[1])^(a[179] & b[2])^(a[178] & b[3])^(a[177] & b[4])^(a[176] & b[5])^(a[175] & b[6])^(a[174] & b[7])^(a[173] & b[8])^(a[172] & b[9])^(a[171] & b[10])^(a[170] & b[11])^(a[169] & b[12])^(a[168] & b[13])^(a[167] & b[14])^(a[166] & b[15])^(a[165] & b[16])^(a[164] & b[17])^(a[163] & b[18])^(a[162] & b[19])^(a[161] & b[20])^(a[160] & b[21])^(a[159] & b[22])^(a[158] & b[23])^(a[157] & b[24])^(a[156] & b[25])^(a[155] & b[26])^(a[154] & b[27])^(a[153] & b[28])^(a[152] & b[29])^(a[151] & b[30])^(a[150] & b[31])^(a[149] & b[32])^(a[148] & b[33])^(a[147] & b[34])^(a[146] & b[35])^(a[145] & b[36])^(a[144] & b[37])^(a[143] & b[38])^(a[142] & b[39])^(a[141] & b[40])^(a[140] & b[41])^(a[139] & b[42])^(a[138] & b[43])^(a[137] & b[44])^(a[136] & b[45])^(a[135] & b[46])^(a[134] & b[47])^(a[133] & b[48])^(a[132] & b[49])^(a[131] & b[50])^(a[130] & b[51])^(a[129] & b[52])^(a[128] & b[53])^(a[127] & b[54])^(a[126] & b[55])^(a[125] & b[56])^(a[124] & b[57])^(a[123] & b[58])^(a[122] & b[59])^(a[121] & b[60])^(a[120] & b[61])^(a[119] & b[62])^(a[118] & b[63])^(a[117] & b[64])^(a[116] & b[65])^(a[115] & b[66])^(a[114] & b[67])^(a[113] & b[68])^(a[112] & b[69])^(a[111] & b[70])^(a[110] & b[71])^(a[109] & b[72])^(a[108] & b[73])^(a[107] & b[74])^(a[106] & b[75])^(a[105] & b[76])^(a[104] & b[77])^(a[103] & b[78])^(a[102] & b[79])^(a[101] & b[80])^(a[100] & b[81])^(a[99] & b[82])^(a[98] & b[83])^(a[97] & b[84])^(a[96] & b[85])^(a[95] & b[86])^(a[94] & b[87])^(a[93] & b[88])^(a[92] & b[89])^(a[91] & b[90])^(a[90] & b[91])^(a[89] & b[92])^(a[88] & b[93])^(a[87] & b[94])^(a[86] & b[95])^(a[85] & b[96])^(a[84] & b[97])^(a[83] & b[98])^(a[82] & b[99])^(a[81] & b[100])^(a[80] & b[101])^(a[79] & b[102])^(a[78] & b[103])^(a[77] & b[104])^(a[76] & b[105])^(a[75] & b[106])^(a[74] & b[107])^(a[73] & b[108])^(a[72] & b[109])^(a[71] & b[110])^(a[70] & b[111])^(a[69] & b[112])^(a[68] & b[113])^(a[67] & b[114])^(a[66] & b[115])^(a[65] & b[116])^(a[64] & b[117])^(a[63] & b[118])^(a[62] & b[119])^(a[61] & b[120])^(a[60] & b[121])^(a[59] & b[122])^(a[58] & b[123])^(a[57] & b[124])^(a[56] & b[125])^(a[55] & b[126])^(a[54] & b[127])^(a[53] & b[128])^(a[52] & b[129])^(a[51] & b[130])^(a[50] & b[131])^(a[49] & b[132])^(a[48] & b[133])^(a[47] & b[134])^(a[46] & b[135])^(a[45] & b[136])^(a[44] & b[137])^(a[43] & b[138])^(a[42] & b[139])^(a[41] & b[140])^(a[40] & b[141])^(a[39] & b[142])^(a[38] & b[143])^(a[37] & b[144])^(a[36] & b[145])^(a[35] & b[146])^(a[34] & b[147])^(a[33] & b[148])^(a[32] & b[149])^(a[31] & b[150])^(a[30] & b[151])^(a[29] & b[152])^(a[28] & b[153])^(a[27] & b[154])^(a[26] & b[155])^(a[25] & b[156])^(a[24] & b[157])^(a[23] & b[158])^(a[22] & b[159])^(a[21] & b[160])^(a[20] & b[161])^(a[19] & b[162])^(a[18] & b[163])^(a[17] & b[164])^(a[16] & b[165])^(a[15] & b[166])^(a[14] & b[167])^(a[13] & b[168])^(a[12] & b[169])^(a[11] & b[170])^(a[10] & b[171])^(a[9] & b[172])^(a[8] & b[173])^(a[7] & b[174])^(a[6] & b[175])^(a[5] & b[176])^(a[4] & b[177])^(a[3] & b[178])^(a[2] & b[179])^(a[1] & b[180])^(a[0] & b[181]);
assign y[182] = (a[182] & b[0])^(a[181] & b[1])^(a[180] & b[2])^(a[179] & b[3])^(a[178] & b[4])^(a[177] & b[5])^(a[176] & b[6])^(a[175] & b[7])^(a[174] & b[8])^(a[173] & b[9])^(a[172] & b[10])^(a[171] & b[11])^(a[170] & b[12])^(a[169] & b[13])^(a[168] & b[14])^(a[167] & b[15])^(a[166] & b[16])^(a[165] & b[17])^(a[164] & b[18])^(a[163] & b[19])^(a[162] & b[20])^(a[161] & b[21])^(a[160] & b[22])^(a[159] & b[23])^(a[158] & b[24])^(a[157] & b[25])^(a[156] & b[26])^(a[155] & b[27])^(a[154] & b[28])^(a[153] & b[29])^(a[152] & b[30])^(a[151] & b[31])^(a[150] & b[32])^(a[149] & b[33])^(a[148] & b[34])^(a[147] & b[35])^(a[146] & b[36])^(a[145] & b[37])^(a[144] & b[38])^(a[143] & b[39])^(a[142] & b[40])^(a[141] & b[41])^(a[140] & b[42])^(a[139] & b[43])^(a[138] & b[44])^(a[137] & b[45])^(a[136] & b[46])^(a[135] & b[47])^(a[134] & b[48])^(a[133] & b[49])^(a[132] & b[50])^(a[131] & b[51])^(a[130] & b[52])^(a[129] & b[53])^(a[128] & b[54])^(a[127] & b[55])^(a[126] & b[56])^(a[125] & b[57])^(a[124] & b[58])^(a[123] & b[59])^(a[122] & b[60])^(a[121] & b[61])^(a[120] & b[62])^(a[119] & b[63])^(a[118] & b[64])^(a[117] & b[65])^(a[116] & b[66])^(a[115] & b[67])^(a[114] & b[68])^(a[113] & b[69])^(a[112] & b[70])^(a[111] & b[71])^(a[110] & b[72])^(a[109] & b[73])^(a[108] & b[74])^(a[107] & b[75])^(a[106] & b[76])^(a[105] & b[77])^(a[104] & b[78])^(a[103] & b[79])^(a[102] & b[80])^(a[101] & b[81])^(a[100] & b[82])^(a[99] & b[83])^(a[98] & b[84])^(a[97] & b[85])^(a[96] & b[86])^(a[95] & b[87])^(a[94] & b[88])^(a[93] & b[89])^(a[92] & b[90])^(a[91] & b[91])^(a[90] & b[92])^(a[89] & b[93])^(a[88] & b[94])^(a[87] & b[95])^(a[86] & b[96])^(a[85] & b[97])^(a[84] & b[98])^(a[83] & b[99])^(a[82] & b[100])^(a[81] & b[101])^(a[80] & b[102])^(a[79] & b[103])^(a[78] & b[104])^(a[77] & b[105])^(a[76] & b[106])^(a[75] & b[107])^(a[74] & b[108])^(a[73] & b[109])^(a[72] & b[110])^(a[71] & b[111])^(a[70] & b[112])^(a[69] & b[113])^(a[68] & b[114])^(a[67] & b[115])^(a[66] & b[116])^(a[65] & b[117])^(a[64] & b[118])^(a[63] & b[119])^(a[62] & b[120])^(a[61] & b[121])^(a[60] & b[122])^(a[59] & b[123])^(a[58] & b[124])^(a[57] & b[125])^(a[56] & b[126])^(a[55] & b[127])^(a[54] & b[128])^(a[53] & b[129])^(a[52] & b[130])^(a[51] & b[131])^(a[50] & b[132])^(a[49] & b[133])^(a[48] & b[134])^(a[47] & b[135])^(a[46] & b[136])^(a[45] & b[137])^(a[44] & b[138])^(a[43] & b[139])^(a[42] & b[140])^(a[41] & b[141])^(a[40] & b[142])^(a[39] & b[143])^(a[38] & b[144])^(a[37] & b[145])^(a[36] & b[146])^(a[35] & b[147])^(a[34] & b[148])^(a[33] & b[149])^(a[32] & b[150])^(a[31] & b[151])^(a[30] & b[152])^(a[29] & b[153])^(a[28] & b[154])^(a[27] & b[155])^(a[26] & b[156])^(a[25] & b[157])^(a[24] & b[158])^(a[23] & b[159])^(a[22] & b[160])^(a[21] & b[161])^(a[20] & b[162])^(a[19] & b[163])^(a[18] & b[164])^(a[17] & b[165])^(a[16] & b[166])^(a[15] & b[167])^(a[14] & b[168])^(a[13] & b[169])^(a[12] & b[170])^(a[11] & b[171])^(a[10] & b[172])^(a[9] & b[173])^(a[8] & b[174])^(a[7] & b[175])^(a[6] & b[176])^(a[5] & b[177])^(a[4] & b[178])^(a[3] & b[179])^(a[2] & b[180])^(a[1] & b[181])^(a[0] & b[182]);
assign y[183] = (a[183] & b[0])^(a[182] & b[1])^(a[181] & b[2])^(a[180] & b[3])^(a[179] & b[4])^(a[178] & b[5])^(a[177] & b[6])^(a[176] & b[7])^(a[175] & b[8])^(a[174] & b[9])^(a[173] & b[10])^(a[172] & b[11])^(a[171] & b[12])^(a[170] & b[13])^(a[169] & b[14])^(a[168] & b[15])^(a[167] & b[16])^(a[166] & b[17])^(a[165] & b[18])^(a[164] & b[19])^(a[163] & b[20])^(a[162] & b[21])^(a[161] & b[22])^(a[160] & b[23])^(a[159] & b[24])^(a[158] & b[25])^(a[157] & b[26])^(a[156] & b[27])^(a[155] & b[28])^(a[154] & b[29])^(a[153] & b[30])^(a[152] & b[31])^(a[151] & b[32])^(a[150] & b[33])^(a[149] & b[34])^(a[148] & b[35])^(a[147] & b[36])^(a[146] & b[37])^(a[145] & b[38])^(a[144] & b[39])^(a[143] & b[40])^(a[142] & b[41])^(a[141] & b[42])^(a[140] & b[43])^(a[139] & b[44])^(a[138] & b[45])^(a[137] & b[46])^(a[136] & b[47])^(a[135] & b[48])^(a[134] & b[49])^(a[133] & b[50])^(a[132] & b[51])^(a[131] & b[52])^(a[130] & b[53])^(a[129] & b[54])^(a[128] & b[55])^(a[127] & b[56])^(a[126] & b[57])^(a[125] & b[58])^(a[124] & b[59])^(a[123] & b[60])^(a[122] & b[61])^(a[121] & b[62])^(a[120] & b[63])^(a[119] & b[64])^(a[118] & b[65])^(a[117] & b[66])^(a[116] & b[67])^(a[115] & b[68])^(a[114] & b[69])^(a[113] & b[70])^(a[112] & b[71])^(a[111] & b[72])^(a[110] & b[73])^(a[109] & b[74])^(a[108] & b[75])^(a[107] & b[76])^(a[106] & b[77])^(a[105] & b[78])^(a[104] & b[79])^(a[103] & b[80])^(a[102] & b[81])^(a[101] & b[82])^(a[100] & b[83])^(a[99] & b[84])^(a[98] & b[85])^(a[97] & b[86])^(a[96] & b[87])^(a[95] & b[88])^(a[94] & b[89])^(a[93] & b[90])^(a[92] & b[91])^(a[91] & b[92])^(a[90] & b[93])^(a[89] & b[94])^(a[88] & b[95])^(a[87] & b[96])^(a[86] & b[97])^(a[85] & b[98])^(a[84] & b[99])^(a[83] & b[100])^(a[82] & b[101])^(a[81] & b[102])^(a[80] & b[103])^(a[79] & b[104])^(a[78] & b[105])^(a[77] & b[106])^(a[76] & b[107])^(a[75] & b[108])^(a[74] & b[109])^(a[73] & b[110])^(a[72] & b[111])^(a[71] & b[112])^(a[70] & b[113])^(a[69] & b[114])^(a[68] & b[115])^(a[67] & b[116])^(a[66] & b[117])^(a[65] & b[118])^(a[64] & b[119])^(a[63] & b[120])^(a[62] & b[121])^(a[61] & b[122])^(a[60] & b[123])^(a[59] & b[124])^(a[58] & b[125])^(a[57] & b[126])^(a[56] & b[127])^(a[55] & b[128])^(a[54] & b[129])^(a[53] & b[130])^(a[52] & b[131])^(a[51] & b[132])^(a[50] & b[133])^(a[49] & b[134])^(a[48] & b[135])^(a[47] & b[136])^(a[46] & b[137])^(a[45] & b[138])^(a[44] & b[139])^(a[43] & b[140])^(a[42] & b[141])^(a[41] & b[142])^(a[40] & b[143])^(a[39] & b[144])^(a[38] & b[145])^(a[37] & b[146])^(a[36] & b[147])^(a[35] & b[148])^(a[34] & b[149])^(a[33] & b[150])^(a[32] & b[151])^(a[31] & b[152])^(a[30] & b[153])^(a[29] & b[154])^(a[28] & b[155])^(a[27] & b[156])^(a[26] & b[157])^(a[25] & b[158])^(a[24] & b[159])^(a[23] & b[160])^(a[22] & b[161])^(a[21] & b[162])^(a[20] & b[163])^(a[19] & b[164])^(a[18] & b[165])^(a[17] & b[166])^(a[16] & b[167])^(a[15] & b[168])^(a[14] & b[169])^(a[13] & b[170])^(a[12] & b[171])^(a[11] & b[172])^(a[10] & b[173])^(a[9] & b[174])^(a[8] & b[175])^(a[7] & b[176])^(a[6] & b[177])^(a[5] & b[178])^(a[4] & b[179])^(a[3] & b[180])^(a[2] & b[181])^(a[1] & b[182])^(a[0] & b[183]);
assign y[184] = (a[184] & b[0])^(a[183] & b[1])^(a[182] & b[2])^(a[181] & b[3])^(a[180] & b[4])^(a[179] & b[5])^(a[178] & b[6])^(a[177] & b[7])^(a[176] & b[8])^(a[175] & b[9])^(a[174] & b[10])^(a[173] & b[11])^(a[172] & b[12])^(a[171] & b[13])^(a[170] & b[14])^(a[169] & b[15])^(a[168] & b[16])^(a[167] & b[17])^(a[166] & b[18])^(a[165] & b[19])^(a[164] & b[20])^(a[163] & b[21])^(a[162] & b[22])^(a[161] & b[23])^(a[160] & b[24])^(a[159] & b[25])^(a[158] & b[26])^(a[157] & b[27])^(a[156] & b[28])^(a[155] & b[29])^(a[154] & b[30])^(a[153] & b[31])^(a[152] & b[32])^(a[151] & b[33])^(a[150] & b[34])^(a[149] & b[35])^(a[148] & b[36])^(a[147] & b[37])^(a[146] & b[38])^(a[145] & b[39])^(a[144] & b[40])^(a[143] & b[41])^(a[142] & b[42])^(a[141] & b[43])^(a[140] & b[44])^(a[139] & b[45])^(a[138] & b[46])^(a[137] & b[47])^(a[136] & b[48])^(a[135] & b[49])^(a[134] & b[50])^(a[133] & b[51])^(a[132] & b[52])^(a[131] & b[53])^(a[130] & b[54])^(a[129] & b[55])^(a[128] & b[56])^(a[127] & b[57])^(a[126] & b[58])^(a[125] & b[59])^(a[124] & b[60])^(a[123] & b[61])^(a[122] & b[62])^(a[121] & b[63])^(a[120] & b[64])^(a[119] & b[65])^(a[118] & b[66])^(a[117] & b[67])^(a[116] & b[68])^(a[115] & b[69])^(a[114] & b[70])^(a[113] & b[71])^(a[112] & b[72])^(a[111] & b[73])^(a[110] & b[74])^(a[109] & b[75])^(a[108] & b[76])^(a[107] & b[77])^(a[106] & b[78])^(a[105] & b[79])^(a[104] & b[80])^(a[103] & b[81])^(a[102] & b[82])^(a[101] & b[83])^(a[100] & b[84])^(a[99] & b[85])^(a[98] & b[86])^(a[97] & b[87])^(a[96] & b[88])^(a[95] & b[89])^(a[94] & b[90])^(a[93] & b[91])^(a[92] & b[92])^(a[91] & b[93])^(a[90] & b[94])^(a[89] & b[95])^(a[88] & b[96])^(a[87] & b[97])^(a[86] & b[98])^(a[85] & b[99])^(a[84] & b[100])^(a[83] & b[101])^(a[82] & b[102])^(a[81] & b[103])^(a[80] & b[104])^(a[79] & b[105])^(a[78] & b[106])^(a[77] & b[107])^(a[76] & b[108])^(a[75] & b[109])^(a[74] & b[110])^(a[73] & b[111])^(a[72] & b[112])^(a[71] & b[113])^(a[70] & b[114])^(a[69] & b[115])^(a[68] & b[116])^(a[67] & b[117])^(a[66] & b[118])^(a[65] & b[119])^(a[64] & b[120])^(a[63] & b[121])^(a[62] & b[122])^(a[61] & b[123])^(a[60] & b[124])^(a[59] & b[125])^(a[58] & b[126])^(a[57] & b[127])^(a[56] & b[128])^(a[55] & b[129])^(a[54] & b[130])^(a[53] & b[131])^(a[52] & b[132])^(a[51] & b[133])^(a[50] & b[134])^(a[49] & b[135])^(a[48] & b[136])^(a[47] & b[137])^(a[46] & b[138])^(a[45] & b[139])^(a[44] & b[140])^(a[43] & b[141])^(a[42] & b[142])^(a[41] & b[143])^(a[40] & b[144])^(a[39] & b[145])^(a[38] & b[146])^(a[37] & b[147])^(a[36] & b[148])^(a[35] & b[149])^(a[34] & b[150])^(a[33] & b[151])^(a[32] & b[152])^(a[31] & b[153])^(a[30] & b[154])^(a[29] & b[155])^(a[28] & b[156])^(a[27] & b[157])^(a[26] & b[158])^(a[25] & b[159])^(a[24] & b[160])^(a[23] & b[161])^(a[22] & b[162])^(a[21] & b[163])^(a[20] & b[164])^(a[19] & b[165])^(a[18] & b[166])^(a[17] & b[167])^(a[16] & b[168])^(a[15] & b[169])^(a[14] & b[170])^(a[13] & b[171])^(a[12] & b[172])^(a[11] & b[173])^(a[10] & b[174])^(a[9] & b[175])^(a[8] & b[176])^(a[7] & b[177])^(a[6] & b[178])^(a[5] & b[179])^(a[4] & b[180])^(a[3] & b[181])^(a[2] & b[182])^(a[1] & b[183])^(a[0] & b[184]);
assign y[185] = (a[185] & b[0])^(a[184] & b[1])^(a[183] & b[2])^(a[182] & b[3])^(a[181] & b[4])^(a[180] & b[5])^(a[179] & b[6])^(a[178] & b[7])^(a[177] & b[8])^(a[176] & b[9])^(a[175] & b[10])^(a[174] & b[11])^(a[173] & b[12])^(a[172] & b[13])^(a[171] & b[14])^(a[170] & b[15])^(a[169] & b[16])^(a[168] & b[17])^(a[167] & b[18])^(a[166] & b[19])^(a[165] & b[20])^(a[164] & b[21])^(a[163] & b[22])^(a[162] & b[23])^(a[161] & b[24])^(a[160] & b[25])^(a[159] & b[26])^(a[158] & b[27])^(a[157] & b[28])^(a[156] & b[29])^(a[155] & b[30])^(a[154] & b[31])^(a[153] & b[32])^(a[152] & b[33])^(a[151] & b[34])^(a[150] & b[35])^(a[149] & b[36])^(a[148] & b[37])^(a[147] & b[38])^(a[146] & b[39])^(a[145] & b[40])^(a[144] & b[41])^(a[143] & b[42])^(a[142] & b[43])^(a[141] & b[44])^(a[140] & b[45])^(a[139] & b[46])^(a[138] & b[47])^(a[137] & b[48])^(a[136] & b[49])^(a[135] & b[50])^(a[134] & b[51])^(a[133] & b[52])^(a[132] & b[53])^(a[131] & b[54])^(a[130] & b[55])^(a[129] & b[56])^(a[128] & b[57])^(a[127] & b[58])^(a[126] & b[59])^(a[125] & b[60])^(a[124] & b[61])^(a[123] & b[62])^(a[122] & b[63])^(a[121] & b[64])^(a[120] & b[65])^(a[119] & b[66])^(a[118] & b[67])^(a[117] & b[68])^(a[116] & b[69])^(a[115] & b[70])^(a[114] & b[71])^(a[113] & b[72])^(a[112] & b[73])^(a[111] & b[74])^(a[110] & b[75])^(a[109] & b[76])^(a[108] & b[77])^(a[107] & b[78])^(a[106] & b[79])^(a[105] & b[80])^(a[104] & b[81])^(a[103] & b[82])^(a[102] & b[83])^(a[101] & b[84])^(a[100] & b[85])^(a[99] & b[86])^(a[98] & b[87])^(a[97] & b[88])^(a[96] & b[89])^(a[95] & b[90])^(a[94] & b[91])^(a[93] & b[92])^(a[92] & b[93])^(a[91] & b[94])^(a[90] & b[95])^(a[89] & b[96])^(a[88] & b[97])^(a[87] & b[98])^(a[86] & b[99])^(a[85] & b[100])^(a[84] & b[101])^(a[83] & b[102])^(a[82] & b[103])^(a[81] & b[104])^(a[80] & b[105])^(a[79] & b[106])^(a[78] & b[107])^(a[77] & b[108])^(a[76] & b[109])^(a[75] & b[110])^(a[74] & b[111])^(a[73] & b[112])^(a[72] & b[113])^(a[71] & b[114])^(a[70] & b[115])^(a[69] & b[116])^(a[68] & b[117])^(a[67] & b[118])^(a[66] & b[119])^(a[65] & b[120])^(a[64] & b[121])^(a[63] & b[122])^(a[62] & b[123])^(a[61] & b[124])^(a[60] & b[125])^(a[59] & b[126])^(a[58] & b[127])^(a[57] & b[128])^(a[56] & b[129])^(a[55] & b[130])^(a[54] & b[131])^(a[53] & b[132])^(a[52] & b[133])^(a[51] & b[134])^(a[50] & b[135])^(a[49] & b[136])^(a[48] & b[137])^(a[47] & b[138])^(a[46] & b[139])^(a[45] & b[140])^(a[44] & b[141])^(a[43] & b[142])^(a[42] & b[143])^(a[41] & b[144])^(a[40] & b[145])^(a[39] & b[146])^(a[38] & b[147])^(a[37] & b[148])^(a[36] & b[149])^(a[35] & b[150])^(a[34] & b[151])^(a[33] & b[152])^(a[32] & b[153])^(a[31] & b[154])^(a[30] & b[155])^(a[29] & b[156])^(a[28] & b[157])^(a[27] & b[158])^(a[26] & b[159])^(a[25] & b[160])^(a[24] & b[161])^(a[23] & b[162])^(a[22] & b[163])^(a[21] & b[164])^(a[20] & b[165])^(a[19] & b[166])^(a[18] & b[167])^(a[17] & b[168])^(a[16] & b[169])^(a[15] & b[170])^(a[14] & b[171])^(a[13] & b[172])^(a[12] & b[173])^(a[11] & b[174])^(a[10] & b[175])^(a[9] & b[176])^(a[8] & b[177])^(a[7] & b[178])^(a[6] & b[179])^(a[5] & b[180])^(a[4] & b[181])^(a[3] & b[182])^(a[2] & b[183])^(a[1] & b[184])^(a[0] & b[185]);
assign y[186] = (a[186] & b[0])^(a[185] & b[1])^(a[184] & b[2])^(a[183] & b[3])^(a[182] & b[4])^(a[181] & b[5])^(a[180] & b[6])^(a[179] & b[7])^(a[178] & b[8])^(a[177] & b[9])^(a[176] & b[10])^(a[175] & b[11])^(a[174] & b[12])^(a[173] & b[13])^(a[172] & b[14])^(a[171] & b[15])^(a[170] & b[16])^(a[169] & b[17])^(a[168] & b[18])^(a[167] & b[19])^(a[166] & b[20])^(a[165] & b[21])^(a[164] & b[22])^(a[163] & b[23])^(a[162] & b[24])^(a[161] & b[25])^(a[160] & b[26])^(a[159] & b[27])^(a[158] & b[28])^(a[157] & b[29])^(a[156] & b[30])^(a[155] & b[31])^(a[154] & b[32])^(a[153] & b[33])^(a[152] & b[34])^(a[151] & b[35])^(a[150] & b[36])^(a[149] & b[37])^(a[148] & b[38])^(a[147] & b[39])^(a[146] & b[40])^(a[145] & b[41])^(a[144] & b[42])^(a[143] & b[43])^(a[142] & b[44])^(a[141] & b[45])^(a[140] & b[46])^(a[139] & b[47])^(a[138] & b[48])^(a[137] & b[49])^(a[136] & b[50])^(a[135] & b[51])^(a[134] & b[52])^(a[133] & b[53])^(a[132] & b[54])^(a[131] & b[55])^(a[130] & b[56])^(a[129] & b[57])^(a[128] & b[58])^(a[127] & b[59])^(a[126] & b[60])^(a[125] & b[61])^(a[124] & b[62])^(a[123] & b[63])^(a[122] & b[64])^(a[121] & b[65])^(a[120] & b[66])^(a[119] & b[67])^(a[118] & b[68])^(a[117] & b[69])^(a[116] & b[70])^(a[115] & b[71])^(a[114] & b[72])^(a[113] & b[73])^(a[112] & b[74])^(a[111] & b[75])^(a[110] & b[76])^(a[109] & b[77])^(a[108] & b[78])^(a[107] & b[79])^(a[106] & b[80])^(a[105] & b[81])^(a[104] & b[82])^(a[103] & b[83])^(a[102] & b[84])^(a[101] & b[85])^(a[100] & b[86])^(a[99] & b[87])^(a[98] & b[88])^(a[97] & b[89])^(a[96] & b[90])^(a[95] & b[91])^(a[94] & b[92])^(a[93] & b[93])^(a[92] & b[94])^(a[91] & b[95])^(a[90] & b[96])^(a[89] & b[97])^(a[88] & b[98])^(a[87] & b[99])^(a[86] & b[100])^(a[85] & b[101])^(a[84] & b[102])^(a[83] & b[103])^(a[82] & b[104])^(a[81] & b[105])^(a[80] & b[106])^(a[79] & b[107])^(a[78] & b[108])^(a[77] & b[109])^(a[76] & b[110])^(a[75] & b[111])^(a[74] & b[112])^(a[73] & b[113])^(a[72] & b[114])^(a[71] & b[115])^(a[70] & b[116])^(a[69] & b[117])^(a[68] & b[118])^(a[67] & b[119])^(a[66] & b[120])^(a[65] & b[121])^(a[64] & b[122])^(a[63] & b[123])^(a[62] & b[124])^(a[61] & b[125])^(a[60] & b[126])^(a[59] & b[127])^(a[58] & b[128])^(a[57] & b[129])^(a[56] & b[130])^(a[55] & b[131])^(a[54] & b[132])^(a[53] & b[133])^(a[52] & b[134])^(a[51] & b[135])^(a[50] & b[136])^(a[49] & b[137])^(a[48] & b[138])^(a[47] & b[139])^(a[46] & b[140])^(a[45] & b[141])^(a[44] & b[142])^(a[43] & b[143])^(a[42] & b[144])^(a[41] & b[145])^(a[40] & b[146])^(a[39] & b[147])^(a[38] & b[148])^(a[37] & b[149])^(a[36] & b[150])^(a[35] & b[151])^(a[34] & b[152])^(a[33] & b[153])^(a[32] & b[154])^(a[31] & b[155])^(a[30] & b[156])^(a[29] & b[157])^(a[28] & b[158])^(a[27] & b[159])^(a[26] & b[160])^(a[25] & b[161])^(a[24] & b[162])^(a[23] & b[163])^(a[22] & b[164])^(a[21] & b[165])^(a[20] & b[166])^(a[19] & b[167])^(a[18] & b[168])^(a[17] & b[169])^(a[16] & b[170])^(a[15] & b[171])^(a[14] & b[172])^(a[13] & b[173])^(a[12] & b[174])^(a[11] & b[175])^(a[10] & b[176])^(a[9] & b[177])^(a[8] & b[178])^(a[7] & b[179])^(a[6] & b[180])^(a[5] & b[181])^(a[4] & b[182])^(a[3] & b[183])^(a[2] & b[184])^(a[1] & b[185])^(a[0] & b[186]);
assign y[187] = (a[187] & b[0])^(a[186] & b[1])^(a[185] & b[2])^(a[184] & b[3])^(a[183] & b[4])^(a[182] & b[5])^(a[181] & b[6])^(a[180] & b[7])^(a[179] & b[8])^(a[178] & b[9])^(a[177] & b[10])^(a[176] & b[11])^(a[175] & b[12])^(a[174] & b[13])^(a[173] & b[14])^(a[172] & b[15])^(a[171] & b[16])^(a[170] & b[17])^(a[169] & b[18])^(a[168] & b[19])^(a[167] & b[20])^(a[166] & b[21])^(a[165] & b[22])^(a[164] & b[23])^(a[163] & b[24])^(a[162] & b[25])^(a[161] & b[26])^(a[160] & b[27])^(a[159] & b[28])^(a[158] & b[29])^(a[157] & b[30])^(a[156] & b[31])^(a[155] & b[32])^(a[154] & b[33])^(a[153] & b[34])^(a[152] & b[35])^(a[151] & b[36])^(a[150] & b[37])^(a[149] & b[38])^(a[148] & b[39])^(a[147] & b[40])^(a[146] & b[41])^(a[145] & b[42])^(a[144] & b[43])^(a[143] & b[44])^(a[142] & b[45])^(a[141] & b[46])^(a[140] & b[47])^(a[139] & b[48])^(a[138] & b[49])^(a[137] & b[50])^(a[136] & b[51])^(a[135] & b[52])^(a[134] & b[53])^(a[133] & b[54])^(a[132] & b[55])^(a[131] & b[56])^(a[130] & b[57])^(a[129] & b[58])^(a[128] & b[59])^(a[127] & b[60])^(a[126] & b[61])^(a[125] & b[62])^(a[124] & b[63])^(a[123] & b[64])^(a[122] & b[65])^(a[121] & b[66])^(a[120] & b[67])^(a[119] & b[68])^(a[118] & b[69])^(a[117] & b[70])^(a[116] & b[71])^(a[115] & b[72])^(a[114] & b[73])^(a[113] & b[74])^(a[112] & b[75])^(a[111] & b[76])^(a[110] & b[77])^(a[109] & b[78])^(a[108] & b[79])^(a[107] & b[80])^(a[106] & b[81])^(a[105] & b[82])^(a[104] & b[83])^(a[103] & b[84])^(a[102] & b[85])^(a[101] & b[86])^(a[100] & b[87])^(a[99] & b[88])^(a[98] & b[89])^(a[97] & b[90])^(a[96] & b[91])^(a[95] & b[92])^(a[94] & b[93])^(a[93] & b[94])^(a[92] & b[95])^(a[91] & b[96])^(a[90] & b[97])^(a[89] & b[98])^(a[88] & b[99])^(a[87] & b[100])^(a[86] & b[101])^(a[85] & b[102])^(a[84] & b[103])^(a[83] & b[104])^(a[82] & b[105])^(a[81] & b[106])^(a[80] & b[107])^(a[79] & b[108])^(a[78] & b[109])^(a[77] & b[110])^(a[76] & b[111])^(a[75] & b[112])^(a[74] & b[113])^(a[73] & b[114])^(a[72] & b[115])^(a[71] & b[116])^(a[70] & b[117])^(a[69] & b[118])^(a[68] & b[119])^(a[67] & b[120])^(a[66] & b[121])^(a[65] & b[122])^(a[64] & b[123])^(a[63] & b[124])^(a[62] & b[125])^(a[61] & b[126])^(a[60] & b[127])^(a[59] & b[128])^(a[58] & b[129])^(a[57] & b[130])^(a[56] & b[131])^(a[55] & b[132])^(a[54] & b[133])^(a[53] & b[134])^(a[52] & b[135])^(a[51] & b[136])^(a[50] & b[137])^(a[49] & b[138])^(a[48] & b[139])^(a[47] & b[140])^(a[46] & b[141])^(a[45] & b[142])^(a[44] & b[143])^(a[43] & b[144])^(a[42] & b[145])^(a[41] & b[146])^(a[40] & b[147])^(a[39] & b[148])^(a[38] & b[149])^(a[37] & b[150])^(a[36] & b[151])^(a[35] & b[152])^(a[34] & b[153])^(a[33] & b[154])^(a[32] & b[155])^(a[31] & b[156])^(a[30] & b[157])^(a[29] & b[158])^(a[28] & b[159])^(a[27] & b[160])^(a[26] & b[161])^(a[25] & b[162])^(a[24] & b[163])^(a[23] & b[164])^(a[22] & b[165])^(a[21] & b[166])^(a[20] & b[167])^(a[19] & b[168])^(a[18] & b[169])^(a[17] & b[170])^(a[16] & b[171])^(a[15] & b[172])^(a[14] & b[173])^(a[13] & b[174])^(a[12] & b[175])^(a[11] & b[176])^(a[10] & b[177])^(a[9] & b[178])^(a[8] & b[179])^(a[7] & b[180])^(a[6] & b[181])^(a[5] & b[182])^(a[4] & b[183])^(a[3] & b[184])^(a[2] & b[185])^(a[1] & b[186])^(a[0] & b[187]);
assign y[188] = (a[188] & b[0])^(a[187] & b[1])^(a[186] & b[2])^(a[185] & b[3])^(a[184] & b[4])^(a[183] & b[5])^(a[182] & b[6])^(a[181] & b[7])^(a[180] & b[8])^(a[179] & b[9])^(a[178] & b[10])^(a[177] & b[11])^(a[176] & b[12])^(a[175] & b[13])^(a[174] & b[14])^(a[173] & b[15])^(a[172] & b[16])^(a[171] & b[17])^(a[170] & b[18])^(a[169] & b[19])^(a[168] & b[20])^(a[167] & b[21])^(a[166] & b[22])^(a[165] & b[23])^(a[164] & b[24])^(a[163] & b[25])^(a[162] & b[26])^(a[161] & b[27])^(a[160] & b[28])^(a[159] & b[29])^(a[158] & b[30])^(a[157] & b[31])^(a[156] & b[32])^(a[155] & b[33])^(a[154] & b[34])^(a[153] & b[35])^(a[152] & b[36])^(a[151] & b[37])^(a[150] & b[38])^(a[149] & b[39])^(a[148] & b[40])^(a[147] & b[41])^(a[146] & b[42])^(a[145] & b[43])^(a[144] & b[44])^(a[143] & b[45])^(a[142] & b[46])^(a[141] & b[47])^(a[140] & b[48])^(a[139] & b[49])^(a[138] & b[50])^(a[137] & b[51])^(a[136] & b[52])^(a[135] & b[53])^(a[134] & b[54])^(a[133] & b[55])^(a[132] & b[56])^(a[131] & b[57])^(a[130] & b[58])^(a[129] & b[59])^(a[128] & b[60])^(a[127] & b[61])^(a[126] & b[62])^(a[125] & b[63])^(a[124] & b[64])^(a[123] & b[65])^(a[122] & b[66])^(a[121] & b[67])^(a[120] & b[68])^(a[119] & b[69])^(a[118] & b[70])^(a[117] & b[71])^(a[116] & b[72])^(a[115] & b[73])^(a[114] & b[74])^(a[113] & b[75])^(a[112] & b[76])^(a[111] & b[77])^(a[110] & b[78])^(a[109] & b[79])^(a[108] & b[80])^(a[107] & b[81])^(a[106] & b[82])^(a[105] & b[83])^(a[104] & b[84])^(a[103] & b[85])^(a[102] & b[86])^(a[101] & b[87])^(a[100] & b[88])^(a[99] & b[89])^(a[98] & b[90])^(a[97] & b[91])^(a[96] & b[92])^(a[95] & b[93])^(a[94] & b[94])^(a[93] & b[95])^(a[92] & b[96])^(a[91] & b[97])^(a[90] & b[98])^(a[89] & b[99])^(a[88] & b[100])^(a[87] & b[101])^(a[86] & b[102])^(a[85] & b[103])^(a[84] & b[104])^(a[83] & b[105])^(a[82] & b[106])^(a[81] & b[107])^(a[80] & b[108])^(a[79] & b[109])^(a[78] & b[110])^(a[77] & b[111])^(a[76] & b[112])^(a[75] & b[113])^(a[74] & b[114])^(a[73] & b[115])^(a[72] & b[116])^(a[71] & b[117])^(a[70] & b[118])^(a[69] & b[119])^(a[68] & b[120])^(a[67] & b[121])^(a[66] & b[122])^(a[65] & b[123])^(a[64] & b[124])^(a[63] & b[125])^(a[62] & b[126])^(a[61] & b[127])^(a[60] & b[128])^(a[59] & b[129])^(a[58] & b[130])^(a[57] & b[131])^(a[56] & b[132])^(a[55] & b[133])^(a[54] & b[134])^(a[53] & b[135])^(a[52] & b[136])^(a[51] & b[137])^(a[50] & b[138])^(a[49] & b[139])^(a[48] & b[140])^(a[47] & b[141])^(a[46] & b[142])^(a[45] & b[143])^(a[44] & b[144])^(a[43] & b[145])^(a[42] & b[146])^(a[41] & b[147])^(a[40] & b[148])^(a[39] & b[149])^(a[38] & b[150])^(a[37] & b[151])^(a[36] & b[152])^(a[35] & b[153])^(a[34] & b[154])^(a[33] & b[155])^(a[32] & b[156])^(a[31] & b[157])^(a[30] & b[158])^(a[29] & b[159])^(a[28] & b[160])^(a[27] & b[161])^(a[26] & b[162])^(a[25] & b[163])^(a[24] & b[164])^(a[23] & b[165])^(a[22] & b[166])^(a[21] & b[167])^(a[20] & b[168])^(a[19] & b[169])^(a[18] & b[170])^(a[17] & b[171])^(a[16] & b[172])^(a[15] & b[173])^(a[14] & b[174])^(a[13] & b[175])^(a[12] & b[176])^(a[11] & b[177])^(a[10] & b[178])^(a[9] & b[179])^(a[8] & b[180])^(a[7] & b[181])^(a[6] & b[182])^(a[5] & b[183])^(a[4] & b[184])^(a[3] & b[185])^(a[2] & b[186])^(a[1] & b[187])^(a[0] & b[188]);
assign y[189] = (a[189] & b[0])^(a[188] & b[1])^(a[187] & b[2])^(a[186] & b[3])^(a[185] & b[4])^(a[184] & b[5])^(a[183] & b[6])^(a[182] & b[7])^(a[181] & b[8])^(a[180] & b[9])^(a[179] & b[10])^(a[178] & b[11])^(a[177] & b[12])^(a[176] & b[13])^(a[175] & b[14])^(a[174] & b[15])^(a[173] & b[16])^(a[172] & b[17])^(a[171] & b[18])^(a[170] & b[19])^(a[169] & b[20])^(a[168] & b[21])^(a[167] & b[22])^(a[166] & b[23])^(a[165] & b[24])^(a[164] & b[25])^(a[163] & b[26])^(a[162] & b[27])^(a[161] & b[28])^(a[160] & b[29])^(a[159] & b[30])^(a[158] & b[31])^(a[157] & b[32])^(a[156] & b[33])^(a[155] & b[34])^(a[154] & b[35])^(a[153] & b[36])^(a[152] & b[37])^(a[151] & b[38])^(a[150] & b[39])^(a[149] & b[40])^(a[148] & b[41])^(a[147] & b[42])^(a[146] & b[43])^(a[145] & b[44])^(a[144] & b[45])^(a[143] & b[46])^(a[142] & b[47])^(a[141] & b[48])^(a[140] & b[49])^(a[139] & b[50])^(a[138] & b[51])^(a[137] & b[52])^(a[136] & b[53])^(a[135] & b[54])^(a[134] & b[55])^(a[133] & b[56])^(a[132] & b[57])^(a[131] & b[58])^(a[130] & b[59])^(a[129] & b[60])^(a[128] & b[61])^(a[127] & b[62])^(a[126] & b[63])^(a[125] & b[64])^(a[124] & b[65])^(a[123] & b[66])^(a[122] & b[67])^(a[121] & b[68])^(a[120] & b[69])^(a[119] & b[70])^(a[118] & b[71])^(a[117] & b[72])^(a[116] & b[73])^(a[115] & b[74])^(a[114] & b[75])^(a[113] & b[76])^(a[112] & b[77])^(a[111] & b[78])^(a[110] & b[79])^(a[109] & b[80])^(a[108] & b[81])^(a[107] & b[82])^(a[106] & b[83])^(a[105] & b[84])^(a[104] & b[85])^(a[103] & b[86])^(a[102] & b[87])^(a[101] & b[88])^(a[100] & b[89])^(a[99] & b[90])^(a[98] & b[91])^(a[97] & b[92])^(a[96] & b[93])^(a[95] & b[94])^(a[94] & b[95])^(a[93] & b[96])^(a[92] & b[97])^(a[91] & b[98])^(a[90] & b[99])^(a[89] & b[100])^(a[88] & b[101])^(a[87] & b[102])^(a[86] & b[103])^(a[85] & b[104])^(a[84] & b[105])^(a[83] & b[106])^(a[82] & b[107])^(a[81] & b[108])^(a[80] & b[109])^(a[79] & b[110])^(a[78] & b[111])^(a[77] & b[112])^(a[76] & b[113])^(a[75] & b[114])^(a[74] & b[115])^(a[73] & b[116])^(a[72] & b[117])^(a[71] & b[118])^(a[70] & b[119])^(a[69] & b[120])^(a[68] & b[121])^(a[67] & b[122])^(a[66] & b[123])^(a[65] & b[124])^(a[64] & b[125])^(a[63] & b[126])^(a[62] & b[127])^(a[61] & b[128])^(a[60] & b[129])^(a[59] & b[130])^(a[58] & b[131])^(a[57] & b[132])^(a[56] & b[133])^(a[55] & b[134])^(a[54] & b[135])^(a[53] & b[136])^(a[52] & b[137])^(a[51] & b[138])^(a[50] & b[139])^(a[49] & b[140])^(a[48] & b[141])^(a[47] & b[142])^(a[46] & b[143])^(a[45] & b[144])^(a[44] & b[145])^(a[43] & b[146])^(a[42] & b[147])^(a[41] & b[148])^(a[40] & b[149])^(a[39] & b[150])^(a[38] & b[151])^(a[37] & b[152])^(a[36] & b[153])^(a[35] & b[154])^(a[34] & b[155])^(a[33] & b[156])^(a[32] & b[157])^(a[31] & b[158])^(a[30] & b[159])^(a[29] & b[160])^(a[28] & b[161])^(a[27] & b[162])^(a[26] & b[163])^(a[25] & b[164])^(a[24] & b[165])^(a[23] & b[166])^(a[22] & b[167])^(a[21] & b[168])^(a[20] & b[169])^(a[19] & b[170])^(a[18] & b[171])^(a[17] & b[172])^(a[16] & b[173])^(a[15] & b[174])^(a[14] & b[175])^(a[13] & b[176])^(a[12] & b[177])^(a[11] & b[178])^(a[10] & b[179])^(a[9] & b[180])^(a[8] & b[181])^(a[7] & b[182])^(a[6] & b[183])^(a[5] & b[184])^(a[4] & b[185])^(a[3] & b[186])^(a[2] & b[187])^(a[1] & b[188])^(a[0] & b[189]);
assign y[190] = (a[190] & b[0])^(a[189] & b[1])^(a[188] & b[2])^(a[187] & b[3])^(a[186] & b[4])^(a[185] & b[5])^(a[184] & b[6])^(a[183] & b[7])^(a[182] & b[8])^(a[181] & b[9])^(a[180] & b[10])^(a[179] & b[11])^(a[178] & b[12])^(a[177] & b[13])^(a[176] & b[14])^(a[175] & b[15])^(a[174] & b[16])^(a[173] & b[17])^(a[172] & b[18])^(a[171] & b[19])^(a[170] & b[20])^(a[169] & b[21])^(a[168] & b[22])^(a[167] & b[23])^(a[166] & b[24])^(a[165] & b[25])^(a[164] & b[26])^(a[163] & b[27])^(a[162] & b[28])^(a[161] & b[29])^(a[160] & b[30])^(a[159] & b[31])^(a[158] & b[32])^(a[157] & b[33])^(a[156] & b[34])^(a[155] & b[35])^(a[154] & b[36])^(a[153] & b[37])^(a[152] & b[38])^(a[151] & b[39])^(a[150] & b[40])^(a[149] & b[41])^(a[148] & b[42])^(a[147] & b[43])^(a[146] & b[44])^(a[145] & b[45])^(a[144] & b[46])^(a[143] & b[47])^(a[142] & b[48])^(a[141] & b[49])^(a[140] & b[50])^(a[139] & b[51])^(a[138] & b[52])^(a[137] & b[53])^(a[136] & b[54])^(a[135] & b[55])^(a[134] & b[56])^(a[133] & b[57])^(a[132] & b[58])^(a[131] & b[59])^(a[130] & b[60])^(a[129] & b[61])^(a[128] & b[62])^(a[127] & b[63])^(a[126] & b[64])^(a[125] & b[65])^(a[124] & b[66])^(a[123] & b[67])^(a[122] & b[68])^(a[121] & b[69])^(a[120] & b[70])^(a[119] & b[71])^(a[118] & b[72])^(a[117] & b[73])^(a[116] & b[74])^(a[115] & b[75])^(a[114] & b[76])^(a[113] & b[77])^(a[112] & b[78])^(a[111] & b[79])^(a[110] & b[80])^(a[109] & b[81])^(a[108] & b[82])^(a[107] & b[83])^(a[106] & b[84])^(a[105] & b[85])^(a[104] & b[86])^(a[103] & b[87])^(a[102] & b[88])^(a[101] & b[89])^(a[100] & b[90])^(a[99] & b[91])^(a[98] & b[92])^(a[97] & b[93])^(a[96] & b[94])^(a[95] & b[95])^(a[94] & b[96])^(a[93] & b[97])^(a[92] & b[98])^(a[91] & b[99])^(a[90] & b[100])^(a[89] & b[101])^(a[88] & b[102])^(a[87] & b[103])^(a[86] & b[104])^(a[85] & b[105])^(a[84] & b[106])^(a[83] & b[107])^(a[82] & b[108])^(a[81] & b[109])^(a[80] & b[110])^(a[79] & b[111])^(a[78] & b[112])^(a[77] & b[113])^(a[76] & b[114])^(a[75] & b[115])^(a[74] & b[116])^(a[73] & b[117])^(a[72] & b[118])^(a[71] & b[119])^(a[70] & b[120])^(a[69] & b[121])^(a[68] & b[122])^(a[67] & b[123])^(a[66] & b[124])^(a[65] & b[125])^(a[64] & b[126])^(a[63] & b[127])^(a[62] & b[128])^(a[61] & b[129])^(a[60] & b[130])^(a[59] & b[131])^(a[58] & b[132])^(a[57] & b[133])^(a[56] & b[134])^(a[55] & b[135])^(a[54] & b[136])^(a[53] & b[137])^(a[52] & b[138])^(a[51] & b[139])^(a[50] & b[140])^(a[49] & b[141])^(a[48] & b[142])^(a[47] & b[143])^(a[46] & b[144])^(a[45] & b[145])^(a[44] & b[146])^(a[43] & b[147])^(a[42] & b[148])^(a[41] & b[149])^(a[40] & b[150])^(a[39] & b[151])^(a[38] & b[152])^(a[37] & b[153])^(a[36] & b[154])^(a[35] & b[155])^(a[34] & b[156])^(a[33] & b[157])^(a[32] & b[158])^(a[31] & b[159])^(a[30] & b[160])^(a[29] & b[161])^(a[28] & b[162])^(a[27] & b[163])^(a[26] & b[164])^(a[25] & b[165])^(a[24] & b[166])^(a[23] & b[167])^(a[22] & b[168])^(a[21] & b[169])^(a[20] & b[170])^(a[19] & b[171])^(a[18] & b[172])^(a[17] & b[173])^(a[16] & b[174])^(a[15] & b[175])^(a[14] & b[176])^(a[13] & b[177])^(a[12] & b[178])^(a[11] & b[179])^(a[10] & b[180])^(a[9] & b[181])^(a[8] & b[182])^(a[7] & b[183])^(a[6] & b[184])^(a[5] & b[185])^(a[4] & b[186])^(a[3] & b[187])^(a[2] & b[188])^(a[1] & b[189])^(a[0] & b[190]);
assign y[191] = (a[191] & b[0])^(a[190] & b[1])^(a[189] & b[2])^(a[188] & b[3])^(a[187] & b[4])^(a[186] & b[5])^(a[185] & b[6])^(a[184] & b[7])^(a[183] & b[8])^(a[182] & b[9])^(a[181] & b[10])^(a[180] & b[11])^(a[179] & b[12])^(a[178] & b[13])^(a[177] & b[14])^(a[176] & b[15])^(a[175] & b[16])^(a[174] & b[17])^(a[173] & b[18])^(a[172] & b[19])^(a[171] & b[20])^(a[170] & b[21])^(a[169] & b[22])^(a[168] & b[23])^(a[167] & b[24])^(a[166] & b[25])^(a[165] & b[26])^(a[164] & b[27])^(a[163] & b[28])^(a[162] & b[29])^(a[161] & b[30])^(a[160] & b[31])^(a[159] & b[32])^(a[158] & b[33])^(a[157] & b[34])^(a[156] & b[35])^(a[155] & b[36])^(a[154] & b[37])^(a[153] & b[38])^(a[152] & b[39])^(a[151] & b[40])^(a[150] & b[41])^(a[149] & b[42])^(a[148] & b[43])^(a[147] & b[44])^(a[146] & b[45])^(a[145] & b[46])^(a[144] & b[47])^(a[143] & b[48])^(a[142] & b[49])^(a[141] & b[50])^(a[140] & b[51])^(a[139] & b[52])^(a[138] & b[53])^(a[137] & b[54])^(a[136] & b[55])^(a[135] & b[56])^(a[134] & b[57])^(a[133] & b[58])^(a[132] & b[59])^(a[131] & b[60])^(a[130] & b[61])^(a[129] & b[62])^(a[128] & b[63])^(a[127] & b[64])^(a[126] & b[65])^(a[125] & b[66])^(a[124] & b[67])^(a[123] & b[68])^(a[122] & b[69])^(a[121] & b[70])^(a[120] & b[71])^(a[119] & b[72])^(a[118] & b[73])^(a[117] & b[74])^(a[116] & b[75])^(a[115] & b[76])^(a[114] & b[77])^(a[113] & b[78])^(a[112] & b[79])^(a[111] & b[80])^(a[110] & b[81])^(a[109] & b[82])^(a[108] & b[83])^(a[107] & b[84])^(a[106] & b[85])^(a[105] & b[86])^(a[104] & b[87])^(a[103] & b[88])^(a[102] & b[89])^(a[101] & b[90])^(a[100] & b[91])^(a[99] & b[92])^(a[98] & b[93])^(a[97] & b[94])^(a[96] & b[95])^(a[95] & b[96])^(a[94] & b[97])^(a[93] & b[98])^(a[92] & b[99])^(a[91] & b[100])^(a[90] & b[101])^(a[89] & b[102])^(a[88] & b[103])^(a[87] & b[104])^(a[86] & b[105])^(a[85] & b[106])^(a[84] & b[107])^(a[83] & b[108])^(a[82] & b[109])^(a[81] & b[110])^(a[80] & b[111])^(a[79] & b[112])^(a[78] & b[113])^(a[77] & b[114])^(a[76] & b[115])^(a[75] & b[116])^(a[74] & b[117])^(a[73] & b[118])^(a[72] & b[119])^(a[71] & b[120])^(a[70] & b[121])^(a[69] & b[122])^(a[68] & b[123])^(a[67] & b[124])^(a[66] & b[125])^(a[65] & b[126])^(a[64] & b[127])^(a[63] & b[128])^(a[62] & b[129])^(a[61] & b[130])^(a[60] & b[131])^(a[59] & b[132])^(a[58] & b[133])^(a[57] & b[134])^(a[56] & b[135])^(a[55] & b[136])^(a[54] & b[137])^(a[53] & b[138])^(a[52] & b[139])^(a[51] & b[140])^(a[50] & b[141])^(a[49] & b[142])^(a[48] & b[143])^(a[47] & b[144])^(a[46] & b[145])^(a[45] & b[146])^(a[44] & b[147])^(a[43] & b[148])^(a[42] & b[149])^(a[41] & b[150])^(a[40] & b[151])^(a[39] & b[152])^(a[38] & b[153])^(a[37] & b[154])^(a[36] & b[155])^(a[35] & b[156])^(a[34] & b[157])^(a[33] & b[158])^(a[32] & b[159])^(a[31] & b[160])^(a[30] & b[161])^(a[29] & b[162])^(a[28] & b[163])^(a[27] & b[164])^(a[26] & b[165])^(a[25] & b[166])^(a[24] & b[167])^(a[23] & b[168])^(a[22] & b[169])^(a[21] & b[170])^(a[20] & b[171])^(a[19] & b[172])^(a[18] & b[173])^(a[17] & b[174])^(a[16] & b[175])^(a[15] & b[176])^(a[14] & b[177])^(a[13] & b[178])^(a[12] & b[179])^(a[11] & b[180])^(a[10] & b[181])^(a[9] & b[182])^(a[8] & b[183])^(a[7] & b[184])^(a[6] & b[185])^(a[5] & b[186])^(a[4] & b[187])^(a[3] & b[188])^(a[2] & b[189])^(a[1] & b[190])^(a[0] & b[191]);
assign y[192] = (a[192] & b[0])^(a[191] & b[1])^(a[190] & b[2])^(a[189] & b[3])^(a[188] & b[4])^(a[187] & b[5])^(a[186] & b[6])^(a[185] & b[7])^(a[184] & b[8])^(a[183] & b[9])^(a[182] & b[10])^(a[181] & b[11])^(a[180] & b[12])^(a[179] & b[13])^(a[178] & b[14])^(a[177] & b[15])^(a[176] & b[16])^(a[175] & b[17])^(a[174] & b[18])^(a[173] & b[19])^(a[172] & b[20])^(a[171] & b[21])^(a[170] & b[22])^(a[169] & b[23])^(a[168] & b[24])^(a[167] & b[25])^(a[166] & b[26])^(a[165] & b[27])^(a[164] & b[28])^(a[163] & b[29])^(a[162] & b[30])^(a[161] & b[31])^(a[160] & b[32])^(a[159] & b[33])^(a[158] & b[34])^(a[157] & b[35])^(a[156] & b[36])^(a[155] & b[37])^(a[154] & b[38])^(a[153] & b[39])^(a[152] & b[40])^(a[151] & b[41])^(a[150] & b[42])^(a[149] & b[43])^(a[148] & b[44])^(a[147] & b[45])^(a[146] & b[46])^(a[145] & b[47])^(a[144] & b[48])^(a[143] & b[49])^(a[142] & b[50])^(a[141] & b[51])^(a[140] & b[52])^(a[139] & b[53])^(a[138] & b[54])^(a[137] & b[55])^(a[136] & b[56])^(a[135] & b[57])^(a[134] & b[58])^(a[133] & b[59])^(a[132] & b[60])^(a[131] & b[61])^(a[130] & b[62])^(a[129] & b[63])^(a[128] & b[64])^(a[127] & b[65])^(a[126] & b[66])^(a[125] & b[67])^(a[124] & b[68])^(a[123] & b[69])^(a[122] & b[70])^(a[121] & b[71])^(a[120] & b[72])^(a[119] & b[73])^(a[118] & b[74])^(a[117] & b[75])^(a[116] & b[76])^(a[115] & b[77])^(a[114] & b[78])^(a[113] & b[79])^(a[112] & b[80])^(a[111] & b[81])^(a[110] & b[82])^(a[109] & b[83])^(a[108] & b[84])^(a[107] & b[85])^(a[106] & b[86])^(a[105] & b[87])^(a[104] & b[88])^(a[103] & b[89])^(a[102] & b[90])^(a[101] & b[91])^(a[100] & b[92])^(a[99] & b[93])^(a[98] & b[94])^(a[97] & b[95])^(a[96] & b[96])^(a[95] & b[97])^(a[94] & b[98])^(a[93] & b[99])^(a[92] & b[100])^(a[91] & b[101])^(a[90] & b[102])^(a[89] & b[103])^(a[88] & b[104])^(a[87] & b[105])^(a[86] & b[106])^(a[85] & b[107])^(a[84] & b[108])^(a[83] & b[109])^(a[82] & b[110])^(a[81] & b[111])^(a[80] & b[112])^(a[79] & b[113])^(a[78] & b[114])^(a[77] & b[115])^(a[76] & b[116])^(a[75] & b[117])^(a[74] & b[118])^(a[73] & b[119])^(a[72] & b[120])^(a[71] & b[121])^(a[70] & b[122])^(a[69] & b[123])^(a[68] & b[124])^(a[67] & b[125])^(a[66] & b[126])^(a[65] & b[127])^(a[64] & b[128])^(a[63] & b[129])^(a[62] & b[130])^(a[61] & b[131])^(a[60] & b[132])^(a[59] & b[133])^(a[58] & b[134])^(a[57] & b[135])^(a[56] & b[136])^(a[55] & b[137])^(a[54] & b[138])^(a[53] & b[139])^(a[52] & b[140])^(a[51] & b[141])^(a[50] & b[142])^(a[49] & b[143])^(a[48] & b[144])^(a[47] & b[145])^(a[46] & b[146])^(a[45] & b[147])^(a[44] & b[148])^(a[43] & b[149])^(a[42] & b[150])^(a[41] & b[151])^(a[40] & b[152])^(a[39] & b[153])^(a[38] & b[154])^(a[37] & b[155])^(a[36] & b[156])^(a[35] & b[157])^(a[34] & b[158])^(a[33] & b[159])^(a[32] & b[160])^(a[31] & b[161])^(a[30] & b[162])^(a[29] & b[163])^(a[28] & b[164])^(a[27] & b[165])^(a[26] & b[166])^(a[25] & b[167])^(a[24] & b[168])^(a[23] & b[169])^(a[22] & b[170])^(a[21] & b[171])^(a[20] & b[172])^(a[19] & b[173])^(a[18] & b[174])^(a[17] & b[175])^(a[16] & b[176])^(a[15] & b[177])^(a[14] & b[178])^(a[13] & b[179])^(a[12] & b[180])^(a[11] & b[181])^(a[10] & b[182])^(a[9] & b[183])^(a[8] & b[184])^(a[7] & b[185])^(a[6] & b[186])^(a[5] & b[187])^(a[4] & b[188])^(a[3] & b[189])^(a[2] & b[190])^(a[1] & b[191])^(a[0] & b[192]);
assign y[193] = (a[193] & b[0])^(a[192] & b[1])^(a[191] & b[2])^(a[190] & b[3])^(a[189] & b[4])^(a[188] & b[5])^(a[187] & b[6])^(a[186] & b[7])^(a[185] & b[8])^(a[184] & b[9])^(a[183] & b[10])^(a[182] & b[11])^(a[181] & b[12])^(a[180] & b[13])^(a[179] & b[14])^(a[178] & b[15])^(a[177] & b[16])^(a[176] & b[17])^(a[175] & b[18])^(a[174] & b[19])^(a[173] & b[20])^(a[172] & b[21])^(a[171] & b[22])^(a[170] & b[23])^(a[169] & b[24])^(a[168] & b[25])^(a[167] & b[26])^(a[166] & b[27])^(a[165] & b[28])^(a[164] & b[29])^(a[163] & b[30])^(a[162] & b[31])^(a[161] & b[32])^(a[160] & b[33])^(a[159] & b[34])^(a[158] & b[35])^(a[157] & b[36])^(a[156] & b[37])^(a[155] & b[38])^(a[154] & b[39])^(a[153] & b[40])^(a[152] & b[41])^(a[151] & b[42])^(a[150] & b[43])^(a[149] & b[44])^(a[148] & b[45])^(a[147] & b[46])^(a[146] & b[47])^(a[145] & b[48])^(a[144] & b[49])^(a[143] & b[50])^(a[142] & b[51])^(a[141] & b[52])^(a[140] & b[53])^(a[139] & b[54])^(a[138] & b[55])^(a[137] & b[56])^(a[136] & b[57])^(a[135] & b[58])^(a[134] & b[59])^(a[133] & b[60])^(a[132] & b[61])^(a[131] & b[62])^(a[130] & b[63])^(a[129] & b[64])^(a[128] & b[65])^(a[127] & b[66])^(a[126] & b[67])^(a[125] & b[68])^(a[124] & b[69])^(a[123] & b[70])^(a[122] & b[71])^(a[121] & b[72])^(a[120] & b[73])^(a[119] & b[74])^(a[118] & b[75])^(a[117] & b[76])^(a[116] & b[77])^(a[115] & b[78])^(a[114] & b[79])^(a[113] & b[80])^(a[112] & b[81])^(a[111] & b[82])^(a[110] & b[83])^(a[109] & b[84])^(a[108] & b[85])^(a[107] & b[86])^(a[106] & b[87])^(a[105] & b[88])^(a[104] & b[89])^(a[103] & b[90])^(a[102] & b[91])^(a[101] & b[92])^(a[100] & b[93])^(a[99] & b[94])^(a[98] & b[95])^(a[97] & b[96])^(a[96] & b[97])^(a[95] & b[98])^(a[94] & b[99])^(a[93] & b[100])^(a[92] & b[101])^(a[91] & b[102])^(a[90] & b[103])^(a[89] & b[104])^(a[88] & b[105])^(a[87] & b[106])^(a[86] & b[107])^(a[85] & b[108])^(a[84] & b[109])^(a[83] & b[110])^(a[82] & b[111])^(a[81] & b[112])^(a[80] & b[113])^(a[79] & b[114])^(a[78] & b[115])^(a[77] & b[116])^(a[76] & b[117])^(a[75] & b[118])^(a[74] & b[119])^(a[73] & b[120])^(a[72] & b[121])^(a[71] & b[122])^(a[70] & b[123])^(a[69] & b[124])^(a[68] & b[125])^(a[67] & b[126])^(a[66] & b[127])^(a[65] & b[128])^(a[64] & b[129])^(a[63] & b[130])^(a[62] & b[131])^(a[61] & b[132])^(a[60] & b[133])^(a[59] & b[134])^(a[58] & b[135])^(a[57] & b[136])^(a[56] & b[137])^(a[55] & b[138])^(a[54] & b[139])^(a[53] & b[140])^(a[52] & b[141])^(a[51] & b[142])^(a[50] & b[143])^(a[49] & b[144])^(a[48] & b[145])^(a[47] & b[146])^(a[46] & b[147])^(a[45] & b[148])^(a[44] & b[149])^(a[43] & b[150])^(a[42] & b[151])^(a[41] & b[152])^(a[40] & b[153])^(a[39] & b[154])^(a[38] & b[155])^(a[37] & b[156])^(a[36] & b[157])^(a[35] & b[158])^(a[34] & b[159])^(a[33] & b[160])^(a[32] & b[161])^(a[31] & b[162])^(a[30] & b[163])^(a[29] & b[164])^(a[28] & b[165])^(a[27] & b[166])^(a[26] & b[167])^(a[25] & b[168])^(a[24] & b[169])^(a[23] & b[170])^(a[22] & b[171])^(a[21] & b[172])^(a[20] & b[173])^(a[19] & b[174])^(a[18] & b[175])^(a[17] & b[176])^(a[16] & b[177])^(a[15] & b[178])^(a[14] & b[179])^(a[13] & b[180])^(a[12] & b[181])^(a[11] & b[182])^(a[10] & b[183])^(a[9] & b[184])^(a[8] & b[185])^(a[7] & b[186])^(a[6] & b[187])^(a[5] & b[188])^(a[4] & b[189])^(a[3] & b[190])^(a[2] & b[191])^(a[1] & b[192])^(a[0] & b[193]);
assign y[194] = (a[194] & b[0])^(a[193] & b[1])^(a[192] & b[2])^(a[191] & b[3])^(a[190] & b[4])^(a[189] & b[5])^(a[188] & b[6])^(a[187] & b[7])^(a[186] & b[8])^(a[185] & b[9])^(a[184] & b[10])^(a[183] & b[11])^(a[182] & b[12])^(a[181] & b[13])^(a[180] & b[14])^(a[179] & b[15])^(a[178] & b[16])^(a[177] & b[17])^(a[176] & b[18])^(a[175] & b[19])^(a[174] & b[20])^(a[173] & b[21])^(a[172] & b[22])^(a[171] & b[23])^(a[170] & b[24])^(a[169] & b[25])^(a[168] & b[26])^(a[167] & b[27])^(a[166] & b[28])^(a[165] & b[29])^(a[164] & b[30])^(a[163] & b[31])^(a[162] & b[32])^(a[161] & b[33])^(a[160] & b[34])^(a[159] & b[35])^(a[158] & b[36])^(a[157] & b[37])^(a[156] & b[38])^(a[155] & b[39])^(a[154] & b[40])^(a[153] & b[41])^(a[152] & b[42])^(a[151] & b[43])^(a[150] & b[44])^(a[149] & b[45])^(a[148] & b[46])^(a[147] & b[47])^(a[146] & b[48])^(a[145] & b[49])^(a[144] & b[50])^(a[143] & b[51])^(a[142] & b[52])^(a[141] & b[53])^(a[140] & b[54])^(a[139] & b[55])^(a[138] & b[56])^(a[137] & b[57])^(a[136] & b[58])^(a[135] & b[59])^(a[134] & b[60])^(a[133] & b[61])^(a[132] & b[62])^(a[131] & b[63])^(a[130] & b[64])^(a[129] & b[65])^(a[128] & b[66])^(a[127] & b[67])^(a[126] & b[68])^(a[125] & b[69])^(a[124] & b[70])^(a[123] & b[71])^(a[122] & b[72])^(a[121] & b[73])^(a[120] & b[74])^(a[119] & b[75])^(a[118] & b[76])^(a[117] & b[77])^(a[116] & b[78])^(a[115] & b[79])^(a[114] & b[80])^(a[113] & b[81])^(a[112] & b[82])^(a[111] & b[83])^(a[110] & b[84])^(a[109] & b[85])^(a[108] & b[86])^(a[107] & b[87])^(a[106] & b[88])^(a[105] & b[89])^(a[104] & b[90])^(a[103] & b[91])^(a[102] & b[92])^(a[101] & b[93])^(a[100] & b[94])^(a[99] & b[95])^(a[98] & b[96])^(a[97] & b[97])^(a[96] & b[98])^(a[95] & b[99])^(a[94] & b[100])^(a[93] & b[101])^(a[92] & b[102])^(a[91] & b[103])^(a[90] & b[104])^(a[89] & b[105])^(a[88] & b[106])^(a[87] & b[107])^(a[86] & b[108])^(a[85] & b[109])^(a[84] & b[110])^(a[83] & b[111])^(a[82] & b[112])^(a[81] & b[113])^(a[80] & b[114])^(a[79] & b[115])^(a[78] & b[116])^(a[77] & b[117])^(a[76] & b[118])^(a[75] & b[119])^(a[74] & b[120])^(a[73] & b[121])^(a[72] & b[122])^(a[71] & b[123])^(a[70] & b[124])^(a[69] & b[125])^(a[68] & b[126])^(a[67] & b[127])^(a[66] & b[128])^(a[65] & b[129])^(a[64] & b[130])^(a[63] & b[131])^(a[62] & b[132])^(a[61] & b[133])^(a[60] & b[134])^(a[59] & b[135])^(a[58] & b[136])^(a[57] & b[137])^(a[56] & b[138])^(a[55] & b[139])^(a[54] & b[140])^(a[53] & b[141])^(a[52] & b[142])^(a[51] & b[143])^(a[50] & b[144])^(a[49] & b[145])^(a[48] & b[146])^(a[47] & b[147])^(a[46] & b[148])^(a[45] & b[149])^(a[44] & b[150])^(a[43] & b[151])^(a[42] & b[152])^(a[41] & b[153])^(a[40] & b[154])^(a[39] & b[155])^(a[38] & b[156])^(a[37] & b[157])^(a[36] & b[158])^(a[35] & b[159])^(a[34] & b[160])^(a[33] & b[161])^(a[32] & b[162])^(a[31] & b[163])^(a[30] & b[164])^(a[29] & b[165])^(a[28] & b[166])^(a[27] & b[167])^(a[26] & b[168])^(a[25] & b[169])^(a[24] & b[170])^(a[23] & b[171])^(a[22] & b[172])^(a[21] & b[173])^(a[20] & b[174])^(a[19] & b[175])^(a[18] & b[176])^(a[17] & b[177])^(a[16] & b[178])^(a[15] & b[179])^(a[14] & b[180])^(a[13] & b[181])^(a[12] & b[182])^(a[11] & b[183])^(a[10] & b[184])^(a[9] & b[185])^(a[8] & b[186])^(a[7] & b[187])^(a[6] & b[188])^(a[5] & b[189])^(a[4] & b[190])^(a[3] & b[191])^(a[2] & b[192])^(a[1] & b[193])^(a[0] & b[194]);
assign y[195] = (a[195] & b[0])^(a[194] & b[1])^(a[193] & b[2])^(a[192] & b[3])^(a[191] & b[4])^(a[190] & b[5])^(a[189] & b[6])^(a[188] & b[7])^(a[187] & b[8])^(a[186] & b[9])^(a[185] & b[10])^(a[184] & b[11])^(a[183] & b[12])^(a[182] & b[13])^(a[181] & b[14])^(a[180] & b[15])^(a[179] & b[16])^(a[178] & b[17])^(a[177] & b[18])^(a[176] & b[19])^(a[175] & b[20])^(a[174] & b[21])^(a[173] & b[22])^(a[172] & b[23])^(a[171] & b[24])^(a[170] & b[25])^(a[169] & b[26])^(a[168] & b[27])^(a[167] & b[28])^(a[166] & b[29])^(a[165] & b[30])^(a[164] & b[31])^(a[163] & b[32])^(a[162] & b[33])^(a[161] & b[34])^(a[160] & b[35])^(a[159] & b[36])^(a[158] & b[37])^(a[157] & b[38])^(a[156] & b[39])^(a[155] & b[40])^(a[154] & b[41])^(a[153] & b[42])^(a[152] & b[43])^(a[151] & b[44])^(a[150] & b[45])^(a[149] & b[46])^(a[148] & b[47])^(a[147] & b[48])^(a[146] & b[49])^(a[145] & b[50])^(a[144] & b[51])^(a[143] & b[52])^(a[142] & b[53])^(a[141] & b[54])^(a[140] & b[55])^(a[139] & b[56])^(a[138] & b[57])^(a[137] & b[58])^(a[136] & b[59])^(a[135] & b[60])^(a[134] & b[61])^(a[133] & b[62])^(a[132] & b[63])^(a[131] & b[64])^(a[130] & b[65])^(a[129] & b[66])^(a[128] & b[67])^(a[127] & b[68])^(a[126] & b[69])^(a[125] & b[70])^(a[124] & b[71])^(a[123] & b[72])^(a[122] & b[73])^(a[121] & b[74])^(a[120] & b[75])^(a[119] & b[76])^(a[118] & b[77])^(a[117] & b[78])^(a[116] & b[79])^(a[115] & b[80])^(a[114] & b[81])^(a[113] & b[82])^(a[112] & b[83])^(a[111] & b[84])^(a[110] & b[85])^(a[109] & b[86])^(a[108] & b[87])^(a[107] & b[88])^(a[106] & b[89])^(a[105] & b[90])^(a[104] & b[91])^(a[103] & b[92])^(a[102] & b[93])^(a[101] & b[94])^(a[100] & b[95])^(a[99] & b[96])^(a[98] & b[97])^(a[97] & b[98])^(a[96] & b[99])^(a[95] & b[100])^(a[94] & b[101])^(a[93] & b[102])^(a[92] & b[103])^(a[91] & b[104])^(a[90] & b[105])^(a[89] & b[106])^(a[88] & b[107])^(a[87] & b[108])^(a[86] & b[109])^(a[85] & b[110])^(a[84] & b[111])^(a[83] & b[112])^(a[82] & b[113])^(a[81] & b[114])^(a[80] & b[115])^(a[79] & b[116])^(a[78] & b[117])^(a[77] & b[118])^(a[76] & b[119])^(a[75] & b[120])^(a[74] & b[121])^(a[73] & b[122])^(a[72] & b[123])^(a[71] & b[124])^(a[70] & b[125])^(a[69] & b[126])^(a[68] & b[127])^(a[67] & b[128])^(a[66] & b[129])^(a[65] & b[130])^(a[64] & b[131])^(a[63] & b[132])^(a[62] & b[133])^(a[61] & b[134])^(a[60] & b[135])^(a[59] & b[136])^(a[58] & b[137])^(a[57] & b[138])^(a[56] & b[139])^(a[55] & b[140])^(a[54] & b[141])^(a[53] & b[142])^(a[52] & b[143])^(a[51] & b[144])^(a[50] & b[145])^(a[49] & b[146])^(a[48] & b[147])^(a[47] & b[148])^(a[46] & b[149])^(a[45] & b[150])^(a[44] & b[151])^(a[43] & b[152])^(a[42] & b[153])^(a[41] & b[154])^(a[40] & b[155])^(a[39] & b[156])^(a[38] & b[157])^(a[37] & b[158])^(a[36] & b[159])^(a[35] & b[160])^(a[34] & b[161])^(a[33] & b[162])^(a[32] & b[163])^(a[31] & b[164])^(a[30] & b[165])^(a[29] & b[166])^(a[28] & b[167])^(a[27] & b[168])^(a[26] & b[169])^(a[25] & b[170])^(a[24] & b[171])^(a[23] & b[172])^(a[22] & b[173])^(a[21] & b[174])^(a[20] & b[175])^(a[19] & b[176])^(a[18] & b[177])^(a[17] & b[178])^(a[16] & b[179])^(a[15] & b[180])^(a[14] & b[181])^(a[13] & b[182])^(a[12] & b[183])^(a[11] & b[184])^(a[10] & b[185])^(a[9] & b[186])^(a[8] & b[187])^(a[7] & b[188])^(a[6] & b[189])^(a[5] & b[190])^(a[4] & b[191])^(a[3] & b[192])^(a[2] & b[193])^(a[1] & b[194])^(a[0] & b[195]);
assign y[196] = (a[196] & b[0])^(a[195] & b[1])^(a[194] & b[2])^(a[193] & b[3])^(a[192] & b[4])^(a[191] & b[5])^(a[190] & b[6])^(a[189] & b[7])^(a[188] & b[8])^(a[187] & b[9])^(a[186] & b[10])^(a[185] & b[11])^(a[184] & b[12])^(a[183] & b[13])^(a[182] & b[14])^(a[181] & b[15])^(a[180] & b[16])^(a[179] & b[17])^(a[178] & b[18])^(a[177] & b[19])^(a[176] & b[20])^(a[175] & b[21])^(a[174] & b[22])^(a[173] & b[23])^(a[172] & b[24])^(a[171] & b[25])^(a[170] & b[26])^(a[169] & b[27])^(a[168] & b[28])^(a[167] & b[29])^(a[166] & b[30])^(a[165] & b[31])^(a[164] & b[32])^(a[163] & b[33])^(a[162] & b[34])^(a[161] & b[35])^(a[160] & b[36])^(a[159] & b[37])^(a[158] & b[38])^(a[157] & b[39])^(a[156] & b[40])^(a[155] & b[41])^(a[154] & b[42])^(a[153] & b[43])^(a[152] & b[44])^(a[151] & b[45])^(a[150] & b[46])^(a[149] & b[47])^(a[148] & b[48])^(a[147] & b[49])^(a[146] & b[50])^(a[145] & b[51])^(a[144] & b[52])^(a[143] & b[53])^(a[142] & b[54])^(a[141] & b[55])^(a[140] & b[56])^(a[139] & b[57])^(a[138] & b[58])^(a[137] & b[59])^(a[136] & b[60])^(a[135] & b[61])^(a[134] & b[62])^(a[133] & b[63])^(a[132] & b[64])^(a[131] & b[65])^(a[130] & b[66])^(a[129] & b[67])^(a[128] & b[68])^(a[127] & b[69])^(a[126] & b[70])^(a[125] & b[71])^(a[124] & b[72])^(a[123] & b[73])^(a[122] & b[74])^(a[121] & b[75])^(a[120] & b[76])^(a[119] & b[77])^(a[118] & b[78])^(a[117] & b[79])^(a[116] & b[80])^(a[115] & b[81])^(a[114] & b[82])^(a[113] & b[83])^(a[112] & b[84])^(a[111] & b[85])^(a[110] & b[86])^(a[109] & b[87])^(a[108] & b[88])^(a[107] & b[89])^(a[106] & b[90])^(a[105] & b[91])^(a[104] & b[92])^(a[103] & b[93])^(a[102] & b[94])^(a[101] & b[95])^(a[100] & b[96])^(a[99] & b[97])^(a[98] & b[98])^(a[97] & b[99])^(a[96] & b[100])^(a[95] & b[101])^(a[94] & b[102])^(a[93] & b[103])^(a[92] & b[104])^(a[91] & b[105])^(a[90] & b[106])^(a[89] & b[107])^(a[88] & b[108])^(a[87] & b[109])^(a[86] & b[110])^(a[85] & b[111])^(a[84] & b[112])^(a[83] & b[113])^(a[82] & b[114])^(a[81] & b[115])^(a[80] & b[116])^(a[79] & b[117])^(a[78] & b[118])^(a[77] & b[119])^(a[76] & b[120])^(a[75] & b[121])^(a[74] & b[122])^(a[73] & b[123])^(a[72] & b[124])^(a[71] & b[125])^(a[70] & b[126])^(a[69] & b[127])^(a[68] & b[128])^(a[67] & b[129])^(a[66] & b[130])^(a[65] & b[131])^(a[64] & b[132])^(a[63] & b[133])^(a[62] & b[134])^(a[61] & b[135])^(a[60] & b[136])^(a[59] & b[137])^(a[58] & b[138])^(a[57] & b[139])^(a[56] & b[140])^(a[55] & b[141])^(a[54] & b[142])^(a[53] & b[143])^(a[52] & b[144])^(a[51] & b[145])^(a[50] & b[146])^(a[49] & b[147])^(a[48] & b[148])^(a[47] & b[149])^(a[46] & b[150])^(a[45] & b[151])^(a[44] & b[152])^(a[43] & b[153])^(a[42] & b[154])^(a[41] & b[155])^(a[40] & b[156])^(a[39] & b[157])^(a[38] & b[158])^(a[37] & b[159])^(a[36] & b[160])^(a[35] & b[161])^(a[34] & b[162])^(a[33] & b[163])^(a[32] & b[164])^(a[31] & b[165])^(a[30] & b[166])^(a[29] & b[167])^(a[28] & b[168])^(a[27] & b[169])^(a[26] & b[170])^(a[25] & b[171])^(a[24] & b[172])^(a[23] & b[173])^(a[22] & b[174])^(a[21] & b[175])^(a[20] & b[176])^(a[19] & b[177])^(a[18] & b[178])^(a[17] & b[179])^(a[16] & b[180])^(a[15] & b[181])^(a[14] & b[182])^(a[13] & b[183])^(a[12] & b[184])^(a[11] & b[185])^(a[10] & b[186])^(a[9] & b[187])^(a[8] & b[188])^(a[7] & b[189])^(a[6] & b[190])^(a[5] & b[191])^(a[4] & b[192])^(a[3] & b[193])^(a[2] & b[194])^(a[1] & b[195])^(a[0] & b[196]);
assign y[197] = (a[197] & b[0])^(a[196] & b[1])^(a[195] & b[2])^(a[194] & b[3])^(a[193] & b[4])^(a[192] & b[5])^(a[191] & b[6])^(a[190] & b[7])^(a[189] & b[8])^(a[188] & b[9])^(a[187] & b[10])^(a[186] & b[11])^(a[185] & b[12])^(a[184] & b[13])^(a[183] & b[14])^(a[182] & b[15])^(a[181] & b[16])^(a[180] & b[17])^(a[179] & b[18])^(a[178] & b[19])^(a[177] & b[20])^(a[176] & b[21])^(a[175] & b[22])^(a[174] & b[23])^(a[173] & b[24])^(a[172] & b[25])^(a[171] & b[26])^(a[170] & b[27])^(a[169] & b[28])^(a[168] & b[29])^(a[167] & b[30])^(a[166] & b[31])^(a[165] & b[32])^(a[164] & b[33])^(a[163] & b[34])^(a[162] & b[35])^(a[161] & b[36])^(a[160] & b[37])^(a[159] & b[38])^(a[158] & b[39])^(a[157] & b[40])^(a[156] & b[41])^(a[155] & b[42])^(a[154] & b[43])^(a[153] & b[44])^(a[152] & b[45])^(a[151] & b[46])^(a[150] & b[47])^(a[149] & b[48])^(a[148] & b[49])^(a[147] & b[50])^(a[146] & b[51])^(a[145] & b[52])^(a[144] & b[53])^(a[143] & b[54])^(a[142] & b[55])^(a[141] & b[56])^(a[140] & b[57])^(a[139] & b[58])^(a[138] & b[59])^(a[137] & b[60])^(a[136] & b[61])^(a[135] & b[62])^(a[134] & b[63])^(a[133] & b[64])^(a[132] & b[65])^(a[131] & b[66])^(a[130] & b[67])^(a[129] & b[68])^(a[128] & b[69])^(a[127] & b[70])^(a[126] & b[71])^(a[125] & b[72])^(a[124] & b[73])^(a[123] & b[74])^(a[122] & b[75])^(a[121] & b[76])^(a[120] & b[77])^(a[119] & b[78])^(a[118] & b[79])^(a[117] & b[80])^(a[116] & b[81])^(a[115] & b[82])^(a[114] & b[83])^(a[113] & b[84])^(a[112] & b[85])^(a[111] & b[86])^(a[110] & b[87])^(a[109] & b[88])^(a[108] & b[89])^(a[107] & b[90])^(a[106] & b[91])^(a[105] & b[92])^(a[104] & b[93])^(a[103] & b[94])^(a[102] & b[95])^(a[101] & b[96])^(a[100] & b[97])^(a[99] & b[98])^(a[98] & b[99])^(a[97] & b[100])^(a[96] & b[101])^(a[95] & b[102])^(a[94] & b[103])^(a[93] & b[104])^(a[92] & b[105])^(a[91] & b[106])^(a[90] & b[107])^(a[89] & b[108])^(a[88] & b[109])^(a[87] & b[110])^(a[86] & b[111])^(a[85] & b[112])^(a[84] & b[113])^(a[83] & b[114])^(a[82] & b[115])^(a[81] & b[116])^(a[80] & b[117])^(a[79] & b[118])^(a[78] & b[119])^(a[77] & b[120])^(a[76] & b[121])^(a[75] & b[122])^(a[74] & b[123])^(a[73] & b[124])^(a[72] & b[125])^(a[71] & b[126])^(a[70] & b[127])^(a[69] & b[128])^(a[68] & b[129])^(a[67] & b[130])^(a[66] & b[131])^(a[65] & b[132])^(a[64] & b[133])^(a[63] & b[134])^(a[62] & b[135])^(a[61] & b[136])^(a[60] & b[137])^(a[59] & b[138])^(a[58] & b[139])^(a[57] & b[140])^(a[56] & b[141])^(a[55] & b[142])^(a[54] & b[143])^(a[53] & b[144])^(a[52] & b[145])^(a[51] & b[146])^(a[50] & b[147])^(a[49] & b[148])^(a[48] & b[149])^(a[47] & b[150])^(a[46] & b[151])^(a[45] & b[152])^(a[44] & b[153])^(a[43] & b[154])^(a[42] & b[155])^(a[41] & b[156])^(a[40] & b[157])^(a[39] & b[158])^(a[38] & b[159])^(a[37] & b[160])^(a[36] & b[161])^(a[35] & b[162])^(a[34] & b[163])^(a[33] & b[164])^(a[32] & b[165])^(a[31] & b[166])^(a[30] & b[167])^(a[29] & b[168])^(a[28] & b[169])^(a[27] & b[170])^(a[26] & b[171])^(a[25] & b[172])^(a[24] & b[173])^(a[23] & b[174])^(a[22] & b[175])^(a[21] & b[176])^(a[20] & b[177])^(a[19] & b[178])^(a[18] & b[179])^(a[17] & b[180])^(a[16] & b[181])^(a[15] & b[182])^(a[14] & b[183])^(a[13] & b[184])^(a[12] & b[185])^(a[11] & b[186])^(a[10] & b[187])^(a[9] & b[188])^(a[8] & b[189])^(a[7] & b[190])^(a[6] & b[191])^(a[5] & b[192])^(a[4] & b[193])^(a[3] & b[194])^(a[2] & b[195])^(a[1] & b[196])^(a[0] & b[197]);
assign y[198] = (a[198] & b[0])^(a[197] & b[1])^(a[196] & b[2])^(a[195] & b[3])^(a[194] & b[4])^(a[193] & b[5])^(a[192] & b[6])^(a[191] & b[7])^(a[190] & b[8])^(a[189] & b[9])^(a[188] & b[10])^(a[187] & b[11])^(a[186] & b[12])^(a[185] & b[13])^(a[184] & b[14])^(a[183] & b[15])^(a[182] & b[16])^(a[181] & b[17])^(a[180] & b[18])^(a[179] & b[19])^(a[178] & b[20])^(a[177] & b[21])^(a[176] & b[22])^(a[175] & b[23])^(a[174] & b[24])^(a[173] & b[25])^(a[172] & b[26])^(a[171] & b[27])^(a[170] & b[28])^(a[169] & b[29])^(a[168] & b[30])^(a[167] & b[31])^(a[166] & b[32])^(a[165] & b[33])^(a[164] & b[34])^(a[163] & b[35])^(a[162] & b[36])^(a[161] & b[37])^(a[160] & b[38])^(a[159] & b[39])^(a[158] & b[40])^(a[157] & b[41])^(a[156] & b[42])^(a[155] & b[43])^(a[154] & b[44])^(a[153] & b[45])^(a[152] & b[46])^(a[151] & b[47])^(a[150] & b[48])^(a[149] & b[49])^(a[148] & b[50])^(a[147] & b[51])^(a[146] & b[52])^(a[145] & b[53])^(a[144] & b[54])^(a[143] & b[55])^(a[142] & b[56])^(a[141] & b[57])^(a[140] & b[58])^(a[139] & b[59])^(a[138] & b[60])^(a[137] & b[61])^(a[136] & b[62])^(a[135] & b[63])^(a[134] & b[64])^(a[133] & b[65])^(a[132] & b[66])^(a[131] & b[67])^(a[130] & b[68])^(a[129] & b[69])^(a[128] & b[70])^(a[127] & b[71])^(a[126] & b[72])^(a[125] & b[73])^(a[124] & b[74])^(a[123] & b[75])^(a[122] & b[76])^(a[121] & b[77])^(a[120] & b[78])^(a[119] & b[79])^(a[118] & b[80])^(a[117] & b[81])^(a[116] & b[82])^(a[115] & b[83])^(a[114] & b[84])^(a[113] & b[85])^(a[112] & b[86])^(a[111] & b[87])^(a[110] & b[88])^(a[109] & b[89])^(a[108] & b[90])^(a[107] & b[91])^(a[106] & b[92])^(a[105] & b[93])^(a[104] & b[94])^(a[103] & b[95])^(a[102] & b[96])^(a[101] & b[97])^(a[100] & b[98])^(a[99] & b[99])^(a[98] & b[100])^(a[97] & b[101])^(a[96] & b[102])^(a[95] & b[103])^(a[94] & b[104])^(a[93] & b[105])^(a[92] & b[106])^(a[91] & b[107])^(a[90] & b[108])^(a[89] & b[109])^(a[88] & b[110])^(a[87] & b[111])^(a[86] & b[112])^(a[85] & b[113])^(a[84] & b[114])^(a[83] & b[115])^(a[82] & b[116])^(a[81] & b[117])^(a[80] & b[118])^(a[79] & b[119])^(a[78] & b[120])^(a[77] & b[121])^(a[76] & b[122])^(a[75] & b[123])^(a[74] & b[124])^(a[73] & b[125])^(a[72] & b[126])^(a[71] & b[127])^(a[70] & b[128])^(a[69] & b[129])^(a[68] & b[130])^(a[67] & b[131])^(a[66] & b[132])^(a[65] & b[133])^(a[64] & b[134])^(a[63] & b[135])^(a[62] & b[136])^(a[61] & b[137])^(a[60] & b[138])^(a[59] & b[139])^(a[58] & b[140])^(a[57] & b[141])^(a[56] & b[142])^(a[55] & b[143])^(a[54] & b[144])^(a[53] & b[145])^(a[52] & b[146])^(a[51] & b[147])^(a[50] & b[148])^(a[49] & b[149])^(a[48] & b[150])^(a[47] & b[151])^(a[46] & b[152])^(a[45] & b[153])^(a[44] & b[154])^(a[43] & b[155])^(a[42] & b[156])^(a[41] & b[157])^(a[40] & b[158])^(a[39] & b[159])^(a[38] & b[160])^(a[37] & b[161])^(a[36] & b[162])^(a[35] & b[163])^(a[34] & b[164])^(a[33] & b[165])^(a[32] & b[166])^(a[31] & b[167])^(a[30] & b[168])^(a[29] & b[169])^(a[28] & b[170])^(a[27] & b[171])^(a[26] & b[172])^(a[25] & b[173])^(a[24] & b[174])^(a[23] & b[175])^(a[22] & b[176])^(a[21] & b[177])^(a[20] & b[178])^(a[19] & b[179])^(a[18] & b[180])^(a[17] & b[181])^(a[16] & b[182])^(a[15] & b[183])^(a[14] & b[184])^(a[13] & b[185])^(a[12] & b[186])^(a[11] & b[187])^(a[10] & b[188])^(a[9] & b[189])^(a[8] & b[190])^(a[7] & b[191])^(a[6] & b[192])^(a[5] & b[193])^(a[4] & b[194])^(a[3] & b[195])^(a[2] & b[196])^(a[1] & b[197])^(a[0] & b[198]);
assign y[199] = (a[199] & b[0])^(a[198] & b[1])^(a[197] & b[2])^(a[196] & b[3])^(a[195] & b[4])^(a[194] & b[5])^(a[193] & b[6])^(a[192] & b[7])^(a[191] & b[8])^(a[190] & b[9])^(a[189] & b[10])^(a[188] & b[11])^(a[187] & b[12])^(a[186] & b[13])^(a[185] & b[14])^(a[184] & b[15])^(a[183] & b[16])^(a[182] & b[17])^(a[181] & b[18])^(a[180] & b[19])^(a[179] & b[20])^(a[178] & b[21])^(a[177] & b[22])^(a[176] & b[23])^(a[175] & b[24])^(a[174] & b[25])^(a[173] & b[26])^(a[172] & b[27])^(a[171] & b[28])^(a[170] & b[29])^(a[169] & b[30])^(a[168] & b[31])^(a[167] & b[32])^(a[166] & b[33])^(a[165] & b[34])^(a[164] & b[35])^(a[163] & b[36])^(a[162] & b[37])^(a[161] & b[38])^(a[160] & b[39])^(a[159] & b[40])^(a[158] & b[41])^(a[157] & b[42])^(a[156] & b[43])^(a[155] & b[44])^(a[154] & b[45])^(a[153] & b[46])^(a[152] & b[47])^(a[151] & b[48])^(a[150] & b[49])^(a[149] & b[50])^(a[148] & b[51])^(a[147] & b[52])^(a[146] & b[53])^(a[145] & b[54])^(a[144] & b[55])^(a[143] & b[56])^(a[142] & b[57])^(a[141] & b[58])^(a[140] & b[59])^(a[139] & b[60])^(a[138] & b[61])^(a[137] & b[62])^(a[136] & b[63])^(a[135] & b[64])^(a[134] & b[65])^(a[133] & b[66])^(a[132] & b[67])^(a[131] & b[68])^(a[130] & b[69])^(a[129] & b[70])^(a[128] & b[71])^(a[127] & b[72])^(a[126] & b[73])^(a[125] & b[74])^(a[124] & b[75])^(a[123] & b[76])^(a[122] & b[77])^(a[121] & b[78])^(a[120] & b[79])^(a[119] & b[80])^(a[118] & b[81])^(a[117] & b[82])^(a[116] & b[83])^(a[115] & b[84])^(a[114] & b[85])^(a[113] & b[86])^(a[112] & b[87])^(a[111] & b[88])^(a[110] & b[89])^(a[109] & b[90])^(a[108] & b[91])^(a[107] & b[92])^(a[106] & b[93])^(a[105] & b[94])^(a[104] & b[95])^(a[103] & b[96])^(a[102] & b[97])^(a[101] & b[98])^(a[100] & b[99])^(a[99] & b[100])^(a[98] & b[101])^(a[97] & b[102])^(a[96] & b[103])^(a[95] & b[104])^(a[94] & b[105])^(a[93] & b[106])^(a[92] & b[107])^(a[91] & b[108])^(a[90] & b[109])^(a[89] & b[110])^(a[88] & b[111])^(a[87] & b[112])^(a[86] & b[113])^(a[85] & b[114])^(a[84] & b[115])^(a[83] & b[116])^(a[82] & b[117])^(a[81] & b[118])^(a[80] & b[119])^(a[79] & b[120])^(a[78] & b[121])^(a[77] & b[122])^(a[76] & b[123])^(a[75] & b[124])^(a[74] & b[125])^(a[73] & b[126])^(a[72] & b[127])^(a[71] & b[128])^(a[70] & b[129])^(a[69] & b[130])^(a[68] & b[131])^(a[67] & b[132])^(a[66] & b[133])^(a[65] & b[134])^(a[64] & b[135])^(a[63] & b[136])^(a[62] & b[137])^(a[61] & b[138])^(a[60] & b[139])^(a[59] & b[140])^(a[58] & b[141])^(a[57] & b[142])^(a[56] & b[143])^(a[55] & b[144])^(a[54] & b[145])^(a[53] & b[146])^(a[52] & b[147])^(a[51] & b[148])^(a[50] & b[149])^(a[49] & b[150])^(a[48] & b[151])^(a[47] & b[152])^(a[46] & b[153])^(a[45] & b[154])^(a[44] & b[155])^(a[43] & b[156])^(a[42] & b[157])^(a[41] & b[158])^(a[40] & b[159])^(a[39] & b[160])^(a[38] & b[161])^(a[37] & b[162])^(a[36] & b[163])^(a[35] & b[164])^(a[34] & b[165])^(a[33] & b[166])^(a[32] & b[167])^(a[31] & b[168])^(a[30] & b[169])^(a[29] & b[170])^(a[28] & b[171])^(a[27] & b[172])^(a[26] & b[173])^(a[25] & b[174])^(a[24] & b[175])^(a[23] & b[176])^(a[22] & b[177])^(a[21] & b[178])^(a[20] & b[179])^(a[19] & b[180])^(a[18] & b[181])^(a[17] & b[182])^(a[16] & b[183])^(a[15] & b[184])^(a[14] & b[185])^(a[13] & b[186])^(a[12] & b[187])^(a[11] & b[188])^(a[10] & b[189])^(a[9] & b[190])^(a[8] & b[191])^(a[7] & b[192])^(a[6] & b[193])^(a[5] & b[194])^(a[4] & b[195])^(a[3] & b[196])^(a[2] & b[197])^(a[1] & b[198])^(a[0] & b[199]);
assign y[200] = (a[200] & b[0])^(a[199] & b[1])^(a[198] & b[2])^(a[197] & b[3])^(a[196] & b[4])^(a[195] & b[5])^(a[194] & b[6])^(a[193] & b[7])^(a[192] & b[8])^(a[191] & b[9])^(a[190] & b[10])^(a[189] & b[11])^(a[188] & b[12])^(a[187] & b[13])^(a[186] & b[14])^(a[185] & b[15])^(a[184] & b[16])^(a[183] & b[17])^(a[182] & b[18])^(a[181] & b[19])^(a[180] & b[20])^(a[179] & b[21])^(a[178] & b[22])^(a[177] & b[23])^(a[176] & b[24])^(a[175] & b[25])^(a[174] & b[26])^(a[173] & b[27])^(a[172] & b[28])^(a[171] & b[29])^(a[170] & b[30])^(a[169] & b[31])^(a[168] & b[32])^(a[167] & b[33])^(a[166] & b[34])^(a[165] & b[35])^(a[164] & b[36])^(a[163] & b[37])^(a[162] & b[38])^(a[161] & b[39])^(a[160] & b[40])^(a[159] & b[41])^(a[158] & b[42])^(a[157] & b[43])^(a[156] & b[44])^(a[155] & b[45])^(a[154] & b[46])^(a[153] & b[47])^(a[152] & b[48])^(a[151] & b[49])^(a[150] & b[50])^(a[149] & b[51])^(a[148] & b[52])^(a[147] & b[53])^(a[146] & b[54])^(a[145] & b[55])^(a[144] & b[56])^(a[143] & b[57])^(a[142] & b[58])^(a[141] & b[59])^(a[140] & b[60])^(a[139] & b[61])^(a[138] & b[62])^(a[137] & b[63])^(a[136] & b[64])^(a[135] & b[65])^(a[134] & b[66])^(a[133] & b[67])^(a[132] & b[68])^(a[131] & b[69])^(a[130] & b[70])^(a[129] & b[71])^(a[128] & b[72])^(a[127] & b[73])^(a[126] & b[74])^(a[125] & b[75])^(a[124] & b[76])^(a[123] & b[77])^(a[122] & b[78])^(a[121] & b[79])^(a[120] & b[80])^(a[119] & b[81])^(a[118] & b[82])^(a[117] & b[83])^(a[116] & b[84])^(a[115] & b[85])^(a[114] & b[86])^(a[113] & b[87])^(a[112] & b[88])^(a[111] & b[89])^(a[110] & b[90])^(a[109] & b[91])^(a[108] & b[92])^(a[107] & b[93])^(a[106] & b[94])^(a[105] & b[95])^(a[104] & b[96])^(a[103] & b[97])^(a[102] & b[98])^(a[101] & b[99])^(a[100] & b[100])^(a[99] & b[101])^(a[98] & b[102])^(a[97] & b[103])^(a[96] & b[104])^(a[95] & b[105])^(a[94] & b[106])^(a[93] & b[107])^(a[92] & b[108])^(a[91] & b[109])^(a[90] & b[110])^(a[89] & b[111])^(a[88] & b[112])^(a[87] & b[113])^(a[86] & b[114])^(a[85] & b[115])^(a[84] & b[116])^(a[83] & b[117])^(a[82] & b[118])^(a[81] & b[119])^(a[80] & b[120])^(a[79] & b[121])^(a[78] & b[122])^(a[77] & b[123])^(a[76] & b[124])^(a[75] & b[125])^(a[74] & b[126])^(a[73] & b[127])^(a[72] & b[128])^(a[71] & b[129])^(a[70] & b[130])^(a[69] & b[131])^(a[68] & b[132])^(a[67] & b[133])^(a[66] & b[134])^(a[65] & b[135])^(a[64] & b[136])^(a[63] & b[137])^(a[62] & b[138])^(a[61] & b[139])^(a[60] & b[140])^(a[59] & b[141])^(a[58] & b[142])^(a[57] & b[143])^(a[56] & b[144])^(a[55] & b[145])^(a[54] & b[146])^(a[53] & b[147])^(a[52] & b[148])^(a[51] & b[149])^(a[50] & b[150])^(a[49] & b[151])^(a[48] & b[152])^(a[47] & b[153])^(a[46] & b[154])^(a[45] & b[155])^(a[44] & b[156])^(a[43] & b[157])^(a[42] & b[158])^(a[41] & b[159])^(a[40] & b[160])^(a[39] & b[161])^(a[38] & b[162])^(a[37] & b[163])^(a[36] & b[164])^(a[35] & b[165])^(a[34] & b[166])^(a[33] & b[167])^(a[32] & b[168])^(a[31] & b[169])^(a[30] & b[170])^(a[29] & b[171])^(a[28] & b[172])^(a[27] & b[173])^(a[26] & b[174])^(a[25] & b[175])^(a[24] & b[176])^(a[23] & b[177])^(a[22] & b[178])^(a[21] & b[179])^(a[20] & b[180])^(a[19] & b[181])^(a[18] & b[182])^(a[17] & b[183])^(a[16] & b[184])^(a[15] & b[185])^(a[14] & b[186])^(a[13] & b[187])^(a[12] & b[188])^(a[11] & b[189])^(a[10] & b[190])^(a[9] & b[191])^(a[8] & b[192])^(a[7] & b[193])^(a[6] & b[194])^(a[5] & b[195])^(a[4] & b[196])^(a[3] & b[197])^(a[2] & b[198])^(a[1] & b[199])^(a[0] & b[200]);
assign y[201] = (a[201] & b[0])^(a[200] & b[1])^(a[199] & b[2])^(a[198] & b[3])^(a[197] & b[4])^(a[196] & b[5])^(a[195] & b[6])^(a[194] & b[7])^(a[193] & b[8])^(a[192] & b[9])^(a[191] & b[10])^(a[190] & b[11])^(a[189] & b[12])^(a[188] & b[13])^(a[187] & b[14])^(a[186] & b[15])^(a[185] & b[16])^(a[184] & b[17])^(a[183] & b[18])^(a[182] & b[19])^(a[181] & b[20])^(a[180] & b[21])^(a[179] & b[22])^(a[178] & b[23])^(a[177] & b[24])^(a[176] & b[25])^(a[175] & b[26])^(a[174] & b[27])^(a[173] & b[28])^(a[172] & b[29])^(a[171] & b[30])^(a[170] & b[31])^(a[169] & b[32])^(a[168] & b[33])^(a[167] & b[34])^(a[166] & b[35])^(a[165] & b[36])^(a[164] & b[37])^(a[163] & b[38])^(a[162] & b[39])^(a[161] & b[40])^(a[160] & b[41])^(a[159] & b[42])^(a[158] & b[43])^(a[157] & b[44])^(a[156] & b[45])^(a[155] & b[46])^(a[154] & b[47])^(a[153] & b[48])^(a[152] & b[49])^(a[151] & b[50])^(a[150] & b[51])^(a[149] & b[52])^(a[148] & b[53])^(a[147] & b[54])^(a[146] & b[55])^(a[145] & b[56])^(a[144] & b[57])^(a[143] & b[58])^(a[142] & b[59])^(a[141] & b[60])^(a[140] & b[61])^(a[139] & b[62])^(a[138] & b[63])^(a[137] & b[64])^(a[136] & b[65])^(a[135] & b[66])^(a[134] & b[67])^(a[133] & b[68])^(a[132] & b[69])^(a[131] & b[70])^(a[130] & b[71])^(a[129] & b[72])^(a[128] & b[73])^(a[127] & b[74])^(a[126] & b[75])^(a[125] & b[76])^(a[124] & b[77])^(a[123] & b[78])^(a[122] & b[79])^(a[121] & b[80])^(a[120] & b[81])^(a[119] & b[82])^(a[118] & b[83])^(a[117] & b[84])^(a[116] & b[85])^(a[115] & b[86])^(a[114] & b[87])^(a[113] & b[88])^(a[112] & b[89])^(a[111] & b[90])^(a[110] & b[91])^(a[109] & b[92])^(a[108] & b[93])^(a[107] & b[94])^(a[106] & b[95])^(a[105] & b[96])^(a[104] & b[97])^(a[103] & b[98])^(a[102] & b[99])^(a[101] & b[100])^(a[100] & b[101])^(a[99] & b[102])^(a[98] & b[103])^(a[97] & b[104])^(a[96] & b[105])^(a[95] & b[106])^(a[94] & b[107])^(a[93] & b[108])^(a[92] & b[109])^(a[91] & b[110])^(a[90] & b[111])^(a[89] & b[112])^(a[88] & b[113])^(a[87] & b[114])^(a[86] & b[115])^(a[85] & b[116])^(a[84] & b[117])^(a[83] & b[118])^(a[82] & b[119])^(a[81] & b[120])^(a[80] & b[121])^(a[79] & b[122])^(a[78] & b[123])^(a[77] & b[124])^(a[76] & b[125])^(a[75] & b[126])^(a[74] & b[127])^(a[73] & b[128])^(a[72] & b[129])^(a[71] & b[130])^(a[70] & b[131])^(a[69] & b[132])^(a[68] & b[133])^(a[67] & b[134])^(a[66] & b[135])^(a[65] & b[136])^(a[64] & b[137])^(a[63] & b[138])^(a[62] & b[139])^(a[61] & b[140])^(a[60] & b[141])^(a[59] & b[142])^(a[58] & b[143])^(a[57] & b[144])^(a[56] & b[145])^(a[55] & b[146])^(a[54] & b[147])^(a[53] & b[148])^(a[52] & b[149])^(a[51] & b[150])^(a[50] & b[151])^(a[49] & b[152])^(a[48] & b[153])^(a[47] & b[154])^(a[46] & b[155])^(a[45] & b[156])^(a[44] & b[157])^(a[43] & b[158])^(a[42] & b[159])^(a[41] & b[160])^(a[40] & b[161])^(a[39] & b[162])^(a[38] & b[163])^(a[37] & b[164])^(a[36] & b[165])^(a[35] & b[166])^(a[34] & b[167])^(a[33] & b[168])^(a[32] & b[169])^(a[31] & b[170])^(a[30] & b[171])^(a[29] & b[172])^(a[28] & b[173])^(a[27] & b[174])^(a[26] & b[175])^(a[25] & b[176])^(a[24] & b[177])^(a[23] & b[178])^(a[22] & b[179])^(a[21] & b[180])^(a[20] & b[181])^(a[19] & b[182])^(a[18] & b[183])^(a[17] & b[184])^(a[16] & b[185])^(a[15] & b[186])^(a[14] & b[187])^(a[13] & b[188])^(a[12] & b[189])^(a[11] & b[190])^(a[10] & b[191])^(a[9] & b[192])^(a[8] & b[193])^(a[7] & b[194])^(a[6] & b[195])^(a[5] & b[196])^(a[4] & b[197])^(a[3] & b[198])^(a[2] & b[199])^(a[1] & b[200])^(a[0] & b[201]);
assign y[202] = (a[202] & b[0])^(a[201] & b[1])^(a[200] & b[2])^(a[199] & b[3])^(a[198] & b[4])^(a[197] & b[5])^(a[196] & b[6])^(a[195] & b[7])^(a[194] & b[8])^(a[193] & b[9])^(a[192] & b[10])^(a[191] & b[11])^(a[190] & b[12])^(a[189] & b[13])^(a[188] & b[14])^(a[187] & b[15])^(a[186] & b[16])^(a[185] & b[17])^(a[184] & b[18])^(a[183] & b[19])^(a[182] & b[20])^(a[181] & b[21])^(a[180] & b[22])^(a[179] & b[23])^(a[178] & b[24])^(a[177] & b[25])^(a[176] & b[26])^(a[175] & b[27])^(a[174] & b[28])^(a[173] & b[29])^(a[172] & b[30])^(a[171] & b[31])^(a[170] & b[32])^(a[169] & b[33])^(a[168] & b[34])^(a[167] & b[35])^(a[166] & b[36])^(a[165] & b[37])^(a[164] & b[38])^(a[163] & b[39])^(a[162] & b[40])^(a[161] & b[41])^(a[160] & b[42])^(a[159] & b[43])^(a[158] & b[44])^(a[157] & b[45])^(a[156] & b[46])^(a[155] & b[47])^(a[154] & b[48])^(a[153] & b[49])^(a[152] & b[50])^(a[151] & b[51])^(a[150] & b[52])^(a[149] & b[53])^(a[148] & b[54])^(a[147] & b[55])^(a[146] & b[56])^(a[145] & b[57])^(a[144] & b[58])^(a[143] & b[59])^(a[142] & b[60])^(a[141] & b[61])^(a[140] & b[62])^(a[139] & b[63])^(a[138] & b[64])^(a[137] & b[65])^(a[136] & b[66])^(a[135] & b[67])^(a[134] & b[68])^(a[133] & b[69])^(a[132] & b[70])^(a[131] & b[71])^(a[130] & b[72])^(a[129] & b[73])^(a[128] & b[74])^(a[127] & b[75])^(a[126] & b[76])^(a[125] & b[77])^(a[124] & b[78])^(a[123] & b[79])^(a[122] & b[80])^(a[121] & b[81])^(a[120] & b[82])^(a[119] & b[83])^(a[118] & b[84])^(a[117] & b[85])^(a[116] & b[86])^(a[115] & b[87])^(a[114] & b[88])^(a[113] & b[89])^(a[112] & b[90])^(a[111] & b[91])^(a[110] & b[92])^(a[109] & b[93])^(a[108] & b[94])^(a[107] & b[95])^(a[106] & b[96])^(a[105] & b[97])^(a[104] & b[98])^(a[103] & b[99])^(a[102] & b[100])^(a[101] & b[101])^(a[100] & b[102])^(a[99] & b[103])^(a[98] & b[104])^(a[97] & b[105])^(a[96] & b[106])^(a[95] & b[107])^(a[94] & b[108])^(a[93] & b[109])^(a[92] & b[110])^(a[91] & b[111])^(a[90] & b[112])^(a[89] & b[113])^(a[88] & b[114])^(a[87] & b[115])^(a[86] & b[116])^(a[85] & b[117])^(a[84] & b[118])^(a[83] & b[119])^(a[82] & b[120])^(a[81] & b[121])^(a[80] & b[122])^(a[79] & b[123])^(a[78] & b[124])^(a[77] & b[125])^(a[76] & b[126])^(a[75] & b[127])^(a[74] & b[128])^(a[73] & b[129])^(a[72] & b[130])^(a[71] & b[131])^(a[70] & b[132])^(a[69] & b[133])^(a[68] & b[134])^(a[67] & b[135])^(a[66] & b[136])^(a[65] & b[137])^(a[64] & b[138])^(a[63] & b[139])^(a[62] & b[140])^(a[61] & b[141])^(a[60] & b[142])^(a[59] & b[143])^(a[58] & b[144])^(a[57] & b[145])^(a[56] & b[146])^(a[55] & b[147])^(a[54] & b[148])^(a[53] & b[149])^(a[52] & b[150])^(a[51] & b[151])^(a[50] & b[152])^(a[49] & b[153])^(a[48] & b[154])^(a[47] & b[155])^(a[46] & b[156])^(a[45] & b[157])^(a[44] & b[158])^(a[43] & b[159])^(a[42] & b[160])^(a[41] & b[161])^(a[40] & b[162])^(a[39] & b[163])^(a[38] & b[164])^(a[37] & b[165])^(a[36] & b[166])^(a[35] & b[167])^(a[34] & b[168])^(a[33] & b[169])^(a[32] & b[170])^(a[31] & b[171])^(a[30] & b[172])^(a[29] & b[173])^(a[28] & b[174])^(a[27] & b[175])^(a[26] & b[176])^(a[25] & b[177])^(a[24] & b[178])^(a[23] & b[179])^(a[22] & b[180])^(a[21] & b[181])^(a[20] & b[182])^(a[19] & b[183])^(a[18] & b[184])^(a[17] & b[185])^(a[16] & b[186])^(a[15] & b[187])^(a[14] & b[188])^(a[13] & b[189])^(a[12] & b[190])^(a[11] & b[191])^(a[10] & b[192])^(a[9] & b[193])^(a[8] & b[194])^(a[7] & b[195])^(a[6] & b[196])^(a[5] & b[197])^(a[4] & b[198])^(a[3] & b[199])^(a[2] & b[200])^(a[1] & b[201])^(a[0] & b[202]);
assign y[203] = (a[203] & b[0])^(a[202] & b[1])^(a[201] & b[2])^(a[200] & b[3])^(a[199] & b[4])^(a[198] & b[5])^(a[197] & b[6])^(a[196] & b[7])^(a[195] & b[8])^(a[194] & b[9])^(a[193] & b[10])^(a[192] & b[11])^(a[191] & b[12])^(a[190] & b[13])^(a[189] & b[14])^(a[188] & b[15])^(a[187] & b[16])^(a[186] & b[17])^(a[185] & b[18])^(a[184] & b[19])^(a[183] & b[20])^(a[182] & b[21])^(a[181] & b[22])^(a[180] & b[23])^(a[179] & b[24])^(a[178] & b[25])^(a[177] & b[26])^(a[176] & b[27])^(a[175] & b[28])^(a[174] & b[29])^(a[173] & b[30])^(a[172] & b[31])^(a[171] & b[32])^(a[170] & b[33])^(a[169] & b[34])^(a[168] & b[35])^(a[167] & b[36])^(a[166] & b[37])^(a[165] & b[38])^(a[164] & b[39])^(a[163] & b[40])^(a[162] & b[41])^(a[161] & b[42])^(a[160] & b[43])^(a[159] & b[44])^(a[158] & b[45])^(a[157] & b[46])^(a[156] & b[47])^(a[155] & b[48])^(a[154] & b[49])^(a[153] & b[50])^(a[152] & b[51])^(a[151] & b[52])^(a[150] & b[53])^(a[149] & b[54])^(a[148] & b[55])^(a[147] & b[56])^(a[146] & b[57])^(a[145] & b[58])^(a[144] & b[59])^(a[143] & b[60])^(a[142] & b[61])^(a[141] & b[62])^(a[140] & b[63])^(a[139] & b[64])^(a[138] & b[65])^(a[137] & b[66])^(a[136] & b[67])^(a[135] & b[68])^(a[134] & b[69])^(a[133] & b[70])^(a[132] & b[71])^(a[131] & b[72])^(a[130] & b[73])^(a[129] & b[74])^(a[128] & b[75])^(a[127] & b[76])^(a[126] & b[77])^(a[125] & b[78])^(a[124] & b[79])^(a[123] & b[80])^(a[122] & b[81])^(a[121] & b[82])^(a[120] & b[83])^(a[119] & b[84])^(a[118] & b[85])^(a[117] & b[86])^(a[116] & b[87])^(a[115] & b[88])^(a[114] & b[89])^(a[113] & b[90])^(a[112] & b[91])^(a[111] & b[92])^(a[110] & b[93])^(a[109] & b[94])^(a[108] & b[95])^(a[107] & b[96])^(a[106] & b[97])^(a[105] & b[98])^(a[104] & b[99])^(a[103] & b[100])^(a[102] & b[101])^(a[101] & b[102])^(a[100] & b[103])^(a[99] & b[104])^(a[98] & b[105])^(a[97] & b[106])^(a[96] & b[107])^(a[95] & b[108])^(a[94] & b[109])^(a[93] & b[110])^(a[92] & b[111])^(a[91] & b[112])^(a[90] & b[113])^(a[89] & b[114])^(a[88] & b[115])^(a[87] & b[116])^(a[86] & b[117])^(a[85] & b[118])^(a[84] & b[119])^(a[83] & b[120])^(a[82] & b[121])^(a[81] & b[122])^(a[80] & b[123])^(a[79] & b[124])^(a[78] & b[125])^(a[77] & b[126])^(a[76] & b[127])^(a[75] & b[128])^(a[74] & b[129])^(a[73] & b[130])^(a[72] & b[131])^(a[71] & b[132])^(a[70] & b[133])^(a[69] & b[134])^(a[68] & b[135])^(a[67] & b[136])^(a[66] & b[137])^(a[65] & b[138])^(a[64] & b[139])^(a[63] & b[140])^(a[62] & b[141])^(a[61] & b[142])^(a[60] & b[143])^(a[59] & b[144])^(a[58] & b[145])^(a[57] & b[146])^(a[56] & b[147])^(a[55] & b[148])^(a[54] & b[149])^(a[53] & b[150])^(a[52] & b[151])^(a[51] & b[152])^(a[50] & b[153])^(a[49] & b[154])^(a[48] & b[155])^(a[47] & b[156])^(a[46] & b[157])^(a[45] & b[158])^(a[44] & b[159])^(a[43] & b[160])^(a[42] & b[161])^(a[41] & b[162])^(a[40] & b[163])^(a[39] & b[164])^(a[38] & b[165])^(a[37] & b[166])^(a[36] & b[167])^(a[35] & b[168])^(a[34] & b[169])^(a[33] & b[170])^(a[32] & b[171])^(a[31] & b[172])^(a[30] & b[173])^(a[29] & b[174])^(a[28] & b[175])^(a[27] & b[176])^(a[26] & b[177])^(a[25] & b[178])^(a[24] & b[179])^(a[23] & b[180])^(a[22] & b[181])^(a[21] & b[182])^(a[20] & b[183])^(a[19] & b[184])^(a[18] & b[185])^(a[17] & b[186])^(a[16] & b[187])^(a[15] & b[188])^(a[14] & b[189])^(a[13] & b[190])^(a[12] & b[191])^(a[11] & b[192])^(a[10] & b[193])^(a[9] & b[194])^(a[8] & b[195])^(a[7] & b[196])^(a[6] & b[197])^(a[5] & b[198])^(a[4] & b[199])^(a[3] & b[200])^(a[2] & b[201])^(a[1] & b[202])^(a[0] & b[203]);
assign y[204] = (a[204] & b[0])^(a[203] & b[1])^(a[202] & b[2])^(a[201] & b[3])^(a[200] & b[4])^(a[199] & b[5])^(a[198] & b[6])^(a[197] & b[7])^(a[196] & b[8])^(a[195] & b[9])^(a[194] & b[10])^(a[193] & b[11])^(a[192] & b[12])^(a[191] & b[13])^(a[190] & b[14])^(a[189] & b[15])^(a[188] & b[16])^(a[187] & b[17])^(a[186] & b[18])^(a[185] & b[19])^(a[184] & b[20])^(a[183] & b[21])^(a[182] & b[22])^(a[181] & b[23])^(a[180] & b[24])^(a[179] & b[25])^(a[178] & b[26])^(a[177] & b[27])^(a[176] & b[28])^(a[175] & b[29])^(a[174] & b[30])^(a[173] & b[31])^(a[172] & b[32])^(a[171] & b[33])^(a[170] & b[34])^(a[169] & b[35])^(a[168] & b[36])^(a[167] & b[37])^(a[166] & b[38])^(a[165] & b[39])^(a[164] & b[40])^(a[163] & b[41])^(a[162] & b[42])^(a[161] & b[43])^(a[160] & b[44])^(a[159] & b[45])^(a[158] & b[46])^(a[157] & b[47])^(a[156] & b[48])^(a[155] & b[49])^(a[154] & b[50])^(a[153] & b[51])^(a[152] & b[52])^(a[151] & b[53])^(a[150] & b[54])^(a[149] & b[55])^(a[148] & b[56])^(a[147] & b[57])^(a[146] & b[58])^(a[145] & b[59])^(a[144] & b[60])^(a[143] & b[61])^(a[142] & b[62])^(a[141] & b[63])^(a[140] & b[64])^(a[139] & b[65])^(a[138] & b[66])^(a[137] & b[67])^(a[136] & b[68])^(a[135] & b[69])^(a[134] & b[70])^(a[133] & b[71])^(a[132] & b[72])^(a[131] & b[73])^(a[130] & b[74])^(a[129] & b[75])^(a[128] & b[76])^(a[127] & b[77])^(a[126] & b[78])^(a[125] & b[79])^(a[124] & b[80])^(a[123] & b[81])^(a[122] & b[82])^(a[121] & b[83])^(a[120] & b[84])^(a[119] & b[85])^(a[118] & b[86])^(a[117] & b[87])^(a[116] & b[88])^(a[115] & b[89])^(a[114] & b[90])^(a[113] & b[91])^(a[112] & b[92])^(a[111] & b[93])^(a[110] & b[94])^(a[109] & b[95])^(a[108] & b[96])^(a[107] & b[97])^(a[106] & b[98])^(a[105] & b[99])^(a[104] & b[100])^(a[103] & b[101])^(a[102] & b[102])^(a[101] & b[103])^(a[100] & b[104])^(a[99] & b[105])^(a[98] & b[106])^(a[97] & b[107])^(a[96] & b[108])^(a[95] & b[109])^(a[94] & b[110])^(a[93] & b[111])^(a[92] & b[112])^(a[91] & b[113])^(a[90] & b[114])^(a[89] & b[115])^(a[88] & b[116])^(a[87] & b[117])^(a[86] & b[118])^(a[85] & b[119])^(a[84] & b[120])^(a[83] & b[121])^(a[82] & b[122])^(a[81] & b[123])^(a[80] & b[124])^(a[79] & b[125])^(a[78] & b[126])^(a[77] & b[127])^(a[76] & b[128])^(a[75] & b[129])^(a[74] & b[130])^(a[73] & b[131])^(a[72] & b[132])^(a[71] & b[133])^(a[70] & b[134])^(a[69] & b[135])^(a[68] & b[136])^(a[67] & b[137])^(a[66] & b[138])^(a[65] & b[139])^(a[64] & b[140])^(a[63] & b[141])^(a[62] & b[142])^(a[61] & b[143])^(a[60] & b[144])^(a[59] & b[145])^(a[58] & b[146])^(a[57] & b[147])^(a[56] & b[148])^(a[55] & b[149])^(a[54] & b[150])^(a[53] & b[151])^(a[52] & b[152])^(a[51] & b[153])^(a[50] & b[154])^(a[49] & b[155])^(a[48] & b[156])^(a[47] & b[157])^(a[46] & b[158])^(a[45] & b[159])^(a[44] & b[160])^(a[43] & b[161])^(a[42] & b[162])^(a[41] & b[163])^(a[40] & b[164])^(a[39] & b[165])^(a[38] & b[166])^(a[37] & b[167])^(a[36] & b[168])^(a[35] & b[169])^(a[34] & b[170])^(a[33] & b[171])^(a[32] & b[172])^(a[31] & b[173])^(a[30] & b[174])^(a[29] & b[175])^(a[28] & b[176])^(a[27] & b[177])^(a[26] & b[178])^(a[25] & b[179])^(a[24] & b[180])^(a[23] & b[181])^(a[22] & b[182])^(a[21] & b[183])^(a[20] & b[184])^(a[19] & b[185])^(a[18] & b[186])^(a[17] & b[187])^(a[16] & b[188])^(a[15] & b[189])^(a[14] & b[190])^(a[13] & b[191])^(a[12] & b[192])^(a[11] & b[193])^(a[10] & b[194])^(a[9] & b[195])^(a[8] & b[196])^(a[7] & b[197])^(a[6] & b[198])^(a[5] & b[199])^(a[4] & b[200])^(a[3] & b[201])^(a[2] & b[202])^(a[1] & b[203])^(a[0] & b[204]);
assign y[205] = (a[205] & b[0])^(a[204] & b[1])^(a[203] & b[2])^(a[202] & b[3])^(a[201] & b[4])^(a[200] & b[5])^(a[199] & b[6])^(a[198] & b[7])^(a[197] & b[8])^(a[196] & b[9])^(a[195] & b[10])^(a[194] & b[11])^(a[193] & b[12])^(a[192] & b[13])^(a[191] & b[14])^(a[190] & b[15])^(a[189] & b[16])^(a[188] & b[17])^(a[187] & b[18])^(a[186] & b[19])^(a[185] & b[20])^(a[184] & b[21])^(a[183] & b[22])^(a[182] & b[23])^(a[181] & b[24])^(a[180] & b[25])^(a[179] & b[26])^(a[178] & b[27])^(a[177] & b[28])^(a[176] & b[29])^(a[175] & b[30])^(a[174] & b[31])^(a[173] & b[32])^(a[172] & b[33])^(a[171] & b[34])^(a[170] & b[35])^(a[169] & b[36])^(a[168] & b[37])^(a[167] & b[38])^(a[166] & b[39])^(a[165] & b[40])^(a[164] & b[41])^(a[163] & b[42])^(a[162] & b[43])^(a[161] & b[44])^(a[160] & b[45])^(a[159] & b[46])^(a[158] & b[47])^(a[157] & b[48])^(a[156] & b[49])^(a[155] & b[50])^(a[154] & b[51])^(a[153] & b[52])^(a[152] & b[53])^(a[151] & b[54])^(a[150] & b[55])^(a[149] & b[56])^(a[148] & b[57])^(a[147] & b[58])^(a[146] & b[59])^(a[145] & b[60])^(a[144] & b[61])^(a[143] & b[62])^(a[142] & b[63])^(a[141] & b[64])^(a[140] & b[65])^(a[139] & b[66])^(a[138] & b[67])^(a[137] & b[68])^(a[136] & b[69])^(a[135] & b[70])^(a[134] & b[71])^(a[133] & b[72])^(a[132] & b[73])^(a[131] & b[74])^(a[130] & b[75])^(a[129] & b[76])^(a[128] & b[77])^(a[127] & b[78])^(a[126] & b[79])^(a[125] & b[80])^(a[124] & b[81])^(a[123] & b[82])^(a[122] & b[83])^(a[121] & b[84])^(a[120] & b[85])^(a[119] & b[86])^(a[118] & b[87])^(a[117] & b[88])^(a[116] & b[89])^(a[115] & b[90])^(a[114] & b[91])^(a[113] & b[92])^(a[112] & b[93])^(a[111] & b[94])^(a[110] & b[95])^(a[109] & b[96])^(a[108] & b[97])^(a[107] & b[98])^(a[106] & b[99])^(a[105] & b[100])^(a[104] & b[101])^(a[103] & b[102])^(a[102] & b[103])^(a[101] & b[104])^(a[100] & b[105])^(a[99] & b[106])^(a[98] & b[107])^(a[97] & b[108])^(a[96] & b[109])^(a[95] & b[110])^(a[94] & b[111])^(a[93] & b[112])^(a[92] & b[113])^(a[91] & b[114])^(a[90] & b[115])^(a[89] & b[116])^(a[88] & b[117])^(a[87] & b[118])^(a[86] & b[119])^(a[85] & b[120])^(a[84] & b[121])^(a[83] & b[122])^(a[82] & b[123])^(a[81] & b[124])^(a[80] & b[125])^(a[79] & b[126])^(a[78] & b[127])^(a[77] & b[128])^(a[76] & b[129])^(a[75] & b[130])^(a[74] & b[131])^(a[73] & b[132])^(a[72] & b[133])^(a[71] & b[134])^(a[70] & b[135])^(a[69] & b[136])^(a[68] & b[137])^(a[67] & b[138])^(a[66] & b[139])^(a[65] & b[140])^(a[64] & b[141])^(a[63] & b[142])^(a[62] & b[143])^(a[61] & b[144])^(a[60] & b[145])^(a[59] & b[146])^(a[58] & b[147])^(a[57] & b[148])^(a[56] & b[149])^(a[55] & b[150])^(a[54] & b[151])^(a[53] & b[152])^(a[52] & b[153])^(a[51] & b[154])^(a[50] & b[155])^(a[49] & b[156])^(a[48] & b[157])^(a[47] & b[158])^(a[46] & b[159])^(a[45] & b[160])^(a[44] & b[161])^(a[43] & b[162])^(a[42] & b[163])^(a[41] & b[164])^(a[40] & b[165])^(a[39] & b[166])^(a[38] & b[167])^(a[37] & b[168])^(a[36] & b[169])^(a[35] & b[170])^(a[34] & b[171])^(a[33] & b[172])^(a[32] & b[173])^(a[31] & b[174])^(a[30] & b[175])^(a[29] & b[176])^(a[28] & b[177])^(a[27] & b[178])^(a[26] & b[179])^(a[25] & b[180])^(a[24] & b[181])^(a[23] & b[182])^(a[22] & b[183])^(a[21] & b[184])^(a[20] & b[185])^(a[19] & b[186])^(a[18] & b[187])^(a[17] & b[188])^(a[16] & b[189])^(a[15] & b[190])^(a[14] & b[191])^(a[13] & b[192])^(a[12] & b[193])^(a[11] & b[194])^(a[10] & b[195])^(a[9] & b[196])^(a[8] & b[197])^(a[7] & b[198])^(a[6] & b[199])^(a[5] & b[200])^(a[4] & b[201])^(a[3] & b[202])^(a[2] & b[203])^(a[1] & b[204])^(a[0] & b[205]);
assign y[206] = (a[206] & b[0])^(a[205] & b[1])^(a[204] & b[2])^(a[203] & b[3])^(a[202] & b[4])^(a[201] & b[5])^(a[200] & b[6])^(a[199] & b[7])^(a[198] & b[8])^(a[197] & b[9])^(a[196] & b[10])^(a[195] & b[11])^(a[194] & b[12])^(a[193] & b[13])^(a[192] & b[14])^(a[191] & b[15])^(a[190] & b[16])^(a[189] & b[17])^(a[188] & b[18])^(a[187] & b[19])^(a[186] & b[20])^(a[185] & b[21])^(a[184] & b[22])^(a[183] & b[23])^(a[182] & b[24])^(a[181] & b[25])^(a[180] & b[26])^(a[179] & b[27])^(a[178] & b[28])^(a[177] & b[29])^(a[176] & b[30])^(a[175] & b[31])^(a[174] & b[32])^(a[173] & b[33])^(a[172] & b[34])^(a[171] & b[35])^(a[170] & b[36])^(a[169] & b[37])^(a[168] & b[38])^(a[167] & b[39])^(a[166] & b[40])^(a[165] & b[41])^(a[164] & b[42])^(a[163] & b[43])^(a[162] & b[44])^(a[161] & b[45])^(a[160] & b[46])^(a[159] & b[47])^(a[158] & b[48])^(a[157] & b[49])^(a[156] & b[50])^(a[155] & b[51])^(a[154] & b[52])^(a[153] & b[53])^(a[152] & b[54])^(a[151] & b[55])^(a[150] & b[56])^(a[149] & b[57])^(a[148] & b[58])^(a[147] & b[59])^(a[146] & b[60])^(a[145] & b[61])^(a[144] & b[62])^(a[143] & b[63])^(a[142] & b[64])^(a[141] & b[65])^(a[140] & b[66])^(a[139] & b[67])^(a[138] & b[68])^(a[137] & b[69])^(a[136] & b[70])^(a[135] & b[71])^(a[134] & b[72])^(a[133] & b[73])^(a[132] & b[74])^(a[131] & b[75])^(a[130] & b[76])^(a[129] & b[77])^(a[128] & b[78])^(a[127] & b[79])^(a[126] & b[80])^(a[125] & b[81])^(a[124] & b[82])^(a[123] & b[83])^(a[122] & b[84])^(a[121] & b[85])^(a[120] & b[86])^(a[119] & b[87])^(a[118] & b[88])^(a[117] & b[89])^(a[116] & b[90])^(a[115] & b[91])^(a[114] & b[92])^(a[113] & b[93])^(a[112] & b[94])^(a[111] & b[95])^(a[110] & b[96])^(a[109] & b[97])^(a[108] & b[98])^(a[107] & b[99])^(a[106] & b[100])^(a[105] & b[101])^(a[104] & b[102])^(a[103] & b[103])^(a[102] & b[104])^(a[101] & b[105])^(a[100] & b[106])^(a[99] & b[107])^(a[98] & b[108])^(a[97] & b[109])^(a[96] & b[110])^(a[95] & b[111])^(a[94] & b[112])^(a[93] & b[113])^(a[92] & b[114])^(a[91] & b[115])^(a[90] & b[116])^(a[89] & b[117])^(a[88] & b[118])^(a[87] & b[119])^(a[86] & b[120])^(a[85] & b[121])^(a[84] & b[122])^(a[83] & b[123])^(a[82] & b[124])^(a[81] & b[125])^(a[80] & b[126])^(a[79] & b[127])^(a[78] & b[128])^(a[77] & b[129])^(a[76] & b[130])^(a[75] & b[131])^(a[74] & b[132])^(a[73] & b[133])^(a[72] & b[134])^(a[71] & b[135])^(a[70] & b[136])^(a[69] & b[137])^(a[68] & b[138])^(a[67] & b[139])^(a[66] & b[140])^(a[65] & b[141])^(a[64] & b[142])^(a[63] & b[143])^(a[62] & b[144])^(a[61] & b[145])^(a[60] & b[146])^(a[59] & b[147])^(a[58] & b[148])^(a[57] & b[149])^(a[56] & b[150])^(a[55] & b[151])^(a[54] & b[152])^(a[53] & b[153])^(a[52] & b[154])^(a[51] & b[155])^(a[50] & b[156])^(a[49] & b[157])^(a[48] & b[158])^(a[47] & b[159])^(a[46] & b[160])^(a[45] & b[161])^(a[44] & b[162])^(a[43] & b[163])^(a[42] & b[164])^(a[41] & b[165])^(a[40] & b[166])^(a[39] & b[167])^(a[38] & b[168])^(a[37] & b[169])^(a[36] & b[170])^(a[35] & b[171])^(a[34] & b[172])^(a[33] & b[173])^(a[32] & b[174])^(a[31] & b[175])^(a[30] & b[176])^(a[29] & b[177])^(a[28] & b[178])^(a[27] & b[179])^(a[26] & b[180])^(a[25] & b[181])^(a[24] & b[182])^(a[23] & b[183])^(a[22] & b[184])^(a[21] & b[185])^(a[20] & b[186])^(a[19] & b[187])^(a[18] & b[188])^(a[17] & b[189])^(a[16] & b[190])^(a[15] & b[191])^(a[14] & b[192])^(a[13] & b[193])^(a[12] & b[194])^(a[11] & b[195])^(a[10] & b[196])^(a[9] & b[197])^(a[8] & b[198])^(a[7] & b[199])^(a[6] & b[200])^(a[5] & b[201])^(a[4] & b[202])^(a[3] & b[203])^(a[2] & b[204])^(a[1] & b[205])^(a[0] & b[206]);
assign y[207] = (a[207] & b[0])^(a[206] & b[1])^(a[205] & b[2])^(a[204] & b[3])^(a[203] & b[4])^(a[202] & b[5])^(a[201] & b[6])^(a[200] & b[7])^(a[199] & b[8])^(a[198] & b[9])^(a[197] & b[10])^(a[196] & b[11])^(a[195] & b[12])^(a[194] & b[13])^(a[193] & b[14])^(a[192] & b[15])^(a[191] & b[16])^(a[190] & b[17])^(a[189] & b[18])^(a[188] & b[19])^(a[187] & b[20])^(a[186] & b[21])^(a[185] & b[22])^(a[184] & b[23])^(a[183] & b[24])^(a[182] & b[25])^(a[181] & b[26])^(a[180] & b[27])^(a[179] & b[28])^(a[178] & b[29])^(a[177] & b[30])^(a[176] & b[31])^(a[175] & b[32])^(a[174] & b[33])^(a[173] & b[34])^(a[172] & b[35])^(a[171] & b[36])^(a[170] & b[37])^(a[169] & b[38])^(a[168] & b[39])^(a[167] & b[40])^(a[166] & b[41])^(a[165] & b[42])^(a[164] & b[43])^(a[163] & b[44])^(a[162] & b[45])^(a[161] & b[46])^(a[160] & b[47])^(a[159] & b[48])^(a[158] & b[49])^(a[157] & b[50])^(a[156] & b[51])^(a[155] & b[52])^(a[154] & b[53])^(a[153] & b[54])^(a[152] & b[55])^(a[151] & b[56])^(a[150] & b[57])^(a[149] & b[58])^(a[148] & b[59])^(a[147] & b[60])^(a[146] & b[61])^(a[145] & b[62])^(a[144] & b[63])^(a[143] & b[64])^(a[142] & b[65])^(a[141] & b[66])^(a[140] & b[67])^(a[139] & b[68])^(a[138] & b[69])^(a[137] & b[70])^(a[136] & b[71])^(a[135] & b[72])^(a[134] & b[73])^(a[133] & b[74])^(a[132] & b[75])^(a[131] & b[76])^(a[130] & b[77])^(a[129] & b[78])^(a[128] & b[79])^(a[127] & b[80])^(a[126] & b[81])^(a[125] & b[82])^(a[124] & b[83])^(a[123] & b[84])^(a[122] & b[85])^(a[121] & b[86])^(a[120] & b[87])^(a[119] & b[88])^(a[118] & b[89])^(a[117] & b[90])^(a[116] & b[91])^(a[115] & b[92])^(a[114] & b[93])^(a[113] & b[94])^(a[112] & b[95])^(a[111] & b[96])^(a[110] & b[97])^(a[109] & b[98])^(a[108] & b[99])^(a[107] & b[100])^(a[106] & b[101])^(a[105] & b[102])^(a[104] & b[103])^(a[103] & b[104])^(a[102] & b[105])^(a[101] & b[106])^(a[100] & b[107])^(a[99] & b[108])^(a[98] & b[109])^(a[97] & b[110])^(a[96] & b[111])^(a[95] & b[112])^(a[94] & b[113])^(a[93] & b[114])^(a[92] & b[115])^(a[91] & b[116])^(a[90] & b[117])^(a[89] & b[118])^(a[88] & b[119])^(a[87] & b[120])^(a[86] & b[121])^(a[85] & b[122])^(a[84] & b[123])^(a[83] & b[124])^(a[82] & b[125])^(a[81] & b[126])^(a[80] & b[127])^(a[79] & b[128])^(a[78] & b[129])^(a[77] & b[130])^(a[76] & b[131])^(a[75] & b[132])^(a[74] & b[133])^(a[73] & b[134])^(a[72] & b[135])^(a[71] & b[136])^(a[70] & b[137])^(a[69] & b[138])^(a[68] & b[139])^(a[67] & b[140])^(a[66] & b[141])^(a[65] & b[142])^(a[64] & b[143])^(a[63] & b[144])^(a[62] & b[145])^(a[61] & b[146])^(a[60] & b[147])^(a[59] & b[148])^(a[58] & b[149])^(a[57] & b[150])^(a[56] & b[151])^(a[55] & b[152])^(a[54] & b[153])^(a[53] & b[154])^(a[52] & b[155])^(a[51] & b[156])^(a[50] & b[157])^(a[49] & b[158])^(a[48] & b[159])^(a[47] & b[160])^(a[46] & b[161])^(a[45] & b[162])^(a[44] & b[163])^(a[43] & b[164])^(a[42] & b[165])^(a[41] & b[166])^(a[40] & b[167])^(a[39] & b[168])^(a[38] & b[169])^(a[37] & b[170])^(a[36] & b[171])^(a[35] & b[172])^(a[34] & b[173])^(a[33] & b[174])^(a[32] & b[175])^(a[31] & b[176])^(a[30] & b[177])^(a[29] & b[178])^(a[28] & b[179])^(a[27] & b[180])^(a[26] & b[181])^(a[25] & b[182])^(a[24] & b[183])^(a[23] & b[184])^(a[22] & b[185])^(a[21] & b[186])^(a[20] & b[187])^(a[19] & b[188])^(a[18] & b[189])^(a[17] & b[190])^(a[16] & b[191])^(a[15] & b[192])^(a[14] & b[193])^(a[13] & b[194])^(a[12] & b[195])^(a[11] & b[196])^(a[10] & b[197])^(a[9] & b[198])^(a[8] & b[199])^(a[7] & b[200])^(a[6] & b[201])^(a[5] & b[202])^(a[4] & b[203])^(a[3] & b[204])^(a[2] & b[205])^(a[1] & b[206])^(a[0] & b[207]);
assign y[208] = (a[208] & b[0])^(a[207] & b[1])^(a[206] & b[2])^(a[205] & b[3])^(a[204] & b[4])^(a[203] & b[5])^(a[202] & b[6])^(a[201] & b[7])^(a[200] & b[8])^(a[199] & b[9])^(a[198] & b[10])^(a[197] & b[11])^(a[196] & b[12])^(a[195] & b[13])^(a[194] & b[14])^(a[193] & b[15])^(a[192] & b[16])^(a[191] & b[17])^(a[190] & b[18])^(a[189] & b[19])^(a[188] & b[20])^(a[187] & b[21])^(a[186] & b[22])^(a[185] & b[23])^(a[184] & b[24])^(a[183] & b[25])^(a[182] & b[26])^(a[181] & b[27])^(a[180] & b[28])^(a[179] & b[29])^(a[178] & b[30])^(a[177] & b[31])^(a[176] & b[32])^(a[175] & b[33])^(a[174] & b[34])^(a[173] & b[35])^(a[172] & b[36])^(a[171] & b[37])^(a[170] & b[38])^(a[169] & b[39])^(a[168] & b[40])^(a[167] & b[41])^(a[166] & b[42])^(a[165] & b[43])^(a[164] & b[44])^(a[163] & b[45])^(a[162] & b[46])^(a[161] & b[47])^(a[160] & b[48])^(a[159] & b[49])^(a[158] & b[50])^(a[157] & b[51])^(a[156] & b[52])^(a[155] & b[53])^(a[154] & b[54])^(a[153] & b[55])^(a[152] & b[56])^(a[151] & b[57])^(a[150] & b[58])^(a[149] & b[59])^(a[148] & b[60])^(a[147] & b[61])^(a[146] & b[62])^(a[145] & b[63])^(a[144] & b[64])^(a[143] & b[65])^(a[142] & b[66])^(a[141] & b[67])^(a[140] & b[68])^(a[139] & b[69])^(a[138] & b[70])^(a[137] & b[71])^(a[136] & b[72])^(a[135] & b[73])^(a[134] & b[74])^(a[133] & b[75])^(a[132] & b[76])^(a[131] & b[77])^(a[130] & b[78])^(a[129] & b[79])^(a[128] & b[80])^(a[127] & b[81])^(a[126] & b[82])^(a[125] & b[83])^(a[124] & b[84])^(a[123] & b[85])^(a[122] & b[86])^(a[121] & b[87])^(a[120] & b[88])^(a[119] & b[89])^(a[118] & b[90])^(a[117] & b[91])^(a[116] & b[92])^(a[115] & b[93])^(a[114] & b[94])^(a[113] & b[95])^(a[112] & b[96])^(a[111] & b[97])^(a[110] & b[98])^(a[109] & b[99])^(a[108] & b[100])^(a[107] & b[101])^(a[106] & b[102])^(a[105] & b[103])^(a[104] & b[104])^(a[103] & b[105])^(a[102] & b[106])^(a[101] & b[107])^(a[100] & b[108])^(a[99] & b[109])^(a[98] & b[110])^(a[97] & b[111])^(a[96] & b[112])^(a[95] & b[113])^(a[94] & b[114])^(a[93] & b[115])^(a[92] & b[116])^(a[91] & b[117])^(a[90] & b[118])^(a[89] & b[119])^(a[88] & b[120])^(a[87] & b[121])^(a[86] & b[122])^(a[85] & b[123])^(a[84] & b[124])^(a[83] & b[125])^(a[82] & b[126])^(a[81] & b[127])^(a[80] & b[128])^(a[79] & b[129])^(a[78] & b[130])^(a[77] & b[131])^(a[76] & b[132])^(a[75] & b[133])^(a[74] & b[134])^(a[73] & b[135])^(a[72] & b[136])^(a[71] & b[137])^(a[70] & b[138])^(a[69] & b[139])^(a[68] & b[140])^(a[67] & b[141])^(a[66] & b[142])^(a[65] & b[143])^(a[64] & b[144])^(a[63] & b[145])^(a[62] & b[146])^(a[61] & b[147])^(a[60] & b[148])^(a[59] & b[149])^(a[58] & b[150])^(a[57] & b[151])^(a[56] & b[152])^(a[55] & b[153])^(a[54] & b[154])^(a[53] & b[155])^(a[52] & b[156])^(a[51] & b[157])^(a[50] & b[158])^(a[49] & b[159])^(a[48] & b[160])^(a[47] & b[161])^(a[46] & b[162])^(a[45] & b[163])^(a[44] & b[164])^(a[43] & b[165])^(a[42] & b[166])^(a[41] & b[167])^(a[40] & b[168])^(a[39] & b[169])^(a[38] & b[170])^(a[37] & b[171])^(a[36] & b[172])^(a[35] & b[173])^(a[34] & b[174])^(a[33] & b[175])^(a[32] & b[176])^(a[31] & b[177])^(a[30] & b[178])^(a[29] & b[179])^(a[28] & b[180])^(a[27] & b[181])^(a[26] & b[182])^(a[25] & b[183])^(a[24] & b[184])^(a[23] & b[185])^(a[22] & b[186])^(a[21] & b[187])^(a[20] & b[188])^(a[19] & b[189])^(a[18] & b[190])^(a[17] & b[191])^(a[16] & b[192])^(a[15] & b[193])^(a[14] & b[194])^(a[13] & b[195])^(a[12] & b[196])^(a[11] & b[197])^(a[10] & b[198])^(a[9] & b[199])^(a[8] & b[200])^(a[7] & b[201])^(a[6] & b[202])^(a[5] & b[203])^(a[4] & b[204])^(a[3] & b[205])^(a[2] & b[206])^(a[1] & b[207])^(a[0] & b[208]);
assign y[209] = (a[209] & b[0])^(a[208] & b[1])^(a[207] & b[2])^(a[206] & b[3])^(a[205] & b[4])^(a[204] & b[5])^(a[203] & b[6])^(a[202] & b[7])^(a[201] & b[8])^(a[200] & b[9])^(a[199] & b[10])^(a[198] & b[11])^(a[197] & b[12])^(a[196] & b[13])^(a[195] & b[14])^(a[194] & b[15])^(a[193] & b[16])^(a[192] & b[17])^(a[191] & b[18])^(a[190] & b[19])^(a[189] & b[20])^(a[188] & b[21])^(a[187] & b[22])^(a[186] & b[23])^(a[185] & b[24])^(a[184] & b[25])^(a[183] & b[26])^(a[182] & b[27])^(a[181] & b[28])^(a[180] & b[29])^(a[179] & b[30])^(a[178] & b[31])^(a[177] & b[32])^(a[176] & b[33])^(a[175] & b[34])^(a[174] & b[35])^(a[173] & b[36])^(a[172] & b[37])^(a[171] & b[38])^(a[170] & b[39])^(a[169] & b[40])^(a[168] & b[41])^(a[167] & b[42])^(a[166] & b[43])^(a[165] & b[44])^(a[164] & b[45])^(a[163] & b[46])^(a[162] & b[47])^(a[161] & b[48])^(a[160] & b[49])^(a[159] & b[50])^(a[158] & b[51])^(a[157] & b[52])^(a[156] & b[53])^(a[155] & b[54])^(a[154] & b[55])^(a[153] & b[56])^(a[152] & b[57])^(a[151] & b[58])^(a[150] & b[59])^(a[149] & b[60])^(a[148] & b[61])^(a[147] & b[62])^(a[146] & b[63])^(a[145] & b[64])^(a[144] & b[65])^(a[143] & b[66])^(a[142] & b[67])^(a[141] & b[68])^(a[140] & b[69])^(a[139] & b[70])^(a[138] & b[71])^(a[137] & b[72])^(a[136] & b[73])^(a[135] & b[74])^(a[134] & b[75])^(a[133] & b[76])^(a[132] & b[77])^(a[131] & b[78])^(a[130] & b[79])^(a[129] & b[80])^(a[128] & b[81])^(a[127] & b[82])^(a[126] & b[83])^(a[125] & b[84])^(a[124] & b[85])^(a[123] & b[86])^(a[122] & b[87])^(a[121] & b[88])^(a[120] & b[89])^(a[119] & b[90])^(a[118] & b[91])^(a[117] & b[92])^(a[116] & b[93])^(a[115] & b[94])^(a[114] & b[95])^(a[113] & b[96])^(a[112] & b[97])^(a[111] & b[98])^(a[110] & b[99])^(a[109] & b[100])^(a[108] & b[101])^(a[107] & b[102])^(a[106] & b[103])^(a[105] & b[104])^(a[104] & b[105])^(a[103] & b[106])^(a[102] & b[107])^(a[101] & b[108])^(a[100] & b[109])^(a[99] & b[110])^(a[98] & b[111])^(a[97] & b[112])^(a[96] & b[113])^(a[95] & b[114])^(a[94] & b[115])^(a[93] & b[116])^(a[92] & b[117])^(a[91] & b[118])^(a[90] & b[119])^(a[89] & b[120])^(a[88] & b[121])^(a[87] & b[122])^(a[86] & b[123])^(a[85] & b[124])^(a[84] & b[125])^(a[83] & b[126])^(a[82] & b[127])^(a[81] & b[128])^(a[80] & b[129])^(a[79] & b[130])^(a[78] & b[131])^(a[77] & b[132])^(a[76] & b[133])^(a[75] & b[134])^(a[74] & b[135])^(a[73] & b[136])^(a[72] & b[137])^(a[71] & b[138])^(a[70] & b[139])^(a[69] & b[140])^(a[68] & b[141])^(a[67] & b[142])^(a[66] & b[143])^(a[65] & b[144])^(a[64] & b[145])^(a[63] & b[146])^(a[62] & b[147])^(a[61] & b[148])^(a[60] & b[149])^(a[59] & b[150])^(a[58] & b[151])^(a[57] & b[152])^(a[56] & b[153])^(a[55] & b[154])^(a[54] & b[155])^(a[53] & b[156])^(a[52] & b[157])^(a[51] & b[158])^(a[50] & b[159])^(a[49] & b[160])^(a[48] & b[161])^(a[47] & b[162])^(a[46] & b[163])^(a[45] & b[164])^(a[44] & b[165])^(a[43] & b[166])^(a[42] & b[167])^(a[41] & b[168])^(a[40] & b[169])^(a[39] & b[170])^(a[38] & b[171])^(a[37] & b[172])^(a[36] & b[173])^(a[35] & b[174])^(a[34] & b[175])^(a[33] & b[176])^(a[32] & b[177])^(a[31] & b[178])^(a[30] & b[179])^(a[29] & b[180])^(a[28] & b[181])^(a[27] & b[182])^(a[26] & b[183])^(a[25] & b[184])^(a[24] & b[185])^(a[23] & b[186])^(a[22] & b[187])^(a[21] & b[188])^(a[20] & b[189])^(a[19] & b[190])^(a[18] & b[191])^(a[17] & b[192])^(a[16] & b[193])^(a[15] & b[194])^(a[14] & b[195])^(a[13] & b[196])^(a[12] & b[197])^(a[11] & b[198])^(a[10] & b[199])^(a[9] & b[200])^(a[8] & b[201])^(a[7] & b[202])^(a[6] & b[203])^(a[5] & b[204])^(a[4] & b[205])^(a[3] & b[206])^(a[2] & b[207])^(a[1] & b[208])^(a[0] & b[209]);
assign y[210] = (a[210] & b[0])^(a[209] & b[1])^(a[208] & b[2])^(a[207] & b[3])^(a[206] & b[4])^(a[205] & b[5])^(a[204] & b[6])^(a[203] & b[7])^(a[202] & b[8])^(a[201] & b[9])^(a[200] & b[10])^(a[199] & b[11])^(a[198] & b[12])^(a[197] & b[13])^(a[196] & b[14])^(a[195] & b[15])^(a[194] & b[16])^(a[193] & b[17])^(a[192] & b[18])^(a[191] & b[19])^(a[190] & b[20])^(a[189] & b[21])^(a[188] & b[22])^(a[187] & b[23])^(a[186] & b[24])^(a[185] & b[25])^(a[184] & b[26])^(a[183] & b[27])^(a[182] & b[28])^(a[181] & b[29])^(a[180] & b[30])^(a[179] & b[31])^(a[178] & b[32])^(a[177] & b[33])^(a[176] & b[34])^(a[175] & b[35])^(a[174] & b[36])^(a[173] & b[37])^(a[172] & b[38])^(a[171] & b[39])^(a[170] & b[40])^(a[169] & b[41])^(a[168] & b[42])^(a[167] & b[43])^(a[166] & b[44])^(a[165] & b[45])^(a[164] & b[46])^(a[163] & b[47])^(a[162] & b[48])^(a[161] & b[49])^(a[160] & b[50])^(a[159] & b[51])^(a[158] & b[52])^(a[157] & b[53])^(a[156] & b[54])^(a[155] & b[55])^(a[154] & b[56])^(a[153] & b[57])^(a[152] & b[58])^(a[151] & b[59])^(a[150] & b[60])^(a[149] & b[61])^(a[148] & b[62])^(a[147] & b[63])^(a[146] & b[64])^(a[145] & b[65])^(a[144] & b[66])^(a[143] & b[67])^(a[142] & b[68])^(a[141] & b[69])^(a[140] & b[70])^(a[139] & b[71])^(a[138] & b[72])^(a[137] & b[73])^(a[136] & b[74])^(a[135] & b[75])^(a[134] & b[76])^(a[133] & b[77])^(a[132] & b[78])^(a[131] & b[79])^(a[130] & b[80])^(a[129] & b[81])^(a[128] & b[82])^(a[127] & b[83])^(a[126] & b[84])^(a[125] & b[85])^(a[124] & b[86])^(a[123] & b[87])^(a[122] & b[88])^(a[121] & b[89])^(a[120] & b[90])^(a[119] & b[91])^(a[118] & b[92])^(a[117] & b[93])^(a[116] & b[94])^(a[115] & b[95])^(a[114] & b[96])^(a[113] & b[97])^(a[112] & b[98])^(a[111] & b[99])^(a[110] & b[100])^(a[109] & b[101])^(a[108] & b[102])^(a[107] & b[103])^(a[106] & b[104])^(a[105] & b[105])^(a[104] & b[106])^(a[103] & b[107])^(a[102] & b[108])^(a[101] & b[109])^(a[100] & b[110])^(a[99] & b[111])^(a[98] & b[112])^(a[97] & b[113])^(a[96] & b[114])^(a[95] & b[115])^(a[94] & b[116])^(a[93] & b[117])^(a[92] & b[118])^(a[91] & b[119])^(a[90] & b[120])^(a[89] & b[121])^(a[88] & b[122])^(a[87] & b[123])^(a[86] & b[124])^(a[85] & b[125])^(a[84] & b[126])^(a[83] & b[127])^(a[82] & b[128])^(a[81] & b[129])^(a[80] & b[130])^(a[79] & b[131])^(a[78] & b[132])^(a[77] & b[133])^(a[76] & b[134])^(a[75] & b[135])^(a[74] & b[136])^(a[73] & b[137])^(a[72] & b[138])^(a[71] & b[139])^(a[70] & b[140])^(a[69] & b[141])^(a[68] & b[142])^(a[67] & b[143])^(a[66] & b[144])^(a[65] & b[145])^(a[64] & b[146])^(a[63] & b[147])^(a[62] & b[148])^(a[61] & b[149])^(a[60] & b[150])^(a[59] & b[151])^(a[58] & b[152])^(a[57] & b[153])^(a[56] & b[154])^(a[55] & b[155])^(a[54] & b[156])^(a[53] & b[157])^(a[52] & b[158])^(a[51] & b[159])^(a[50] & b[160])^(a[49] & b[161])^(a[48] & b[162])^(a[47] & b[163])^(a[46] & b[164])^(a[45] & b[165])^(a[44] & b[166])^(a[43] & b[167])^(a[42] & b[168])^(a[41] & b[169])^(a[40] & b[170])^(a[39] & b[171])^(a[38] & b[172])^(a[37] & b[173])^(a[36] & b[174])^(a[35] & b[175])^(a[34] & b[176])^(a[33] & b[177])^(a[32] & b[178])^(a[31] & b[179])^(a[30] & b[180])^(a[29] & b[181])^(a[28] & b[182])^(a[27] & b[183])^(a[26] & b[184])^(a[25] & b[185])^(a[24] & b[186])^(a[23] & b[187])^(a[22] & b[188])^(a[21] & b[189])^(a[20] & b[190])^(a[19] & b[191])^(a[18] & b[192])^(a[17] & b[193])^(a[16] & b[194])^(a[15] & b[195])^(a[14] & b[196])^(a[13] & b[197])^(a[12] & b[198])^(a[11] & b[199])^(a[10] & b[200])^(a[9] & b[201])^(a[8] & b[202])^(a[7] & b[203])^(a[6] & b[204])^(a[5] & b[205])^(a[4] & b[206])^(a[3] & b[207])^(a[2] & b[208])^(a[1] & b[209])^(a[0] & b[210]);
assign y[211] = (a[211] & b[0])^(a[210] & b[1])^(a[209] & b[2])^(a[208] & b[3])^(a[207] & b[4])^(a[206] & b[5])^(a[205] & b[6])^(a[204] & b[7])^(a[203] & b[8])^(a[202] & b[9])^(a[201] & b[10])^(a[200] & b[11])^(a[199] & b[12])^(a[198] & b[13])^(a[197] & b[14])^(a[196] & b[15])^(a[195] & b[16])^(a[194] & b[17])^(a[193] & b[18])^(a[192] & b[19])^(a[191] & b[20])^(a[190] & b[21])^(a[189] & b[22])^(a[188] & b[23])^(a[187] & b[24])^(a[186] & b[25])^(a[185] & b[26])^(a[184] & b[27])^(a[183] & b[28])^(a[182] & b[29])^(a[181] & b[30])^(a[180] & b[31])^(a[179] & b[32])^(a[178] & b[33])^(a[177] & b[34])^(a[176] & b[35])^(a[175] & b[36])^(a[174] & b[37])^(a[173] & b[38])^(a[172] & b[39])^(a[171] & b[40])^(a[170] & b[41])^(a[169] & b[42])^(a[168] & b[43])^(a[167] & b[44])^(a[166] & b[45])^(a[165] & b[46])^(a[164] & b[47])^(a[163] & b[48])^(a[162] & b[49])^(a[161] & b[50])^(a[160] & b[51])^(a[159] & b[52])^(a[158] & b[53])^(a[157] & b[54])^(a[156] & b[55])^(a[155] & b[56])^(a[154] & b[57])^(a[153] & b[58])^(a[152] & b[59])^(a[151] & b[60])^(a[150] & b[61])^(a[149] & b[62])^(a[148] & b[63])^(a[147] & b[64])^(a[146] & b[65])^(a[145] & b[66])^(a[144] & b[67])^(a[143] & b[68])^(a[142] & b[69])^(a[141] & b[70])^(a[140] & b[71])^(a[139] & b[72])^(a[138] & b[73])^(a[137] & b[74])^(a[136] & b[75])^(a[135] & b[76])^(a[134] & b[77])^(a[133] & b[78])^(a[132] & b[79])^(a[131] & b[80])^(a[130] & b[81])^(a[129] & b[82])^(a[128] & b[83])^(a[127] & b[84])^(a[126] & b[85])^(a[125] & b[86])^(a[124] & b[87])^(a[123] & b[88])^(a[122] & b[89])^(a[121] & b[90])^(a[120] & b[91])^(a[119] & b[92])^(a[118] & b[93])^(a[117] & b[94])^(a[116] & b[95])^(a[115] & b[96])^(a[114] & b[97])^(a[113] & b[98])^(a[112] & b[99])^(a[111] & b[100])^(a[110] & b[101])^(a[109] & b[102])^(a[108] & b[103])^(a[107] & b[104])^(a[106] & b[105])^(a[105] & b[106])^(a[104] & b[107])^(a[103] & b[108])^(a[102] & b[109])^(a[101] & b[110])^(a[100] & b[111])^(a[99] & b[112])^(a[98] & b[113])^(a[97] & b[114])^(a[96] & b[115])^(a[95] & b[116])^(a[94] & b[117])^(a[93] & b[118])^(a[92] & b[119])^(a[91] & b[120])^(a[90] & b[121])^(a[89] & b[122])^(a[88] & b[123])^(a[87] & b[124])^(a[86] & b[125])^(a[85] & b[126])^(a[84] & b[127])^(a[83] & b[128])^(a[82] & b[129])^(a[81] & b[130])^(a[80] & b[131])^(a[79] & b[132])^(a[78] & b[133])^(a[77] & b[134])^(a[76] & b[135])^(a[75] & b[136])^(a[74] & b[137])^(a[73] & b[138])^(a[72] & b[139])^(a[71] & b[140])^(a[70] & b[141])^(a[69] & b[142])^(a[68] & b[143])^(a[67] & b[144])^(a[66] & b[145])^(a[65] & b[146])^(a[64] & b[147])^(a[63] & b[148])^(a[62] & b[149])^(a[61] & b[150])^(a[60] & b[151])^(a[59] & b[152])^(a[58] & b[153])^(a[57] & b[154])^(a[56] & b[155])^(a[55] & b[156])^(a[54] & b[157])^(a[53] & b[158])^(a[52] & b[159])^(a[51] & b[160])^(a[50] & b[161])^(a[49] & b[162])^(a[48] & b[163])^(a[47] & b[164])^(a[46] & b[165])^(a[45] & b[166])^(a[44] & b[167])^(a[43] & b[168])^(a[42] & b[169])^(a[41] & b[170])^(a[40] & b[171])^(a[39] & b[172])^(a[38] & b[173])^(a[37] & b[174])^(a[36] & b[175])^(a[35] & b[176])^(a[34] & b[177])^(a[33] & b[178])^(a[32] & b[179])^(a[31] & b[180])^(a[30] & b[181])^(a[29] & b[182])^(a[28] & b[183])^(a[27] & b[184])^(a[26] & b[185])^(a[25] & b[186])^(a[24] & b[187])^(a[23] & b[188])^(a[22] & b[189])^(a[21] & b[190])^(a[20] & b[191])^(a[19] & b[192])^(a[18] & b[193])^(a[17] & b[194])^(a[16] & b[195])^(a[15] & b[196])^(a[14] & b[197])^(a[13] & b[198])^(a[12] & b[199])^(a[11] & b[200])^(a[10] & b[201])^(a[9] & b[202])^(a[8] & b[203])^(a[7] & b[204])^(a[6] & b[205])^(a[5] & b[206])^(a[4] & b[207])^(a[3] & b[208])^(a[2] & b[209])^(a[1] & b[210])^(a[0] & b[211]);
assign y[212] = (a[212] & b[0])^(a[211] & b[1])^(a[210] & b[2])^(a[209] & b[3])^(a[208] & b[4])^(a[207] & b[5])^(a[206] & b[6])^(a[205] & b[7])^(a[204] & b[8])^(a[203] & b[9])^(a[202] & b[10])^(a[201] & b[11])^(a[200] & b[12])^(a[199] & b[13])^(a[198] & b[14])^(a[197] & b[15])^(a[196] & b[16])^(a[195] & b[17])^(a[194] & b[18])^(a[193] & b[19])^(a[192] & b[20])^(a[191] & b[21])^(a[190] & b[22])^(a[189] & b[23])^(a[188] & b[24])^(a[187] & b[25])^(a[186] & b[26])^(a[185] & b[27])^(a[184] & b[28])^(a[183] & b[29])^(a[182] & b[30])^(a[181] & b[31])^(a[180] & b[32])^(a[179] & b[33])^(a[178] & b[34])^(a[177] & b[35])^(a[176] & b[36])^(a[175] & b[37])^(a[174] & b[38])^(a[173] & b[39])^(a[172] & b[40])^(a[171] & b[41])^(a[170] & b[42])^(a[169] & b[43])^(a[168] & b[44])^(a[167] & b[45])^(a[166] & b[46])^(a[165] & b[47])^(a[164] & b[48])^(a[163] & b[49])^(a[162] & b[50])^(a[161] & b[51])^(a[160] & b[52])^(a[159] & b[53])^(a[158] & b[54])^(a[157] & b[55])^(a[156] & b[56])^(a[155] & b[57])^(a[154] & b[58])^(a[153] & b[59])^(a[152] & b[60])^(a[151] & b[61])^(a[150] & b[62])^(a[149] & b[63])^(a[148] & b[64])^(a[147] & b[65])^(a[146] & b[66])^(a[145] & b[67])^(a[144] & b[68])^(a[143] & b[69])^(a[142] & b[70])^(a[141] & b[71])^(a[140] & b[72])^(a[139] & b[73])^(a[138] & b[74])^(a[137] & b[75])^(a[136] & b[76])^(a[135] & b[77])^(a[134] & b[78])^(a[133] & b[79])^(a[132] & b[80])^(a[131] & b[81])^(a[130] & b[82])^(a[129] & b[83])^(a[128] & b[84])^(a[127] & b[85])^(a[126] & b[86])^(a[125] & b[87])^(a[124] & b[88])^(a[123] & b[89])^(a[122] & b[90])^(a[121] & b[91])^(a[120] & b[92])^(a[119] & b[93])^(a[118] & b[94])^(a[117] & b[95])^(a[116] & b[96])^(a[115] & b[97])^(a[114] & b[98])^(a[113] & b[99])^(a[112] & b[100])^(a[111] & b[101])^(a[110] & b[102])^(a[109] & b[103])^(a[108] & b[104])^(a[107] & b[105])^(a[106] & b[106])^(a[105] & b[107])^(a[104] & b[108])^(a[103] & b[109])^(a[102] & b[110])^(a[101] & b[111])^(a[100] & b[112])^(a[99] & b[113])^(a[98] & b[114])^(a[97] & b[115])^(a[96] & b[116])^(a[95] & b[117])^(a[94] & b[118])^(a[93] & b[119])^(a[92] & b[120])^(a[91] & b[121])^(a[90] & b[122])^(a[89] & b[123])^(a[88] & b[124])^(a[87] & b[125])^(a[86] & b[126])^(a[85] & b[127])^(a[84] & b[128])^(a[83] & b[129])^(a[82] & b[130])^(a[81] & b[131])^(a[80] & b[132])^(a[79] & b[133])^(a[78] & b[134])^(a[77] & b[135])^(a[76] & b[136])^(a[75] & b[137])^(a[74] & b[138])^(a[73] & b[139])^(a[72] & b[140])^(a[71] & b[141])^(a[70] & b[142])^(a[69] & b[143])^(a[68] & b[144])^(a[67] & b[145])^(a[66] & b[146])^(a[65] & b[147])^(a[64] & b[148])^(a[63] & b[149])^(a[62] & b[150])^(a[61] & b[151])^(a[60] & b[152])^(a[59] & b[153])^(a[58] & b[154])^(a[57] & b[155])^(a[56] & b[156])^(a[55] & b[157])^(a[54] & b[158])^(a[53] & b[159])^(a[52] & b[160])^(a[51] & b[161])^(a[50] & b[162])^(a[49] & b[163])^(a[48] & b[164])^(a[47] & b[165])^(a[46] & b[166])^(a[45] & b[167])^(a[44] & b[168])^(a[43] & b[169])^(a[42] & b[170])^(a[41] & b[171])^(a[40] & b[172])^(a[39] & b[173])^(a[38] & b[174])^(a[37] & b[175])^(a[36] & b[176])^(a[35] & b[177])^(a[34] & b[178])^(a[33] & b[179])^(a[32] & b[180])^(a[31] & b[181])^(a[30] & b[182])^(a[29] & b[183])^(a[28] & b[184])^(a[27] & b[185])^(a[26] & b[186])^(a[25] & b[187])^(a[24] & b[188])^(a[23] & b[189])^(a[22] & b[190])^(a[21] & b[191])^(a[20] & b[192])^(a[19] & b[193])^(a[18] & b[194])^(a[17] & b[195])^(a[16] & b[196])^(a[15] & b[197])^(a[14] & b[198])^(a[13] & b[199])^(a[12] & b[200])^(a[11] & b[201])^(a[10] & b[202])^(a[9] & b[203])^(a[8] & b[204])^(a[7] & b[205])^(a[6] & b[206])^(a[5] & b[207])^(a[4] & b[208])^(a[3] & b[209])^(a[2] & b[210])^(a[1] & b[211])^(a[0] & b[212]);
assign y[213] = (a[213] & b[0])^(a[212] & b[1])^(a[211] & b[2])^(a[210] & b[3])^(a[209] & b[4])^(a[208] & b[5])^(a[207] & b[6])^(a[206] & b[7])^(a[205] & b[8])^(a[204] & b[9])^(a[203] & b[10])^(a[202] & b[11])^(a[201] & b[12])^(a[200] & b[13])^(a[199] & b[14])^(a[198] & b[15])^(a[197] & b[16])^(a[196] & b[17])^(a[195] & b[18])^(a[194] & b[19])^(a[193] & b[20])^(a[192] & b[21])^(a[191] & b[22])^(a[190] & b[23])^(a[189] & b[24])^(a[188] & b[25])^(a[187] & b[26])^(a[186] & b[27])^(a[185] & b[28])^(a[184] & b[29])^(a[183] & b[30])^(a[182] & b[31])^(a[181] & b[32])^(a[180] & b[33])^(a[179] & b[34])^(a[178] & b[35])^(a[177] & b[36])^(a[176] & b[37])^(a[175] & b[38])^(a[174] & b[39])^(a[173] & b[40])^(a[172] & b[41])^(a[171] & b[42])^(a[170] & b[43])^(a[169] & b[44])^(a[168] & b[45])^(a[167] & b[46])^(a[166] & b[47])^(a[165] & b[48])^(a[164] & b[49])^(a[163] & b[50])^(a[162] & b[51])^(a[161] & b[52])^(a[160] & b[53])^(a[159] & b[54])^(a[158] & b[55])^(a[157] & b[56])^(a[156] & b[57])^(a[155] & b[58])^(a[154] & b[59])^(a[153] & b[60])^(a[152] & b[61])^(a[151] & b[62])^(a[150] & b[63])^(a[149] & b[64])^(a[148] & b[65])^(a[147] & b[66])^(a[146] & b[67])^(a[145] & b[68])^(a[144] & b[69])^(a[143] & b[70])^(a[142] & b[71])^(a[141] & b[72])^(a[140] & b[73])^(a[139] & b[74])^(a[138] & b[75])^(a[137] & b[76])^(a[136] & b[77])^(a[135] & b[78])^(a[134] & b[79])^(a[133] & b[80])^(a[132] & b[81])^(a[131] & b[82])^(a[130] & b[83])^(a[129] & b[84])^(a[128] & b[85])^(a[127] & b[86])^(a[126] & b[87])^(a[125] & b[88])^(a[124] & b[89])^(a[123] & b[90])^(a[122] & b[91])^(a[121] & b[92])^(a[120] & b[93])^(a[119] & b[94])^(a[118] & b[95])^(a[117] & b[96])^(a[116] & b[97])^(a[115] & b[98])^(a[114] & b[99])^(a[113] & b[100])^(a[112] & b[101])^(a[111] & b[102])^(a[110] & b[103])^(a[109] & b[104])^(a[108] & b[105])^(a[107] & b[106])^(a[106] & b[107])^(a[105] & b[108])^(a[104] & b[109])^(a[103] & b[110])^(a[102] & b[111])^(a[101] & b[112])^(a[100] & b[113])^(a[99] & b[114])^(a[98] & b[115])^(a[97] & b[116])^(a[96] & b[117])^(a[95] & b[118])^(a[94] & b[119])^(a[93] & b[120])^(a[92] & b[121])^(a[91] & b[122])^(a[90] & b[123])^(a[89] & b[124])^(a[88] & b[125])^(a[87] & b[126])^(a[86] & b[127])^(a[85] & b[128])^(a[84] & b[129])^(a[83] & b[130])^(a[82] & b[131])^(a[81] & b[132])^(a[80] & b[133])^(a[79] & b[134])^(a[78] & b[135])^(a[77] & b[136])^(a[76] & b[137])^(a[75] & b[138])^(a[74] & b[139])^(a[73] & b[140])^(a[72] & b[141])^(a[71] & b[142])^(a[70] & b[143])^(a[69] & b[144])^(a[68] & b[145])^(a[67] & b[146])^(a[66] & b[147])^(a[65] & b[148])^(a[64] & b[149])^(a[63] & b[150])^(a[62] & b[151])^(a[61] & b[152])^(a[60] & b[153])^(a[59] & b[154])^(a[58] & b[155])^(a[57] & b[156])^(a[56] & b[157])^(a[55] & b[158])^(a[54] & b[159])^(a[53] & b[160])^(a[52] & b[161])^(a[51] & b[162])^(a[50] & b[163])^(a[49] & b[164])^(a[48] & b[165])^(a[47] & b[166])^(a[46] & b[167])^(a[45] & b[168])^(a[44] & b[169])^(a[43] & b[170])^(a[42] & b[171])^(a[41] & b[172])^(a[40] & b[173])^(a[39] & b[174])^(a[38] & b[175])^(a[37] & b[176])^(a[36] & b[177])^(a[35] & b[178])^(a[34] & b[179])^(a[33] & b[180])^(a[32] & b[181])^(a[31] & b[182])^(a[30] & b[183])^(a[29] & b[184])^(a[28] & b[185])^(a[27] & b[186])^(a[26] & b[187])^(a[25] & b[188])^(a[24] & b[189])^(a[23] & b[190])^(a[22] & b[191])^(a[21] & b[192])^(a[20] & b[193])^(a[19] & b[194])^(a[18] & b[195])^(a[17] & b[196])^(a[16] & b[197])^(a[15] & b[198])^(a[14] & b[199])^(a[13] & b[200])^(a[12] & b[201])^(a[11] & b[202])^(a[10] & b[203])^(a[9] & b[204])^(a[8] & b[205])^(a[7] & b[206])^(a[6] & b[207])^(a[5] & b[208])^(a[4] & b[209])^(a[3] & b[210])^(a[2] & b[211])^(a[1] & b[212])^(a[0] & b[213]);
assign y[214] = (a[214] & b[0])^(a[213] & b[1])^(a[212] & b[2])^(a[211] & b[3])^(a[210] & b[4])^(a[209] & b[5])^(a[208] & b[6])^(a[207] & b[7])^(a[206] & b[8])^(a[205] & b[9])^(a[204] & b[10])^(a[203] & b[11])^(a[202] & b[12])^(a[201] & b[13])^(a[200] & b[14])^(a[199] & b[15])^(a[198] & b[16])^(a[197] & b[17])^(a[196] & b[18])^(a[195] & b[19])^(a[194] & b[20])^(a[193] & b[21])^(a[192] & b[22])^(a[191] & b[23])^(a[190] & b[24])^(a[189] & b[25])^(a[188] & b[26])^(a[187] & b[27])^(a[186] & b[28])^(a[185] & b[29])^(a[184] & b[30])^(a[183] & b[31])^(a[182] & b[32])^(a[181] & b[33])^(a[180] & b[34])^(a[179] & b[35])^(a[178] & b[36])^(a[177] & b[37])^(a[176] & b[38])^(a[175] & b[39])^(a[174] & b[40])^(a[173] & b[41])^(a[172] & b[42])^(a[171] & b[43])^(a[170] & b[44])^(a[169] & b[45])^(a[168] & b[46])^(a[167] & b[47])^(a[166] & b[48])^(a[165] & b[49])^(a[164] & b[50])^(a[163] & b[51])^(a[162] & b[52])^(a[161] & b[53])^(a[160] & b[54])^(a[159] & b[55])^(a[158] & b[56])^(a[157] & b[57])^(a[156] & b[58])^(a[155] & b[59])^(a[154] & b[60])^(a[153] & b[61])^(a[152] & b[62])^(a[151] & b[63])^(a[150] & b[64])^(a[149] & b[65])^(a[148] & b[66])^(a[147] & b[67])^(a[146] & b[68])^(a[145] & b[69])^(a[144] & b[70])^(a[143] & b[71])^(a[142] & b[72])^(a[141] & b[73])^(a[140] & b[74])^(a[139] & b[75])^(a[138] & b[76])^(a[137] & b[77])^(a[136] & b[78])^(a[135] & b[79])^(a[134] & b[80])^(a[133] & b[81])^(a[132] & b[82])^(a[131] & b[83])^(a[130] & b[84])^(a[129] & b[85])^(a[128] & b[86])^(a[127] & b[87])^(a[126] & b[88])^(a[125] & b[89])^(a[124] & b[90])^(a[123] & b[91])^(a[122] & b[92])^(a[121] & b[93])^(a[120] & b[94])^(a[119] & b[95])^(a[118] & b[96])^(a[117] & b[97])^(a[116] & b[98])^(a[115] & b[99])^(a[114] & b[100])^(a[113] & b[101])^(a[112] & b[102])^(a[111] & b[103])^(a[110] & b[104])^(a[109] & b[105])^(a[108] & b[106])^(a[107] & b[107])^(a[106] & b[108])^(a[105] & b[109])^(a[104] & b[110])^(a[103] & b[111])^(a[102] & b[112])^(a[101] & b[113])^(a[100] & b[114])^(a[99] & b[115])^(a[98] & b[116])^(a[97] & b[117])^(a[96] & b[118])^(a[95] & b[119])^(a[94] & b[120])^(a[93] & b[121])^(a[92] & b[122])^(a[91] & b[123])^(a[90] & b[124])^(a[89] & b[125])^(a[88] & b[126])^(a[87] & b[127])^(a[86] & b[128])^(a[85] & b[129])^(a[84] & b[130])^(a[83] & b[131])^(a[82] & b[132])^(a[81] & b[133])^(a[80] & b[134])^(a[79] & b[135])^(a[78] & b[136])^(a[77] & b[137])^(a[76] & b[138])^(a[75] & b[139])^(a[74] & b[140])^(a[73] & b[141])^(a[72] & b[142])^(a[71] & b[143])^(a[70] & b[144])^(a[69] & b[145])^(a[68] & b[146])^(a[67] & b[147])^(a[66] & b[148])^(a[65] & b[149])^(a[64] & b[150])^(a[63] & b[151])^(a[62] & b[152])^(a[61] & b[153])^(a[60] & b[154])^(a[59] & b[155])^(a[58] & b[156])^(a[57] & b[157])^(a[56] & b[158])^(a[55] & b[159])^(a[54] & b[160])^(a[53] & b[161])^(a[52] & b[162])^(a[51] & b[163])^(a[50] & b[164])^(a[49] & b[165])^(a[48] & b[166])^(a[47] & b[167])^(a[46] & b[168])^(a[45] & b[169])^(a[44] & b[170])^(a[43] & b[171])^(a[42] & b[172])^(a[41] & b[173])^(a[40] & b[174])^(a[39] & b[175])^(a[38] & b[176])^(a[37] & b[177])^(a[36] & b[178])^(a[35] & b[179])^(a[34] & b[180])^(a[33] & b[181])^(a[32] & b[182])^(a[31] & b[183])^(a[30] & b[184])^(a[29] & b[185])^(a[28] & b[186])^(a[27] & b[187])^(a[26] & b[188])^(a[25] & b[189])^(a[24] & b[190])^(a[23] & b[191])^(a[22] & b[192])^(a[21] & b[193])^(a[20] & b[194])^(a[19] & b[195])^(a[18] & b[196])^(a[17] & b[197])^(a[16] & b[198])^(a[15] & b[199])^(a[14] & b[200])^(a[13] & b[201])^(a[12] & b[202])^(a[11] & b[203])^(a[10] & b[204])^(a[9] & b[205])^(a[8] & b[206])^(a[7] & b[207])^(a[6] & b[208])^(a[5] & b[209])^(a[4] & b[210])^(a[3] & b[211])^(a[2] & b[212])^(a[1] & b[213])^(a[0] & b[214]);
assign y[215] = (a[215] & b[0])^(a[214] & b[1])^(a[213] & b[2])^(a[212] & b[3])^(a[211] & b[4])^(a[210] & b[5])^(a[209] & b[6])^(a[208] & b[7])^(a[207] & b[8])^(a[206] & b[9])^(a[205] & b[10])^(a[204] & b[11])^(a[203] & b[12])^(a[202] & b[13])^(a[201] & b[14])^(a[200] & b[15])^(a[199] & b[16])^(a[198] & b[17])^(a[197] & b[18])^(a[196] & b[19])^(a[195] & b[20])^(a[194] & b[21])^(a[193] & b[22])^(a[192] & b[23])^(a[191] & b[24])^(a[190] & b[25])^(a[189] & b[26])^(a[188] & b[27])^(a[187] & b[28])^(a[186] & b[29])^(a[185] & b[30])^(a[184] & b[31])^(a[183] & b[32])^(a[182] & b[33])^(a[181] & b[34])^(a[180] & b[35])^(a[179] & b[36])^(a[178] & b[37])^(a[177] & b[38])^(a[176] & b[39])^(a[175] & b[40])^(a[174] & b[41])^(a[173] & b[42])^(a[172] & b[43])^(a[171] & b[44])^(a[170] & b[45])^(a[169] & b[46])^(a[168] & b[47])^(a[167] & b[48])^(a[166] & b[49])^(a[165] & b[50])^(a[164] & b[51])^(a[163] & b[52])^(a[162] & b[53])^(a[161] & b[54])^(a[160] & b[55])^(a[159] & b[56])^(a[158] & b[57])^(a[157] & b[58])^(a[156] & b[59])^(a[155] & b[60])^(a[154] & b[61])^(a[153] & b[62])^(a[152] & b[63])^(a[151] & b[64])^(a[150] & b[65])^(a[149] & b[66])^(a[148] & b[67])^(a[147] & b[68])^(a[146] & b[69])^(a[145] & b[70])^(a[144] & b[71])^(a[143] & b[72])^(a[142] & b[73])^(a[141] & b[74])^(a[140] & b[75])^(a[139] & b[76])^(a[138] & b[77])^(a[137] & b[78])^(a[136] & b[79])^(a[135] & b[80])^(a[134] & b[81])^(a[133] & b[82])^(a[132] & b[83])^(a[131] & b[84])^(a[130] & b[85])^(a[129] & b[86])^(a[128] & b[87])^(a[127] & b[88])^(a[126] & b[89])^(a[125] & b[90])^(a[124] & b[91])^(a[123] & b[92])^(a[122] & b[93])^(a[121] & b[94])^(a[120] & b[95])^(a[119] & b[96])^(a[118] & b[97])^(a[117] & b[98])^(a[116] & b[99])^(a[115] & b[100])^(a[114] & b[101])^(a[113] & b[102])^(a[112] & b[103])^(a[111] & b[104])^(a[110] & b[105])^(a[109] & b[106])^(a[108] & b[107])^(a[107] & b[108])^(a[106] & b[109])^(a[105] & b[110])^(a[104] & b[111])^(a[103] & b[112])^(a[102] & b[113])^(a[101] & b[114])^(a[100] & b[115])^(a[99] & b[116])^(a[98] & b[117])^(a[97] & b[118])^(a[96] & b[119])^(a[95] & b[120])^(a[94] & b[121])^(a[93] & b[122])^(a[92] & b[123])^(a[91] & b[124])^(a[90] & b[125])^(a[89] & b[126])^(a[88] & b[127])^(a[87] & b[128])^(a[86] & b[129])^(a[85] & b[130])^(a[84] & b[131])^(a[83] & b[132])^(a[82] & b[133])^(a[81] & b[134])^(a[80] & b[135])^(a[79] & b[136])^(a[78] & b[137])^(a[77] & b[138])^(a[76] & b[139])^(a[75] & b[140])^(a[74] & b[141])^(a[73] & b[142])^(a[72] & b[143])^(a[71] & b[144])^(a[70] & b[145])^(a[69] & b[146])^(a[68] & b[147])^(a[67] & b[148])^(a[66] & b[149])^(a[65] & b[150])^(a[64] & b[151])^(a[63] & b[152])^(a[62] & b[153])^(a[61] & b[154])^(a[60] & b[155])^(a[59] & b[156])^(a[58] & b[157])^(a[57] & b[158])^(a[56] & b[159])^(a[55] & b[160])^(a[54] & b[161])^(a[53] & b[162])^(a[52] & b[163])^(a[51] & b[164])^(a[50] & b[165])^(a[49] & b[166])^(a[48] & b[167])^(a[47] & b[168])^(a[46] & b[169])^(a[45] & b[170])^(a[44] & b[171])^(a[43] & b[172])^(a[42] & b[173])^(a[41] & b[174])^(a[40] & b[175])^(a[39] & b[176])^(a[38] & b[177])^(a[37] & b[178])^(a[36] & b[179])^(a[35] & b[180])^(a[34] & b[181])^(a[33] & b[182])^(a[32] & b[183])^(a[31] & b[184])^(a[30] & b[185])^(a[29] & b[186])^(a[28] & b[187])^(a[27] & b[188])^(a[26] & b[189])^(a[25] & b[190])^(a[24] & b[191])^(a[23] & b[192])^(a[22] & b[193])^(a[21] & b[194])^(a[20] & b[195])^(a[19] & b[196])^(a[18] & b[197])^(a[17] & b[198])^(a[16] & b[199])^(a[15] & b[200])^(a[14] & b[201])^(a[13] & b[202])^(a[12] & b[203])^(a[11] & b[204])^(a[10] & b[205])^(a[9] & b[206])^(a[8] & b[207])^(a[7] & b[208])^(a[6] & b[209])^(a[5] & b[210])^(a[4] & b[211])^(a[3] & b[212])^(a[2] & b[213])^(a[1] & b[214])^(a[0] & b[215]);
assign y[216] = (a[216] & b[0])^(a[215] & b[1])^(a[214] & b[2])^(a[213] & b[3])^(a[212] & b[4])^(a[211] & b[5])^(a[210] & b[6])^(a[209] & b[7])^(a[208] & b[8])^(a[207] & b[9])^(a[206] & b[10])^(a[205] & b[11])^(a[204] & b[12])^(a[203] & b[13])^(a[202] & b[14])^(a[201] & b[15])^(a[200] & b[16])^(a[199] & b[17])^(a[198] & b[18])^(a[197] & b[19])^(a[196] & b[20])^(a[195] & b[21])^(a[194] & b[22])^(a[193] & b[23])^(a[192] & b[24])^(a[191] & b[25])^(a[190] & b[26])^(a[189] & b[27])^(a[188] & b[28])^(a[187] & b[29])^(a[186] & b[30])^(a[185] & b[31])^(a[184] & b[32])^(a[183] & b[33])^(a[182] & b[34])^(a[181] & b[35])^(a[180] & b[36])^(a[179] & b[37])^(a[178] & b[38])^(a[177] & b[39])^(a[176] & b[40])^(a[175] & b[41])^(a[174] & b[42])^(a[173] & b[43])^(a[172] & b[44])^(a[171] & b[45])^(a[170] & b[46])^(a[169] & b[47])^(a[168] & b[48])^(a[167] & b[49])^(a[166] & b[50])^(a[165] & b[51])^(a[164] & b[52])^(a[163] & b[53])^(a[162] & b[54])^(a[161] & b[55])^(a[160] & b[56])^(a[159] & b[57])^(a[158] & b[58])^(a[157] & b[59])^(a[156] & b[60])^(a[155] & b[61])^(a[154] & b[62])^(a[153] & b[63])^(a[152] & b[64])^(a[151] & b[65])^(a[150] & b[66])^(a[149] & b[67])^(a[148] & b[68])^(a[147] & b[69])^(a[146] & b[70])^(a[145] & b[71])^(a[144] & b[72])^(a[143] & b[73])^(a[142] & b[74])^(a[141] & b[75])^(a[140] & b[76])^(a[139] & b[77])^(a[138] & b[78])^(a[137] & b[79])^(a[136] & b[80])^(a[135] & b[81])^(a[134] & b[82])^(a[133] & b[83])^(a[132] & b[84])^(a[131] & b[85])^(a[130] & b[86])^(a[129] & b[87])^(a[128] & b[88])^(a[127] & b[89])^(a[126] & b[90])^(a[125] & b[91])^(a[124] & b[92])^(a[123] & b[93])^(a[122] & b[94])^(a[121] & b[95])^(a[120] & b[96])^(a[119] & b[97])^(a[118] & b[98])^(a[117] & b[99])^(a[116] & b[100])^(a[115] & b[101])^(a[114] & b[102])^(a[113] & b[103])^(a[112] & b[104])^(a[111] & b[105])^(a[110] & b[106])^(a[109] & b[107])^(a[108] & b[108])^(a[107] & b[109])^(a[106] & b[110])^(a[105] & b[111])^(a[104] & b[112])^(a[103] & b[113])^(a[102] & b[114])^(a[101] & b[115])^(a[100] & b[116])^(a[99] & b[117])^(a[98] & b[118])^(a[97] & b[119])^(a[96] & b[120])^(a[95] & b[121])^(a[94] & b[122])^(a[93] & b[123])^(a[92] & b[124])^(a[91] & b[125])^(a[90] & b[126])^(a[89] & b[127])^(a[88] & b[128])^(a[87] & b[129])^(a[86] & b[130])^(a[85] & b[131])^(a[84] & b[132])^(a[83] & b[133])^(a[82] & b[134])^(a[81] & b[135])^(a[80] & b[136])^(a[79] & b[137])^(a[78] & b[138])^(a[77] & b[139])^(a[76] & b[140])^(a[75] & b[141])^(a[74] & b[142])^(a[73] & b[143])^(a[72] & b[144])^(a[71] & b[145])^(a[70] & b[146])^(a[69] & b[147])^(a[68] & b[148])^(a[67] & b[149])^(a[66] & b[150])^(a[65] & b[151])^(a[64] & b[152])^(a[63] & b[153])^(a[62] & b[154])^(a[61] & b[155])^(a[60] & b[156])^(a[59] & b[157])^(a[58] & b[158])^(a[57] & b[159])^(a[56] & b[160])^(a[55] & b[161])^(a[54] & b[162])^(a[53] & b[163])^(a[52] & b[164])^(a[51] & b[165])^(a[50] & b[166])^(a[49] & b[167])^(a[48] & b[168])^(a[47] & b[169])^(a[46] & b[170])^(a[45] & b[171])^(a[44] & b[172])^(a[43] & b[173])^(a[42] & b[174])^(a[41] & b[175])^(a[40] & b[176])^(a[39] & b[177])^(a[38] & b[178])^(a[37] & b[179])^(a[36] & b[180])^(a[35] & b[181])^(a[34] & b[182])^(a[33] & b[183])^(a[32] & b[184])^(a[31] & b[185])^(a[30] & b[186])^(a[29] & b[187])^(a[28] & b[188])^(a[27] & b[189])^(a[26] & b[190])^(a[25] & b[191])^(a[24] & b[192])^(a[23] & b[193])^(a[22] & b[194])^(a[21] & b[195])^(a[20] & b[196])^(a[19] & b[197])^(a[18] & b[198])^(a[17] & b[199])^(a[16] & b[200])^(a[15] & b[201])^(a[14] & b[202])^(a[13] & b[203])^(a[12] & b[204])^(a[11] & b[205])^(a[10] & b[206])^(a[9] & b[207])^(a[8] & b[208])^(a[7] & b[209])^(a[6] & b[210])^(a[5] & b[211])^(a[4] & b[212])^(a[3] & b[213])^(a[2] & b[214])^(a[1] & b[215])^(a[0] & b[216]);
assign y[217] = (a[217] & b[0])^(a[216] & b[1])^(a[215] & b[2])^(a[214] & b[3])^(a[213] & b[4])^(a[212] & b[5])^(a[211] & b[6])^(a[210] & b[7])^(a[209] & b[8])^(a[208] & b[9])^(a[207] & b[10])^(a[206] & b[11])^(a[205] & b[12])^(a[204] & b[13])^(a[203] & b[14])^(a[202] & b[15])^(a[201] & b[16])^(a[200] & b[17])^(a[199] & b[18])^(a[198] & b[19])^(a[197] & b[20])^(a[196] & b[21])^(a[195] & b[22])^(a[194] & b[23])^(a[193] & b[24])^(a[192] & b[25])^(a[191] & b[26])^(a[190] & b[27])^(a[189] & b[28])^(a[188] & b[29])^(a[187] & b[30])^(a[186] & b[31])^(a[185] & b[32])^(a[184] & b[33])^(a[183] & b[34])^(a[182] & b[35])^(a[181] & b[36])^(a[180] & b[37])^(a[179] & b[38])^(a[178] & b[39])^(a[177] & b[40])^(a[176] & b[41])^(a[175] & b[42])^(a[174] & b[43])^(a[173] & b[44])^(a[172] & b[45])^(a[171] & b[46])^(a[170] & b[47])^(a[169] & b[48])^(a[168] & b[49])^(a[167] & b[50])^(a[166] & b[51])^(a[165] & b[52])^(a[164] & b[53])^(a[163] & b[54])^(a[162] & b[55])^(a[161] & b[56])^(a[160] & b[57])^(a[159] & b[58])^(a[158] & b[59])^(a[157] & b[60])^(a[156] & b[61])^(a[155] & b[62])^(a[154] & b[63])^(a[153] & b[64])^(a[152] & b[65])^(a[151] & b[66])^(a[150] & b[67])^(a[149] & b[68])^(a[148] & b[69])^(a[147] & b[70])^(a[146] & b[71])^(a[145] & b[72])^(a[144] & b[73])^(a[143] & b[74])^(a[142] & b[75])^(a[141] & b[76])^(a[140] & b[77])^(a[139] & b[78])^(a[138] & b[79])^(a[137] & b[80])^(a[136] & b[81])^(a[135] & b[82])^(a[134] & b[83])^(a[133] & b[84])^(a[132] & b[85])^(a[131] & b[86])^(a[130] & b[87])^(a[129] & b[88])^(a[128] & b[89])^(a[127] & b[90])^(a[126] & b[91])^(a[125] & b[92])^(a[124] & b[93])^(a[123] & b[94])^(a[122] & b[95])^(a[121] & b[96])^(a[120] & b[97])^(a[119] & b[98])^(a[118] & b[99])^(a[117] & b[100])^(a[116] & b[101])^(a[115] & b[102])^(a[114] & b[103])^(a[113] & b[104])^(a[112] & b[105])^(a[111] & b[106])^(a[110] & b[107])^(a[109] & b[108])^(a[108] & b[109])^(a[107] & b[110])^(a[106] & b[111])^(a[105] & b[112])^(a[104] & b[113])^(a[103] & b[114])^(a[102] & b[115])^(a[101] & b[116])^(a[100] & b[117])^(a[99] & b[118])^(a[98] & b[119])^(a[97] & b[120])^(a[96] & b[121])^(a[95] & b[122])^(a[94] & b[123])^(a[93] & b[124])^(a[92] & b[125])^(a[91] & b[126])^(a[90] & b[127])^(a[89] & b[128])^(a[88] & b[129])^(a[87] & b[130])^(a[86] & b[131])^(a[85] & b[132])^(a[84] & b[133])^(a[83] & b[134])^(a[82] & b[135])^(a[81] & b[136])^(a[80] & b[137])^(a[79] & b[138])^(a[78] & b[139])^(a[77] & b[140])^(a[76] & b[141])^(a[75] & b[142])^(a[74] & b[143])^(a[73] & b[144])^(a[72] & b[145])^(a[71] & b[146])^(a[70] & b[147])^(a[69] & b[148])^(a[68] & b[149])^(a[67] & b[150])^(a[66] & b[151])^(a[65] & b[152])^(a[64] & b[153])^(a[63] & b[154])^(a[62] & b[155])^(a[61] & b[156])^(a[60] & b[157])^(a[59] & b[158])^(a[58] & b[159])^(a[57] & b[160])^(a[56] & b[161])^(a[55] & b[162])^(a[54] & b[163])^(a[53] & b[164])^(a[52] & b[165])^(a[51] & b[166])^(a[50] & b[167])^(a[49] & b[168])^(a[48] & b[169])^(a[47] & b[170])^(a[46] & b[171])^(a[45] & b[172])^(a[44] & b[173])^(a[43] & b[174])^(a[42] & b[175])^(a[41] & b[176])^(a[40] & b[177])^(a[39] & b[178])^(a[38] & b[179])^(a[37] & b[180])^(a[36] & b[181])^(a[35] & b[182])^(a[34] & b[183])^(a[33] & b[184])^(a[32] & b[185])^(a[31] & b[186])^(a[30] & b[187])^(a[29] & b[188])^(a[28] & b[189])^(a[27] & b[190])^(a[26] & b[191])^(a[25] & b[192])^(a[24] & b[193])^(a[23] & b[194])^(a[22] & b[195])^(a[21] & b[196])^(a[20] & b[197])^(a[19] & b[198])^(a[18] & b[199])^(a[17] & b[200])^(a[16] & b[201])^(a[15] & b[202])^(a[14] & b[203])^(a[13] & b[204])^(a[12] & b[205])^(a[11] & b[206])^(a[10] & b[207])^(a[9] & b[208])^(a[8] & b[209])^(a[7] & b[210])^(a[6] & b[211])^(a[5] & b[212])^(a[4] & b[213])^(a[3] & b[214])^(a[2] & b[215])^(a[1] & b[216])^(a[0] & b[217]);
assign y[218] = (a[218] & b[0])^(a[217] & b[1])^(a[216] & b[2])^(a[215] & b[3])^(a[214] & b[4])^(a[213] & b[5])^(a[212] & b[6])^(a[211] & b[7])^(a[210] & b[8])^(a[209] & b[9])^(a[208] & b[10])^(a[207] & b[11])^(a[206] & b[12])^(a[205] & b[13])^(a[204] & b[14])^(a[203] & b[15])^(a[202] & b[16])^(a[201] & b[17])^(a[200] & b[18])^(a[199] & b[19])^(a[198] & b[20])^(a[197] & b[21])^(a[196] & b[22])^(a[195] & b[23])^(a[194] & b[24])^(a[193] & b[25])^(a[192] & b[26])^(a[191] & b[27])^(a[190] & b[28])^(a[189] & b[29])^(a[188] & b[30])^(a[187] & b[31])^(a[186] & b[32])^(a[185] & b[33])^(a[184] & b[34])^(a[183] & b[35])^(a[182] & b[36])^(a[181] & b[37])^(a[180] & b[38])^(a[179] & b[39])^(a[178] & b[40])^(a[177] & b[41])^(a[176] & b[42])^(a[175] & b[43])^(a[174] & b[44])^(a[173] & b[45])^(a[172] & b[46])^(a[171] & b[47])^(a[170] & b[48])^(a[169] & b[49])^(a[168] & b[50])^(a[167] & b[51])^(a[166] & b[52])^(a[165] & b[53])^(a[164] & b[54])^(a[163] & b[55])^(a[162] & b[56])^(a[161] & b[57])^(a[160] & b[58])^(a[159] & b[59])^(a[158] & b[60])^(a[157] & b[61])^(a[156] & b[62])^(a[155] & b[63])^(a[154] & b[64])^(a[153] & b[65])^(a[152] & b[66])^(a[151] & b[67])^(a[150] & b[68])^(a[149] & b[69])^(a[148] & b[70])^(a[147] & b[71])^(a[146] & b[72])^(a[145] & b[73])^(a[144] & b[74])^(a[143] & b[75])^(a[142] & b[76])^(a[141] & b[77])^(a[140] & b[78])^(a[139] & b[79])^(a[138] & b[80])^(a[137] & b[81])^(a[136] & b[82])^(a[135] & b[83])^(a[134] & b[84])^(a[133] & b[85])^(a[132] & b[86])^(a[131] & b[87])^(a[130] & b[88])^(a[129] & b[89])^(a[128] & b[90])^(a[127] & b[91])^(a[126] & b[92])^(a[125] & b[93])^(a[124] & b[94])^(a[123] & b[95])^(a[122] & b[96])^(a[121] & b[97])^(a[120] & b[98])^(a[119] & b[99])^(a[118] & b[100])^(a[117] & b[101])^(a[116] & b[102])^(a[115] & b[103])^(a[114] & b[104])^(a[113] & b[105])^(a[112] & b[106])^(a[111] & b[107])^(a[110] & b[108])^(a[109] & b[109])^(a[108] & b[110])^(a[107] & b[111])^(a[106] & b[112])^(a[105] & b[113])^(a[104] & b[114])^(a[103] & b[115])^(a[102] & b[116])^(a[101] & b[117])^(a[100] & b[118])^(a[99] & b[119])^(a[98] & b[120])^(a[97] & b[121])^(a[96] & b[122])^(a[95] & b[123])^(a[94] & b[124])^(a[93] & b[125])^(a[92] & b[126])^(a[91] & b[127])^(a[90] & b[128])^(a[89] & b[129])^(a[88] & b[130])^(a[87] & b[131])^(a[86] & b[132])^(a[85] & b[133])^(a[84] & b[134])^(a[83] & b[135])^(a[82] & b[136])^(a[81] & b[137])^(a[80] & b[138])^(a[79] & b[139])^(a[78] & b[140])^(a[77] & b[141])^(a[76] & b[142])^(a[75] & b[143])^(a[74] & b[144])^(a[73] & b[145])^(a[72] & b[146])^(a[71] & b[147])^(a[70] & b[148])^(a[69] & b[149])^(a[68] & b[150])^(a[67] & b[151])^(a[66] & b[152])^(a[65] & b[153])^(a[64] & b[154])^(a[63] & b[155])^(a[62] & b[156])^(a[61] & b[157])^(a[60] & b[158])^(a[59] & b[159])^(a[58] & b[160])^(a[57] & b[161])^(a[56] & b[162])^(a[55] & b[163])^(a[54] & b[164])^(a[53] & b[165])^(a[52] & b[166])^(a[51] & b[167])^(a[50] & b[168])^(a[49] & b[169])^(a[48] & b[170])^(a[47] & b[171])^(a[46] & b[172])^(a[45] & b[173])^(a[44] & b[174])^(a[43] & b[175])^(a[42] & b[176])^(a[41] & b[177])^(a[40] & b[178])^(a[39] & b[179])^(a[38] & b[180])^(a[37] & b[181])^(a[36] & b[182])^(a[35] & b[183])^(a[34] & b[184])^(a[33] & b[185])^(a[32] & b[186])^(a[31] & b[187])^(a[30] & b[188])^(a[29] & b[189])^(a[28] & b[190])^(a[27] & b[191])^(a[26] & b[192])^(a[25] & b[193])^(a[24] & b[194])^(a[23] & b[195])^(a[22] & b[196])^(a[21] & b[197])^(a[20] & b[198])^(a[19] & b[199])^(a[18] & b[200])^(a[17] & b[201])^(a[16] & b[202])^(a[15] & b[203])^(a[14] & b[204])^(a[13] & b[205])^(a[12] & b[206])^(a[11] & b[207])^(a[10] & b[208])^(a[9] & b[209])^(a[8] & b[210])^(a[7] & b[211])^(a[6] & b[212])^(a[5] & b[213])^(a[4] & b[214])^(a[3] & b[215])^(a[2] & b[216])^(a[1] & b[217])^(a[0] & b[218]);
assign y[219] = (a[219] & b[0])^(a[218] & b[1])^(a[217] & b[2])^(a[216] & b[3])^(a[215] & b[4])^(a[214] & b[5])^(a[213] & b[6])^(a[212] & b[7])^(a[211] & b[8])^(a[210] & b[9])^(a[209] & b[10])^(a[208] & b[11])^(a[207] & b[12])^(a[206] & b[13])^(a[205] & b[14])^(a[204] & b[15])^(a[203] & b[16])^(a[202] & b[17])^(a[201] & b[18])^(a[200] & b[19])^(a[199] & b[20])^(a[198] & b[21])^(a[197] & b[22])^(a[196] & b[23])^(a[195] & b[24])^(a[194] & b[25])^(a[193] & b[26])^(a[192] & b[27])^(a[191] & b[28])^(a[190] & b[29])^(a[189] & b[30])^(a[188] & b[31])^(a[187] & b[32])^(a[186] & b[33])^(a[185] & b[34])^(a[184] & b[35])^(a[183] & b[36])^(a[182] & b[37])^(a[181] & b[38])^(a[180] & b[39])^(a[179] & b[40])^(a[178] & b[41])^(a[177] & b[42])^(a[176] & b[43])^(a[175] & b[44])^(a[174] & b[45])^(a[173] & b[46])^(a[172] & b[47])^(a[171] & b[48])^(a[170] & b[49])^(a[169] & b[50])^(a[168] & b[51])^(a[167] & b[52])^(a[166] & b[53])^(a[165] & b[54])^(a[164] & b[55])^(a[163] & b[56])^(a[162] & b[57])^(a[161] & b[58])^(a[160] & b[59])^(a[159] & b[60])^(a[158] & b[61])^(a[157] & b[62])^(a[156] & b[63])^(a[155] & b[64])^(a[154] & b[65])^(a[153] & b[66])^(a[152] & b[67])^(a[151] & b[68])^(a[150] & b[69])^(a[149] & b[70])^(a[148] & b[71])^(a[147] & b[72])^(a[146] & b[73])^(a[145] & b[74])^(a[144] & b[75])^(a[143] & b[76])^(a[142] & b[77])^(a[141] & b[78])^(a[140] & b[79])^(a[139] & b[80])^(a[138] & b[81])^(a[137] & b[82])^(a[136] & b[83])^(a[135] & b[84])^(a[134] & b[85])^(a[133] & b[86])^(a[132] & b[87])^(a[131] & b[88])^(a[130] & b[89])^(a[129] & b[90])^(a[128] & b[91])^(a[127] & b[92])^(a[126] & b[93])^(a[125] & b[94])^(a[124] & b[95])^(a[123] & b[96])^(a[122] & b[97])^(a[121] & b[98])^(a[120] & b[99])^(a[119] & b[100])^(a[118] & b[101])^(a[117] & b[102])^(a[116] & b[103])^(a[115] & b[104])^(a[114] & b[105])^(a[113] & b[106])^(a[112] & b[107])^(a[111] & b[108])^(a[110] & b[109])^(a[109] & b[110])^(a[108] & b[111])^(a[107] & b[112])^(a[106] & b[113])^(a[105] & b[114])^(a[104] & b[115])^(a[103] & b[116])^(a[102] & b[117])^(a[101] & b[118])^(a[100] & b[119])^(a[99] & b[120])^(a[98] & b[121])^(a[97] & b[122])^(a[96] & b[123])^(a[95] & b[124])^(a[94] & b[125])^(a[93] & b[126])^(a[92] & b[127])^(a[91] & b[128])^(a[90] & b[129])^(a[89] & b[130])^(a[88] & b[131])^(a[87] & b[132])^(a[86] & b[133])^(a[85] & b[134])^(a[84] & b[135])^(a[83] & b[136])^(a[82] & b[137])^(a[81] & b[138])^(a[80] & b[139])^(a[79] & b[140])^(a[78] & b[141])^(a[77] & b[142])^(a[76] & b[143])^(a[75] & b[144])^(a[74] & b[145])^(a[73] & b[146])^(a[72] & b[147])^(a[71] & b[148])^(a[70] & b[149])^(a[69] & b[150])^(a[68] & b[151])^(a[67] & b[152])^(a[66] & b[153])^(a[65] & b[154])^(a[64] & b[155])^(a[63] & b[156])^(a[62] & b[157])^(a[61] & b[158])^(a[60] & b[159])^(a[59] & b[160])^(a[58] & b[161])^(a[57] & b[162])^(a[56] & b[163])^(a[55] & b[164])^(a[54] & b[165])^(a[53] & b[166])^(a[52] & b[167])^(a[51] & b[168])^(a[50] & b[169])^(a[49] & b[170])^(a[48] & b[171])^(a[47] & b[172])^(a[46] & b[173])^(a[45] & b[174])^(a[44] & b[175])^(a[43] & b[176])^(a[42] & b[177])^(a[41] & b[178])^(a[40] & b[179])^(a[39] & b[180])^(a[38] & b[181])^(a[37] & b[182])^(a[36] & b[183])^(a[35] & b[184])^(a[34] & b[185])^(a[33] & b[186])^(a[32] & b[187])^(a[31] & b[188])^(a[30] & b[189])^(a[29] & b[190])^(a[28] & b[191])^(a[27] & b[192])^(a[26] & b[193])^(a[25] & b[194])^(a[24] & b[195])^(a[23] & b[196])^(a[22] & b[197])^(a[21] & b[198])^(a[20] & b[199])^(a[19] & b[200])^(a[18] & b[201])^(a[17] & b[202])^(a[16] & b[203])^(a[15] & b[204])^(a[14] & b[205])^(a[13] & b[206])^(a[12] & b[207])^(a[11] & b[208])^(a[10] & b[209])^(a[9] & b[210])^(a[8] & b[211])^(a[7] & b[212])^(a[6] & b[213])^(a[5] & b[214])^(a[4] & b[215])^(a[3] & b[216])^(a[2] & b[217])^(a[1] & b[218])^(a[0] & b[219]);
assign y[220] = (a[220] & b[0])^(a[219] & b[1])^(a[218] & b[2])^(a[217] & b[3])^(a[216] & b[4])^(a[215] & b[5])^(a[214] & b[6])^(a[213] & b[7])^(a[212] & b[8])^(a[211] & b[9])^(a[210] & b[10])^(a[209] & b[11])^(a[208] & b[12])^(a[207] & b[13])^(a[206] & b[14])^(a[205] & b[15])^(a[204] & b[16])^(a[203] & b[17])^(a[202] & b[18])^(a[201] & b[19])^(a[200] & b[20])^(a[199] & b[21])^(a[198] & b[22])^(a[197] & b[23])^(a[196] & b[24])^(a[195] & b[25])^(a[194] & b[26])^(a[193] & b[27])^(a[192] & b[28])^(a[191] & b[29])^(a[190] & b[30])^(a[189] & b[31])^(a[188] & b[32])^(a[187] & b[33])^(a[186] & b[34])^(a[185] & b[35])^(a[184] & b[36])^(a[183] & b[37])^(a[182] & b[38])^(a[181] & b[39])^(a[180] & b[40])^(a[179] & b[41])^(a[178] & b[42])^(a[177] & b[43])^(a[176] & b[44])^(a[175] & b[45])^(a[174] & b[46])^(a[173] & b[47])^(a[172] & b[48])^(a[171] & b[49])^(a[170] & b[50])^(a[169] & b[51])^(a[168] & b[52])^(a[167] & b[53])^(a[166] & b[54])^(a[165] & b[55])^(a[164] & b[56])^(a[163] & b[57])^(a[162] & b[58])^(a[161] & b[59])^(a[160] & b[60])^(a[159] & b[61])^(a[158] & b[62])^(a[157] & b[63])^(a[156] & b[64])^(a[155] & b[65])^(a[154] & b[66])^(a[153] & b[67])^(a[152] & b[68])^(a[151] & b[69])^(a[150] & b[70])^(a[149] & b[71])^(a[148] & b[72])^(a[147] & b[73])^(a[146] & b[74])^(a[145] & b[75])^(a[144] & b[76])^(a[143] & b[77])^(a[142] & b[78])^(a[141] & b[79])^(a[140] & b[80])^(a[139] & b[81])^(a[138] & b[82])^(a[137] & b[83])^(a[136] & b[84])^(a[135] & b[85])^(a[134] & b[86])^(a[133] & b[87])^(a[132] & b[88])^(a[131] & b[89])^(a[130] & b[90])^(a[129] & b[91])^(a[128] & b[92])^(a[127] & b[93])^(a[126] & b[94])^(a[125] & b[95])^(a[124] & b[96])^(a[123] & b[97])^(a[122] & b[98])^(a[121] & b[99])^(a[120] & b[100])^(a[119] & b[101])^(a[118] & b[102])^(a[117] & b[103])^(a[116] & b[104])^(a[115] & b[105])^(a[114] & b[106])^(a[113] & b[107])^(a[112] & b[108])^(a[111] & b[109])^(a[110] & b[110])^(a[109] & b[111])^(a[108] & b[112])^(a[107] & b[113])^(a[106] & b[114])^(a[105] & b[115])^(a[104] & b[116])^(a[103] & b[117])^(a[102] & b[118])^(a[101] & b[119])^(a[100] & b[120])^(a[99] & b[121])^(a[98] & b[122])^(a[97] & b[123])^(a[96] & b[124])^(a[95] & b[125])^(a[94] & b[126])^(a[93] & b[127])^(a[92] & b[128])^(a[91] & b[129])^(a[90] & b[130])^(a[89] & b[131])^(a[88] & b[132])^(a[87] & b[133])^(a[86] & b[134])^(a[85] & b[135])^(a[84] & b[136])^(a[83] & b[137])^(a[82] & b[138])^(a[81] & b[139])^(a[80] & b[140])^(a[79] & b[141])^(a[78] & b[142])^(a[77] & b[143])^(a[76] & b[144])^(a[75] & b[145])^(a[74] & b[146])^(a[73] & b[147])^(a[72] & b[148])^(a[71] & b[149])^(a[70] & b[150])^(a[69] & b[151])^(a[68] & b[152])^(a[67] & b[153])^(a[66] & b[154])^(a[65] & b[155])^(a[64] & b[156])^(a[63] & b[157])^(a[62] & b[158])^(a[61] & b[159])^(a[60] & b[160])^(a[59] & b[161])^(a[58] & b[162])^(a[57] & b[163])^(a[56] & b[164])^(a[55] & b[165])^(a[54] & b[166])^(a[53] & b[167])^(a[52] & b[168])^(a[51] & b[169])^(a[50] & b[170])^(a[49] & b[171])^(a[48] & b[172])^(a[47] & b[173])^(a[46] & b[174])^(a[45] & b[175])^(a[44] & b[176])^(a[43] & b[177])^(a[42] & b[178])^(a[41] & b[179])^(a[40] & b[180])^(a[39] & b[181])^(a[38] & b[182])^(a[37] & b[183])^(a[36] & b[184])^(a[35] & b[185])^(a[34] & b[186])^(a[33] & b[187])^(a[32] & b[188])^(a[31] & b[189])^(a[30] & b[190])^(a[29] & b[191])^(a[28] & b[192])^(a[27] & b[193])^(a[26] & b[194])^(a[25] & b[195])^(a[24] & b[196])^(a[23] & b[197])^(a[22] & b[198])^(a[21] & b[199])^(a[20] & b[200])^(a[19] & b[201])^(a[18] & b[202])^(a[17] & b[203])^(a[16] & b[204])^(a[15] & b[205])^(a[14] & b[206])^(a[13] & b[207])^(a[12] & b[208])^(a[11] & b[209])^(a[10] & b[210])^(a[9] & b[211])^(a[8] & b[212])^(a[7] & b[213])^(a[6] & b[214])^(a[5] & b[215])^(a[4] & b[216])^(a[3] & b[217])^(a[2] & b[218])^(a[1] & b[219])^(a[0] & b[220]);
assign y[221] = (a[221] & b[0])^(a[220] & b[1])^(a[219] & b[2])^(a[218] & b[3])^(a[217] & b[4])^(a[216] & b[5])^(a[215] & b[6])^(a[214] & b[7])^(a[213] & b[8])^(a[212] & b[9])^(a[211] & b[10])^(a[210] & b[11])^(a[209] & b[12])^(a[208] & b[13])^(a[207] & b[14])^(a[206] & b[15])^(a[205] & b[16])^(a[204] & b[17])^(a[203] & b[18])^(a[202] & b[19])^(a[201] & b[20])^(a[200] & b[21])^(a[199] & b[22])^(a[198] & b[23])^(a[197] & b[24])^(a[196] & b[25])^(a[195] & b[26])^(a[194] & b[27])^(a[193] & b[28])^(a[192] & b[29])^(a[191] & b[30])^(a[190] & b[31])^(a[189] & b[32])^(a[188] & b[33])^(a[187] & b[34])^(a[186] & b[35])^(a[185] & b[36])^(a[184] & b[37])^(a[183] & b[38])^(a[182] & b[39])^(a[181] & b[40])^(a[180] & b[41])^(a[179] & b[42])^(a[178] & b[43])^(a[177] & b[44])^(a[176] & b[45])^(a[175] & b[46])^(a[174] & b[47])^(a[173] & b[48])^(a[172] & b[49])^(a[171] & b[50])^(a[170] & b[51])^(a[169] & b[52])^(a[168] & b[53])^(a[167] & b[54])^(a[166] & b[55])^(a[165] & b[56])^(a[164] & b[57])^(a[163] & b[58])^(a[162] & b[59])^(a[161] & b[60])^(a[160] & b[61])^(a[159] & b[62])^(a[158] & b[63])^(a[157] & b[64])^(a[156] & b[65])^(a[155] & b[66])^(a[154] & b[67])^(a[153] & b[68])^(a[152] & b[69])^(a[151] & b[70])^(a[150] & b[71])^(a[149] & b[72])^(a[148] & b[73])^(a[147] & b[74])^(a[146] & b[75])^(a[145] & b[76])^(a[144] & b[77])^(a[143] & b[78])^(a[142] & b[79])^(a[141] & b[80])^(a[140] & b[81])^(a[139] & b[82])^(a[138] & b[83])^(a[137] & b[84])^(a[136] & b[85])^(a[135] & b[86])^(a[134] & b[87])^(a[133] & b[88])^(a[132] & b[89])^(a[131] & b[90])^(a[130] & b[91])^(a[129] & b[92])^(a[128] & b[93])^(a[127] & b[94])^(a[126] & b[95])^(a[125] & b[96])^(a[124] & b[97])^(a[123] & b[98])^(a[122] & b[99])^(a[121] & b[100])^(a[120] & b[101])^(a[119] & b[102])^(a[118] & b[103])^(a[117] & b[104])^(a[116] & b[105])^(a[115] & b[106])^(a[114] & b[107])^(a[113] & b[108])^(a[112] & b[109])^(a[111] & b[110])^(a[110] & b[111])^(a[109] & b[112])^(a[108] & b[113])^(a[107] & b[114])^(a[106] & b[115])^(a[105] & b[116])^(a[104] & b[117])^(a[103] & b[118])^(a[102] & b[119])^(a[101] & b[120])^(a[100] & b[121])^(a[99] & b[122])^(a[98] & b[123])^(a[97] & b[124])^(a[96] & b[125])^(a[95] & b[126])^(a[94] & b[127])^(a[93] & b[128])^(a[92] & b[129])^(a[91] & b[130])^(a[90] & b[131])^(a[89] & b[132])^(a[88] & b[133])^(a[87] & b[134])^(a[86] & b[135])^(a[85] & b[136])^(a[84] & b[137])^(a[83] & b[138])^(a[82] & b[139])^(a[81] & b[140])^(a[80] & b[141])^(a[79] & b[142])^(a[78] & b[143])^(a[77] & b[144])^(a[76] & b[145])^(a[75] & b[146])^(a[74] & b[147])^(a[73] & b[148])^(a[72] & b[149])^(a[71] & b[150])^(a[70] & b[151])^(a[69] & b[152])^(a[68] & b[153])^(a[67] & b[154])^(a[66] & b[155])^(a[65] & b[156])^(a[64] & b[157])^(a[63] & b[158])^(a[62] & b[159])^(a[61] & b[160])^(a[60] & b[161])^(a[59] & b[162])^(a[58] & b[163])^(a[57] & b[164])^(a[56] & b[165])^(a[55] & b[166])^(a[54] & b[167])^(a[53] & b[168])^(a[52] & b[169])^(a[51] & b[170])^(a[50] & b[171])^(a[49] & b[172])^(a[48] & b[173])^(a[47] & b[174])^(a[46] & b[175])^(a[45] & b[176])^(a[44] & b[177])^(a[43] & b[178])^(a[42] & b[179])^(a[41] & b[180])^(a[40] & b[181])^(a[39] & b[182])^(a[38] & b[183])^(a[37] & b[184])^(a[36] & b[185])^(a[35] & b[186])^(a[34] & b[187])^(a[33] & b[188])^(a[32] & b[189])^(a[31] & b[190])^(a[30] & b[191])^(a[29] & b[192])^(a[28] & b[193])^(a[27] & b[194])^(a[26] & b[195])^(a[25] & b[196])^(a[24] & b[197])^(a[23] & b[198])^(a[22] & b[199])^(a[21] & b[200])^(a[20] & b[201])^(a[19] & b[202])^(a[18] & b[203])^(a[17] & b[204])^(a[16] & b[205])^(a[15] & b[206])^(a[14] & b[207])^(a[13] & b[208])^(a[12] & b[209])^(a[11] & b[210])^(a[10] & b[211])^(a[9] & b[212])^(a[8] & b[213])^(a[7] & b[214])^(a[6] & b[215])^(a[5] & b[216])^(a[4] & b[217])^(a[3] & b[218])^(a[2] & b[219])^(a[1] & b[220])^(a[0] & b[221]);
assign y[222] = (a[222] & b[0])^(a[221] & b[1])^(a[220] & b[2])^(a[219] & b[3])^(a[218] & b[4])^(a[217] & b[5])^(a[216] & b[6])^(a[215] & b[7])^(a[214] & b[8])^(a[213] & b[9])^(a[212] & b[10])^(a[211] & b[11])^(a[210] & b[12])^(a[209] & b[13])^(a[208] & b[14])^(a[207] & b[15])^(a[206] & b[16])^(a[205] & b[17])^(a[204] & b[18])^(a[203] & b[19])^(a[202] & b[20])^(a[201] & b[21])^(a[200] & b[22])^(a[199] & b[23])^(a[198] & b[24])^(a[197] & b[25])^(a[196] & b[26])^(a[195] & b[27])^(a[194] & b[28])^(a[193] & b[29])^(a[192] & b[30])^(a[191] & b[31])^(a[190] & b[32])^(a[189] & b[33])^(a[188] & b[34])^(a[187] & b[35])^(a[186] & b[36])^(a[185] & b[37])^(a[184] & b[38])^(a[183] & b[39])^(a[182] & b[40])^(a[181] & b[41])^(a[180] & b[42])^(a[179] & b[43])^(a[178] & b[44])^(a[177] & b[45])^(a[176] & b[46])^(a[175] & b[47])^(a[174] & b[48])^(a[173] & b[49])^(a[172] & b[50])^(a[171] & b[51])^(a[170] & b[52])^(a[169] & b[53])^(a[168] & b[54])^(a[167] & b[55])^(a[166] & b[56])^(a[165] & b[57])^(a[164] & b[58])^(a[163] & b[59])^(a[162] & b[60])^(a[161] & b[61])^(a[160] & b[62])^(a[159] & b[63])^(a[158] & b[64])^(a[157] & b[65])^(a[156] & b[66])^(a[155] & b[67])^(a[154] & b[68])^(a[153] & b[69])^(a[152] & b[70])^(a[151] & b[71])^(a[150] & b[72])^(a[149] & b[73])^(a[148] & b[74])^(a[147] & b[75])^(a[146] & b[76])^(a[145] & b[77])^(a[144] & b[78])^(a[143] & b[79])^(a[142] & b[80])^(a[141] & b[81])^(a[140] & b[82])^(a[139] & b[83])^(a[138] & b[84])^(a[137] & b[85])^(a[136] & b[86])^(a[135] & b[87])^(a[134] & b[88])^(a[133] & b[89])^(a[132] & b[90])^(a[131] & b[91])^(a[130] & b[92])^(a[129] & b[93])^(a[128] & b[94])^(a[127] & b[95])^(a[126] & b[96])^(a[125] & b[97])^(a[124] & b[98])^(a[123] & b[99])^(a[122] & b[100])^(a[121] & b[101])^(a[120] & b[102])^(a[119] & b[103])^(a[118] & b[104])^(a[117] & b[105])^(a[116] & b[106])^(a[115] & b[107])^(a[114] & b[108])^(a[113] & b[109])^(a[112] & b[110])^(a[111] & b[111])^(a[110] & b[112])^(a[109] & b[113])^(a[108] & b[114])^(a[107] & b[115])^(a[106] & b[116])^(a[105] & b[117])^(a[104] & b[118])^(a[103] & b[119])^(a[102] & b[120])^(a[101] & b[121])^(a[100] & b[122])^(a[99] & b[123])^(a[98] & b[124])^(a[97] & b[125])^(a[96] & b[126])^(a[95] & b[127])^(a[94] & b[128])^(a[93] & b[129])^(a[92] & b[130])^(a[91] & b[131])^(a[90] & b[132])^(a[89] & b[133])^(a[88] & b[134])^(a[87] & b[135])^(a[86] & b[136])^(a[85] & b[137])^(a[84] & b[138])^(a[83] & b[139])^(a[82] & b[140])^(a[81] & b[141])^(a[80] & b[142])^(a[79] & b[143])^(a[78] & b[144])^(a[77] & b[145])^(a[76] & b[146])^(a[75] & b[147])^(a[74] & b[148])^(a[73] & b[149])^(a[72] & b[150])^(a[71] & b[151])^(a[70] & b[152])^(a[69] & b[153])^(a[68] & b[154])^(a[67] & b[155])^(a[66] & b[156])^(a[65] & b[157])^(a[64] & b[158])^(a[63] & b[159])^(a[62] & b[160])^(a[61] & b[161])^(a[60] & b[162])^(a[59] & b[163])^(a[58] & b[164])^(a[57] & b[165])^(a[56] & b[166])^(a[55] & b[167])^(a[54] & b[168])^(a[53] & b[169])^(a[52] & b[170])^(a[51] & b[171])^(a[50] & b[172])^(a[49] & b[173])^(a[48] & b[174])^(a[47] & b[175])^(a[46] & b[176])^(a[45] & b[177])^(a[44] & b[178])^(a[43] & b[179])^(a[42] & b[180])^(a[41] & b[181])^(a[40] & b[182])^(a[39] & b[183])^(a[38] & b[184])^(a[37] & b[185])^(a[36] & b[186])^(a[35] & b[187])^(a[34] & b[188])^(a[33] & b[189])^(a[32] & b[190])^(a[31] & b[191])^(a[30] & b[192])^(a[29] & b[193])^(a[28] & b[194])^(a[27] & b[195])^(a[26] & b[196])^(a[25] & b[197])^(a[24] & b[198])^(a[23] & b[199])^(a[22] & b[200])^(a[21] & b[201])^(a[20] & b[202])^(a[19] & b[203])^(a[18] & b[204])^(a[17] & b[205])^(a[16] & b[206])^(a[15] & b[207])^(a[14] & b[208])^(a[13] & b[209])^(a[12] & b[210])^(a[11] & b[211])^(a[10] & b[212])^(a[9] & b[213])^(a[8] & b[214])^(a[7] & b[215])^(a[6] & b[216])^(a[5] & b[217])^(a[4] & b[218])^(a[3] & b[219])^(a[2] & b[220])^(a[1] & b[221])^(a[0] & b[222]);
assign y[223] = (a[223] & b[0])^(a[222] & b[1])^(a[221] & b[2])^(a[220] & b[3])^(a[219] & b[4])^(a[218] & b[5])^(a[217] & b[6])^(a[216] & b[7])^(a[215] & b[8])^(a[214] & b[9])^(a[213] & b[10])^(a[212] & b[11])^(a[211] & b[12])^(a[210] & b[13])^(a[209] & b[14])^(a[208] & b[15])^(a[207] & b[16])^(a[206] & b[17])^(a[205] & b[18])^(a[204] & b[19])^(a[203] & b[20])^(a[202] & b[21])^(a[201] & b[22])^(a[200] & b[23])^(a[199] & b[24])^(a[198] & b[25])^(a[197] & b[26])^(a[196] & b[27])^(a[195] & b[28])^(a[194] & b[29])^(a[193] & b[30])^(a[192] & b[31])^(a[191] & b[32])^(a[190] & b[33])^(a[189] & b[34])^(a[188] & b[35])^(a[187] & b[36])^(a[186] & b[37])^(a[185] & b[38])^(a[184] & b[39])^(a[183] & b[40])^(a[182] & b[41])^(a[181] & b[42])^(a[180] & b[43])^(a[179] & b[44])^(a[178] & b[45])^(a[177] & b[46])^(a[176] & b[47])^(a[175] & b[48])^(a[174] & b[49])^(a[173] & b[50])^(a[172] & b[51])^(a[171] & b[52])^(a[170] & b[53])^(a[169] & b[54])^(a[168] & b[55])^(a[167] & b[56])^(a[166] & b[57])^(a[165] & b[58])^(a[164] & b[59])^(a[163] & b[60])^(a[162] & b[61])^(a[161] & b[62])^(a[160] & b[63])^(a[159] & b[64])^(a[158] & b[65])^(a[157] & b[66])^(a[156] & b[67])^(a[155] & b[68])^(a[154] & b[69])^(a[153] & b[70])^(a[152] & b[71])^(a[151] & b[72])^(a[150] & b[73])^(a[149] & b[74])^(a[148] & b[75])^(a[147] & b[76])^(a[146] & b[77])^(a[145] & b[78])^(a[144] & b[79])^(a[143] & b[80])^(a[142] & b[81])^(a[141] & b[82])^(a[140] & b[83])^(a[139] & b[84])^(a[138] & b[85])^(a[137] & b[86])^(a[136] & b[87])^(a[135] & b[88])^(a[134] & b[89])^(a[133] & b[90])^(a[132] & b[91])^(a[131] & b[92])^(a[130] & b[93])^(a[129] & b[94])^(a[128] & b[95])^(a[127] & b[96])^(a[126] & b[97])^(a[125] & b[98])^(a[124] & b[99])^(a[123] & b[100])^(a[122] & b[101])^(a[121] & b[102])^(a[120] & b[103])^(a[119] & b[104])^(a[118] & b[105])^(a[117] & b[106])^(a[116] & b[107])^(a[115] & b[108])^(a[114] & b[109])^(a[113] & b[110])^(a[112] & b[111])^(a[111] & b[112])^(a[110] & b[113])^(a[109] & b[114])^(a[108] & b[115])^(a[107] & b[116])^(a[106] & b[117])^(a[105] & b[118])^(a[104] & b[119])^(a[103] & b[120])^(a[102] & b[121])^(a[101] & b[122])^(a[100] & b[123])^(a[99] & b[124])^(a[98] & b[125])^(a[97] & b[126])^(a[96] & b[127])^(a[95] & b[128])^(a[94] & b[129])^(a[93] & b[130])^(a[92] & b[131])^(a[91] & b[132])^(a[90] & b[133])^(a[89] & b[134])^(a[88] & b[135])^(a[87] & b[136])^(a[86] & b[137])^(a[85] & b[138])^(a[84] & b[139])^(a[83] & b[140])^(a[82] & b[141])^(a[81] & b[142])^(a[80] & b[143])^(a[79] & b[144])^(a[78] & b[145])^(a[77] & b[146])^(a[76] & b[147])^(a[75] & b[148])^(a[74] & b[149])^(a[73] & b[150])^(a[72] & b[151])^(a[71] & b[152])^(a[70] & b[153])^(a[69] & b[154])^(a[68] & b[155])^(a[67] & b[156])^(a[66] & b[157])^(a[65] & b[158])^(a[64] & b[159])^(a[63] & b[160])^(a[62] & b[161])^(a[61] & b[162])^(a[60] & b[163])^(a[59] & b[164])^(a[58] & b[165])^(a[57] & b[166])^(a[56] & b[167])^(a[55] & b[168])^(a[54] & b[169])^(a[53] & b[170])^(a[52] & b[171])^(a[51] & b[172])^(a[50] & b[173])^(a[49] & b[174])^(a[48] & b[175])^(a[47] & b[176])^(a[46] & b[177])^(a[45] & b[178])^(a[44] & b[179])^(a[43] & b[180])^(a[42] & b[181])^(a[41] & b[182])^(a[40] & b[183])^(a[39] & b[184])^(a[38] & b[185])^(a[37] & b[186])^(a[36] & b[187])^(a[35] & b[188])^(a[34] & b[189])^(a[33] & b[190])^(a[32] & b[191])^(a[31] & b[192])^(a[30] & b[193])^(a[29] & b[194])^(a[28] & b[195])^(a[27] & b[196])^(a[26] & b[197])^(a[25] & b[198])^(a[24] & b[199])^(a[23] & b[200])^(a[22] & b[201])^(a[21] & b[202])^(a[20] & b[203])^(a[19] & b[204])^(a[18] & b[205])^(a[17] & b[206])^(a[16] & b[207])^(a[15] & b[208])^(a[14] & b[209])^(a[13] & b[210])^(a[12] & b[211])^(a[11] & b[212])^(a[10] & b[213])^(a[9] & b[214])^(a[8] & b[215])^(a[7] & b[216])^(a[6] & b[217])^(a[5] & b[218])^(a[4] & b[219])^(a[3] & b[220])^(a[2] & b[221])^(a[1] & b[222])^(a[0] & b[223]);
assign y[224] = (a[224] & b[0])^(a[223] & b[1])^(a[222] & b[2])^(a[221] & b[3])^(a[220] & b[4])^(a[219] & b[5])^(a[218] & b[6])^(a[217] & b[7])^(a[216] & b[8])^(a[215] & b[9])^(a[214] & b[10])^(a[213] & b[11])^(a[212] & b[12])^(a[211] & b[13])^(a[210] & b[14])^(a[209] & b[15])^(a[208] & b[16])^(a[207] & b[17])^(a[206] & b[18])^(a[205] & b[19])^(a[204] & b[20])^(a[203] & b[21])^(a[202] & b[22])^(a[201] & b[23])^(a[200] & b[24])^(a[199] & b[25])^(a[198] & b[26])^(a[197] & b[27])^(a[196] & b[28])^(a[195] & b[29])^(a[194] & b[30])^(a[193] & b[31])^(a[192] & b[32])^(a[191] & b[33])^(a[190] & b[34])^(a[189] & b[35])^(a[188] & b[36])^(a[187] & b[37])^(a[186] & b[38])^(a[185] & b[39])^(a[184] & b[40])^(a[183] & b[41])^(a[182] & b[42])^(a[181] & b[43])^(a[180] & b[44])^(a[179] & b[45])^(a[178] & b[46])^(a[177] & b[47])^(a[176] & b[48])^(a[175] & b[49])^(a[174] & b[50])^(a[173] & b[51])^(a[172] & b[52])^(a[171] & b[53])^(a[170] & b[54])^(a[169] & b[55])^(a[168] & b[56])^(a[167] & b[57])^(a[166] & b[58])^(a[165] & b[59])^(a[164] & b[60])^(a[163] & b[61])^(a[162] & b[62])^(a[161] & b[63])^(a[160] & b[64])^(a[159] & b[65])^(a[158] & b[66])^(a[157] & b[67])^(a[156] & b[68])^(a[155] & b[69])^(a[154] & b[70])^(a[153] & b[71])^(a[152] & b[72])^(a[151] & b[73])^(a[150] & b[74])^(a[149] & b[75])^(a[148] & b[76])^(a[147] & b[77])^(a[146] & b[78])^(a[145] & b[79])^(a[144] & b[80])^(a[143] & b[81])^(a[142] & b[82])^(a[141] & b[83])^(a[140] & b[84])^(a[139] & b[85])^(a[138] & b[86])^(a[137] & b[87])^(a[136] & b[88])^(a[135] & b[89])^(a[134] & b[90])^(a[133] & b[91])^(a[132] & b[92])^(a[131] & b[93])^(a[130] & b[94])^(a[129] & b[95])^(a[128] & b[96])^(a[127] & b[97])^(a[126] & b[98])^(a[125] & b[99])^(a[124] & b[100])^(a[123] & b[101])^(a[122] & b[102])^(a[121] & b[103])^(a[120] & b[104])^(a[119] & b[105])^(a[118] & b[106])^(a[117] & b[107])^(a[116] & b[108])^(a[115] & b[109])^(a[114] & b[110])^(a[113] & b[111])^(a[112] & b[112])^(a[111] & b[113])^(a[110] & b[114])^(a[109] & b[115])^(a[108] & b[116])^(a[107] & b[117])^(a[106] & b[118])^(a[105] & b[119])^(a[104] & b[120])^(a[103] & b[121])^(a[102] & b[122])^(a[101] & b[123])^(a[100] & b[124])^(a[99] & b[125])^(a[98] & b[126])^(a[97] & b[127])^(a[96] & b[128])^(a[95] & b[129])^(a[94] & b[130])^(a[93] & b[131])^(a[92] & b[132])^(a[91] & b[133])^(a[90] & b[134])^(a[89] & b[135])^(a[88] & b[136])^(a[87] & b[137])^(a[86] & b[138])^(a[85] & b[139])^(a[84] & b[140])^(a[83] & b[141])^(a[82] & b[142])^(a[81] & b[143])^(a[80] & b[144])^(a[79] & b[145])^(a[78] & b[146])^(a[77] & b[147])^(a[76] & b[148])^(a[75] & b[149])^(a[74] & b[150])^(a[73] & b[151])^(a[72] & b[152])^(a[71] & b[153])^(a[70] & b[154])^(a[69] & b[155])^(a[68] & b[156])^(a[67] & b[157])^(a[66] & b[158])^(a[65] & b[159])^(a[64] & b[160])^(a[63] & b[161])^(a[62] & b[162])^(a[61] & b[163])^(a[60] & b[164])^(a[59] & b[165])^(a[58] & b[166])^(a[57] & b[167])^(a[56] & b[168])^(a[55] & b[169])^(a[54] & b[170])^(a[53] & b[171])^(a[52] & b[172])^(a[51] & b[173])^(a[50] & b[174])^(a[49] & b[175])^(a[48] & b[176])^(a[47] & b[177])^(a[46] & b[178])^(a[45] & b[179])^(a[44] & b[180])^(a[43] & b[181])^(a[42] & b[182])^(a[41] & b[183])^(a[40] & b[184])^(a[39] & b[185])^(a[38] & b[186])^(a[37] & b[187])^(a[36] & b[188])^(a[35] & b[189])^(a[34] & b[190])^(a[33] & b[191])^(a[32] & b[192])^(a[31] & b[193])^(a[30] & b[194])^(a[29] & b[195])^(a[28] & b[196])^(a[27] & b[197])^(a[26] & b[198])^(a[25] & b[199])^(a[24] & b[200])^(a[23] & b[201])^(a[22] & b[202])^(a[21] & b[203])^(a[20] & b[204])^(a[19] & b[205])^(a[18] & b[206])^(a[17] & b[207])^(a[16] & b[208])^(a[15] & b[209])^(a[14] & b[210])^(a[13] & b[211])^(a[12] & b[212])^(a[11] & b[213])^(a[10] & b[214])^(a[9] & b[215])^(a[8] & b[216])^(a[7] & b[217])^(a[6] & b[218])^(a[5] & b[219])^(a[4] & b[220])^(a[3] & b[221])^(a[2] & b[222])^(a[1] & b[223])^(a[0] & b[224]);
assign y[225] = (a[225] & b[0])^(a[224] & b[1])^(a[223] & b[2])^(a[222] & b[3])^(a[221] & b[4])^(a[220] & b[5])^(a[219] & b[6])^(a[218] & b[7])^(a[217] & b[8])^(a[216] & b[9])^(a[215] & b[10])^(a[214] & b[11])^(a[213] & b[12])^(a[212] & b[13])^(a[211] & b[14])^(a[210] & b[15])^(a[209] & b[16])^(a[208] & b[17])^(a[207] & b[18])^(a[206] & b[19])^(a[205] & b[20])^(a[204] & b[21])^(a[203] & b[22])^(a[202] & b[23])^(a[201] & b[24])^(a[200] & b[25])^(a[199] & b[26])^(a[198] & b[27])^(a[197] & b[28])^(a[196] & b[29])^(a[195] & b[30])^(a[194] & b[31])^(a[193] & b[32])^(a[192] & b[33])^(a[191] & b[34])^(a[190] & b[35])^(a[189] & b[36])^(a[188] & b[37])^(a[187] & b[38])^(a[186] & b[39])^(a[185] & b[40])^(a[184] & b[41])^(a[183] & b[42])^(a[182] & b[43])^(a[181] & b[44])^(a[180] & b[45])^(a[179] & b[46])^(a[178] & b[47])^(a[177] & b[48])^(a[176] & b[49])^(a[175] & b[50])^(a[174] & b[51])^(a[173] & b[52])^(a[172] & b[53])^(a[171] & b[54])^(a[170] & b[55])^(a[169] & b[56])^(a[168] & b[57])^(a[167] & b[58])^(a[166] & b[59])^(a[165] & b[60])^(a[164] & b[61])^(a[163] & b[62])^(a[162] & b[63])^(a[161] & b[64])^(a[160] & b[65])^(a[159] & b[66])^(a[158] & b[67])^(a[157] & b[68])^(a[156] & b[69])^(a[155] & b[70])^(a[154] & b[71])^(a[153] & b[72])^(a[152] & b[73])^(a[151] & b[74])^(a[150] & b[75])^(a[149] & b[76])^(a[148] & b[77])^(a[147] & b[78])^(a[146] & b[79])^(a[145] & b[80])^(a[144] & b[81])^(a[143] & b[82])^(a[142] & b[83])^(a[141] & b[84])^(a[140] & b[85])^(a[139] & b[86])^(a[138] & b[87])^(a[137] & b[88])^(a[136] & b[89])^(a[135] & b[90])^(a[134] & b[91])^(a[133] & b[92])^(a[132] & b[93])^(a[131] & b[94])^(a[130] & b[95])^(a[129] & b[96])^(a[128] & b[97])^(a[127] & b[98])^(a[126] & b[99])^(a[125] & b[100])^(a[124] & b[101])^(a[123] & b[102])^(a[122] & b[103])^(a[121] & b[104])^(a[120] & b[105])^(a[119] & b[106])^(a[118] & b[107])^(a[117] & b[108])^(a[116] & b[109])^(a[115] & b[110])^(a[114] & b[111])^(a[113] & b[112])^(a[112] & b[113])^(a[111] & b[114])^(a[110] & b[115])^(a[109] & b[116])^(a[108] & b[117])^(a[107] & b[118])^(a[106] & b[119])^(a[105] & b[120])^(a[104] & b[121])^(a[103] & b[122])^(a[102] & b[123])^(a[101] & b[124])^(a[100] & b[125])^(a[99] & b[126])^(a[98] & b[127])^(a[97] & b[128])^(a[96] & b[129])^(a[95] & b[130])^(a[94] & b[131])^(a[93] & b[132])^(a[92] & b[133])^(a[91] & b[134])^(a[90] & b[135])^(a[89] & b[136])^(a[88] & b[137])^(a[87] & b[138])^(a[86] & b[139])^(a[85] & b[140])^(a[84] & b[141])^(a[83] & b[142])^(a[82] & b[143])^(a[81] & b[144])^(a[80] & b[145])^(a[79] & b[146])^(a[78] & b[147])^(a[77] & b[148])^(a[76] & b[149])^(a[75] & b[150])^(a[74] & b[151])^(a[73] & b[152])^(a[72] & b[153])^(a[71] & b[154])^(a[70] & b[155])^(a[69] & b[156])^(a[68] & b[157])^(a[67] & b[158])^(a[66] & b[159])^(a[65] & b[160])^(a[64] & b[161])^(a[63] & b[162])^(a[62] & b[163])^(a[61] & b[164])^(a[60] & b[165])^(a[59] & b[166])^(a[58] & b[167])^(a[57] & b[168])^(a[56] & b[169])^(a[55] & b[170])^(a[54] & b[171])^(a[53] & b[172])^(a[52] & b[173])^(a[51] & b[174])^(a[50] & b[175])^(a[49] & b[176])^(a[48] & b[177])^(a[47] & b[178])^(a[46] & b[179])^(a[45] & b[180])^(a[44] & b[181])^(a[43] & b[182])^(a[42] & b[183])^(a[41] & b[184])^(a[40] & b[185])^(a[39] & b[186])^(a[38] & b[187])^(a[37] & b[188])^(a[36] & b[189])^(a[35] & b[190])^(a[34] & b[191])^(a[33] & b[192])^(a[32] & b[193])^(a[31] & b[194])^(a[30] & b[195])^(a[29] & b[196])^(a[28] & b[197])^(a[27] & b[198])^(a[26] & b[199])^(a[25] & b[200])^(a[24] & b[201])^(a[23] & b[202])^(a[22] & b[203])^(a[21] & b[204])^(a[20] & b[205])^(a[19] & b[206])^(a[18] & b[207])^(a[17] & b[208])^(a[16] & b[209])^(a[15] & b[210])^(a[14] & b[211])^(a[13] & b[212])^(a[12] & b[213])^(a[11] & b[214])^(a[10] & b[215])^(a[9] & b[216])^(a[8] & b[217])^(a[7] & b[218])^(a[6] & b[219])^(a[5] & b[220])^(a[4] & b[221])^(a[3] & b[222])^(a[2] & b[223])^(a[1] & b[224])^(a[0] & b[225]);
assign y[226] = (a[226] & b[0])^(a[225] & b[1])^(a[224] & b[2])^(a[223] & b[3])^(a[222] & b[4])^(a[221] & b[5])^(a[220] & b[6])^(a[219] & b[7])^(a[218] & b[8])^(a[217] & b[9])^(a[216] & b[10])^(a[215] & b[11])^(a[214] & b[12])^(a[213] & b[13])^(a[212] & b[14])^(a[211] & b[15])^(a[210] & b[16])^(a[209] & b[17])^(a[208] & b[18])^(a[207] & b[19])^(a[206] & b[20])^(a[205] & b[21])^(a[204] & b[22])^(a[203] & b[23])^(a[202] & b[24])^(a[201] & b[25])^(a[200] & b[26])^(a[199] & b[27])^(a[198] & b[28])^(a[197] & b[29])^(a[196] & b[30])^(a[195] & b[31])^(a[194] & b[32])^(a[193] & b[33])^(a[192] & b[34])^(a[191] & b[35])^(a[190] & b[36])^(a[189] & b[37])^(a[188] & b[38])^(a[187] & b[39])^(a[186] & b[40])^(a[185] & b[41])^(a[184] & b[42])^(a[183] & b[43])^(a[182] & b[44])^(a[181] & b[45])^(a[180] & b[46])^(a[179] & b[47])^(a[178] & b[48])^(a[177] & b[49])^(a[176] & b[50])^(a[175] & b[51])^(a[174] & b[52])^(a[173] & b[53])^(a[172] & b[54])^(a[171] & b[55])^(a[170] & b[56])^(a[169] & b[57])^(a[168] & b[58])^(a[167] & b[59])^(a[166] & b[60])^(a[165] & b[61])^(a[164] & b[62])^(a[163] & b[63])^(a[162] & b[64])^(a[161] & b[65])^(a[160] & b[66])^(a[159] & b[67])^(a[158] & b[68])^(a[157] & b[69])^(a[156] & b[70])^(a[155] & b[71])^(a[154] & b[72])^(a[153] & b[73])^(a[152] & b[74])^(a[151] & b[75])^(a[150] & b[76])^(a[149] & b[77])^(a[148] & b[78])^(a[147] & b[79])^(a[146] & b[80])^(a[145] & b[81])^(a[144] & b[82])^(a[143] & b[83])^(a[142] & b[84])^(a[141] & b[85])^(a[140] & b[86])^(a[139] & b[87])^(a[138] & b[88])^(a[137] & b[89])^(a[136] & b[90])^(a[135] & b[91])^(a[134] & b[92])^(a[133] & b[93])^(a[132] & b[94])^(a[131] & b[95])^(a[130] & b[96])^(a[129] & b[97])^(a[128] & b[98])^(a[127] & b[99])^(a[126] & b[100])^(a[125] & b[101])^(a[124] & b[102])^(a[123] & b[103])^(a[122] & b[104])^(a[121] & b[105])^(a[120] & b[106])^(a[119] & b[107])^(a[118] & b[108])^(a[117] & b[109])^(a[116] & b[110])^(a[115] & b[111])^(a[114] & b[112])^(a[113] & b[113])^(a[112] & b[114])^(a[111] & b[115])^(a[110] & b[116])^(a[109] & b[117])^(a[108] & b[118])^(a[107] & b[119])^(a[106] & b[120])^(a[105] & b[121])^(a[104] & b[122])^(a[103] & b[123])^(a[102] & b[124])^(a[101] & b[125])^(a[100] & b[126])^(a[99] & b[127])^(a[98] & b[128])^(a[97] & b[129])^(a[96] & b[130])^(a[95] & b[131])^(a[94] & b[132])^(a[93] & b[133])^(a[92] & b[134])^(a[91] & b[135])^(a[90] & b[136])^(a[89] & b[137])^(a[88] & b[138])^(a[87] & b[139])^(a[86] & b[140])^(a[85] & b[141])^(a[84] & b[142])^(a[83] & b[143])^(a[82] & b[144])^(a[81] & b[145])^(a[80] & b[146])^(a[79] & b[147])^(a[78] & b[148])^(a[77] & b[149])^(a[76] & b[150])^(a[75] & b[151])^(a[74] & b[152])^(a[73] & b[153])^(a[72] & b[154])^(a[71] & b[155])^(a[70] & b[156])^(a[69] & b[157])^(a[68] & b[158])^(a[67] & b[159])^(a[66] & b[160])^(a[65] & b[161])^(a[64] & b[162])^(a[63] & b[163])^(a[62] & b[164])^(a[61] & b[165])^(a[60] & b[166])^(a[59] & b[167])^(a[58] & b[168])^(a[57] & b[169])^(a[56] & b[170])^(a[55] & b[171])^(a[54] & b[172])^(a[53] & b[173])^(a[52] & b[174])^(a[51] & b[175])^(a[50] & b[176])^(a[49] & b[177])^(a[48] & b[178])^(a[47] & b[179])^(a[46] & b[180])^(a[45] & b[181])^(a[44] & b[182])^(a[43] & b[183])^(a[42] & b[184])^(a[41] & b[185])^(a[40] & b[186])^(a[39] & b[187])^(a[38] & b[188])^(a[37] & b[189])^(a[36] & b[190])^(a[35] & b[191])^(a[34] & b[192])^(a[33] & b[193])^(a[32] & b[194])^(a[31] & b[195])^(a[30] & b[196])^(a[29] & b[197])^(a[28] & b[198])^(a[27] & b[199])^(a[26] & b[200])^(a[25] & b[201])^(a[24] & b[202])^(a[23] & b[203])^(a[22] & b[204])^(a[21] & b[205])^(a[20] & b[206])^(a[19] & b[207])^(a[18] & b[208])^(a[17] & b[209])^(a[16] & b[210])^(a[15] & b[211])^(a[14] & b[212])^(a[13] & b[213])^(a[12] & b[214])^(a[11] & b[215])^(a[10] & b[216])^(a[9] & b[217])^(a[8] & b[218])^(a[7] & b[219])^(a[6] & b[220])^(a[5] & b[221])^(a[4] & b[222])^(a[3] & b[223])^(a[2] & b[224])^(a[1] & b[225])^(a[0] & b[226]);
assign y[227] = (a[227] & b[0])^(a[226] & b[1])^(a[225] & b[2])^(a[224] & b[3])^(a[223] & b[4])^(a[222] & b[5])^(a[221] & b[6])^(a[220] & b[7])^(a[219] & b[8])^(a[218] & b[9])^(a[217] & b[10])^(a[216] & b[11])^(a[215] & b[12])^(a[214] & b[13])^(a[213] & b[14])^(a[212] & b[15])^(a[211] & b[16])^(a[210] & b[17])^(a[209] & b[18])^(a[208] & b[19])^(a[207] & b[20])^(a[206] & b[21])^(a[205] & b[22])^(a[204] & b[23])^(a[203] & b[24])^(a[202] & b[25])^(a[201] & b[26])^(a[200] & b[27])^(a[199] & b[28])^(a[198] & b[29])^(a[197] & b[30])^(a[196] & b[31])^(a[195] & b[32])^(a[194] & b[33])^(a[193] & b[34])^(a[192] & b[35])^(a[191] & b[36])^(a[190] & b[37])^(a[189] & b[38])^(a[188] & b[39])^(a[187] & b[40])^(a[186] & b[41])^(a[185] & b[42])^(a[184] & b[43])^(a[183] & b[44])^(a[182] & b[45])^(a[181] & b[46])^(a[180] & b[47])^(a[179] & b[48])^(a[178] & b[49])^(a[177] & b[50])^(a[176] & b[51])^(a[175] & b[52])^(a[174] & b[53])^(a[173] & b[54])^(a[172] & b[55])^(a[171] & b[56])^(a[170] & b[57])^(a[169] & b[58])^(a[168] & b[59])^(a[167] & b[60])^(a[166] & b[61])^(a[165] & b[62])^(a[164] & b[63])^(a[163] & b[64])^(a[162] & b[65])^(a[161] & b[66])^(a[160] & b[67])^(a[159] & b[68])^(a[158] & b[69])^(a[157] & b[70])^(a[156] & b[71])^(a[155] & b[72])^(a[154] & b[73])^(a[153] & b[74])^(a[152] & b[75])^(a[151] & b[76])^(a[150] & b[77])^(a[149] & b[78])^(a[148] & b[79])^(a[147] & b[80])^(a[146] & b[81])^(a[145] & b[82])^(a[144] & b[83])^(a[143] & b[84])^(a[142] & b[85])^(a[141] & b[86])^(a[140] & b[87])^(a[139] & b[88])^(a[138] & b[89])^(a[137] & b[90])^(a[136] & b[91])^(a[135] & b[92])^(a[134] & b[93])^(a[133] & b[94])^(a[132] & b[95])^(a[131] & b[96])^(a[130] & b[97])^(a[129] & b[98])^(a[128] & b[99])^(a[127] & b[100])^(a[126] & b[101])^(a[125] & b[102])^(a[124] & b[103])^(a[123] & b[104])^(a[122] & b[105])^(a[121] & b[106])^(a[120] & b[107])^(a[119] & b[108])^(a[118] & b[109])^(a[117] & b[110])^(a[116] & b[111])^(a[115] & b[112])^(a[114] & b[113])^(a[113] & b[114])^(a[112] & b[115])^(a[111] & b[116])^(a[110] & b[117])^(a[109] & b[118])^(a[108] & b[119])^(a[107] & b[120])^(a[106] & b[121])^(a[105] & b[122])^(a[104] & b[123])^(a[103] & b[124])^(a[102] & b[125])^(a[101] & b[126])^(a[100] & b[127])^(a[99] & b[128])^(a[98] & b[129])^(a[97] & b[130])^(a[96] & b[131])^(a[95] & b[132])^(a[94] & b[133])^(a[93] & b[134])^(a[92] & b[135])^(a[91] & b[136])^(a[90] & b[137])^(a[89] & b[138])^(a[88] & b[139])^(a[87] & b[140])^(a[86] & b[141])^(a[85] & b[142])^(a[84] & b[143])^(a[83] & b[144])^(a[82] & b[145])^(a[81] & b[146])^(a[80] & b[147])^(a[79] & b[148])^(a[78] & b[149])^(a[77] & b[150])^(a[76] & b[151])^(a[75] & b[152])^(a[74] & b[153])^(a[73] & b[154])^(a[72] & b[155])^(a[71] & b[156])^(a[70] & b[157])^(a[69] & b[158])^(a[68] & b[159])^(a[67] & b[160])^(a[66] & b[161])^(a[65] & b[162])^(a[64] & b[163])^(a[63] & b[164])^(a[62] & b[165])^(a[61] & b[166])^(a[60] & b[167])^(a[59] & b[168])^(a[58] & b[169])^(a[57] & b[170])^(a[56] & b[171])^(a[55] & b[172])^(a[54] & b[173])^(a[53] & b[174])^(a[52] & b[175])^(a[51] & b[176])^(a[50] & b[177])^(a[49] & b[178])^(a[48] & b[179])^(a[47] & b[180])^(a[46] & b[181])^(a[45] & b[182])^(a[44] & b[183])^(a[43] & b[184])^(a[42] & b[185])^(a[41] & b[186])^(a[40] & b[187])^(a[39] & b[188])^(a[38] & b[189])^(a[37] & b[190])^(a[36] & b[191])^(a[35] & b[192])^(a[34] & b[193])^(a[33] & b[194])^(a[32] & b[195])^(a[31] & b[196])^(a[30] & b[197])^(a[29] & b[198])^(a[28] & b[199])^(a[27] & b[200])^(a[26] & b[201])^(a[25] & b[202])^(a[24] & b[203])^(a[23] & b[204])^(a[22] & b[205])^(a[21] & b[206])^(a[20] & b[207])^(a[19] & b[208])^(a[18] & b[209])^(a[17] & b[210])^(a[16] & b[211])^(a[15] & b[212])^(a[14] & b[213])^(a[13] & b[214])^(a[12] & b[215])^(a[11] & b[216])^(a[10] & b[217])^(a[9] & b[218])^(a[8] & b[219])^(a[7] & b[220])^(a[6] & b[221])^(a[5] & b[222])^(a[4] & b[223])^(a[3] & b[224])^(a[2] & b[225])^(a[1] & b[226])^(a[0] & b[227]);
assign y[228] = (a[228] & b[0])^(a[227] & b[1])^(a[226] & b[2])^(a[225] & b[3])^(a[224] & b[4])^(a[223] & b[5])^(a[222] & b[6])^(a[221] & b[7])^(a[220] & b[8])^(a[219] & b[9])^(a[218] & b[10])^(a[217] & b[11])^(a[216] & b[12])^(a[215] & b[13])^(a[214] & b[14])^(a[213] & b[15])^(a[212] & b[16])^(a[211] & b[17])^(a[210] & b[18])^(a[209] & b[19])^(a[208] & b[20])^(a[207] & b[21])^(a[206] & b[22])^(a[205] & b[23])^(a[204] & b[24])^(a[203] & b[25])^(a[202] & b[26])^(a[201] & b[27])^(a[200] & b[28])^(a[199] & b[29])^(a[198] & b[30])^(a[197] & b[31])^(a[196] & b[32])^(a[195] & b[33])^(a[194] & b[34])^(a[193] & b[35])^(a[192] & b[36])^(a[191] & b[37])^(a[190] & b[38])^(a[189] & b[39])^(a[188] & b[40])^(a[187] & b[41])^(a[186] & b[42])^(a[185] & b[43])^(a[184] & b[44])^(a[183] & b[45])^(a[182] & b[46])^(a[181] & b[47])^(a[180] & b[48])^(a[179] & b[49])^(a[178] & b[50])^(a[177] & b[51])^(a[176] & b[52])^(a[175] & b[53])^(a[174] & b[54])^(a[173] & b[55])^(a[172] & b[56])^(a[171] & b[57])^(a[170] & b[58])^(a[169] & b[59])^(a[168] & b[60])^(a[167] & b[61])^(a[166] & b[62])^(a[165] & b[63])^(a[164] & b[64])^(a[163] & b[65])^(a[162] & b[66])^(a[161] & b[67])^(a[160] & b[68])^(a[159] & b[69])^(a[158] & b[70])^(a[157] & b[71])^(a[156] & b[72])^(a[155] & b[73])^(a[154] & b[74])^(a[153] & b[75])^(a[152] & b[76])^(a[151] & b[77])^(a[150] & b[78])^(a[149] & b[79])^(a[148] & b[80])^(a[147] & b[81])^(a[146] & b[82])^(a[145] & b[83])^(a[144] & b[84])^(a[143] & b[85])^(a[142] & b[86])^(a[141] & b[87])^(a[140] & b[88])^(a[139] & b[89])^(a[138] & b[90])^(a[137] & b[91])^(a[136] & b[92])^(a[135] & b[93])^(a[134] & b[94])^(a[133] & b[95])^(a[132] & b[96])^(a[131] & b[97])^(a[130] & b[98])^(a[129] & b[99])^(a[128] & b[100])^(a[127] & b[101])^(a[126] & b[102])^(a[125] & b[103])^(a[124] & b[104])^(a[123] & b[105])^(a[122] & b[106])^(a[121] & b[107])^(a[120] & b[108])^(a[119] & b[109])^(a[118] & b[110])^(a[117] & b[111])^(a[116] & b[112])^(a[115] & b[113])^(a[114] & b[114])^(a[113] & b[115])^(a[112] & b[116])^(a[111] & b[117])^(a[110] & b[118])^(a[109] & b[119])^(a[108] & b[120])^(a[107] & b[121])^(a[106] & b[122])^(a[105] & b[123])^(a[104] & b[124])^(a[103] & b[125])^(a[102] & b[126])^(a[101] & b[127])^(a[100] & b[128])^(a[99] & b[129])^(a[98] & b[130])^(a[97] & b[131])^(a[96] & b[132])^(a[95] & b[133])^(a[94] & b[134])^(a[93] & b[135])^(a[92] & b[136])^(a[91] & b[137])^(a[90] & b[138])^(a[89] & b[139])^(a[88] & b[140])^(a[87] & b[141])^(a[86] & b[142])^(a[85] & b[143])^(a[84] & b[144])^(a[83] & b[145])^(a[82] & b[146])^(a[81] & b[147])^(a[80] & b[148])^(a[79] & b[149])^(a[78] & b[150])^(a[77] & b[151])^(a[76] & b[152])^(a[75] & b[153])^(a[74] & b[154])^(a[73] & b[155])^(a[72] & b[156])^(a[71] & b[157])^(a[70] & b[158])^(a[69] & b[159])^(a[68] & b[160])^(a[67] & b[161])^(a[66] & b[162])^(a[65] & b[163])^(a[64] & b[164])^(a[63] & b[165])^(a[62] & b[166])^(a[61] & b[167])^(a[60] & b[168])^(a[59] & b[169])^(a[58] & b[170])^(a[57] & b[171])^(a[56] & b[172])^(a[55] & b[173])^(a[54] & b[174])^(a[53] & b[175])^(a[52] & b[176])^(a[51] & b[177])^(a[50] & b[178])^(a[49] & b[179])^(a[48] & b[180])^(a[47] & b[181])^(a[46] & b[182])^(a[45] & b[183])^(a[44] & b[184])^(a[43] & b[185])^(a[42] & b[186])^(a[41] & b[187])^(a[40] & b[188])^(a[39] & b[189])^(a[38] & b[190])^(a[37] & b[191])^(a[36] & b[192])^(a[35] & b[193])^(a[34] & b[194])^(a[33] & b[195])^(a[32] & b[196])^(a[31] & b[197])^(a[30] & b[198])^(a[29] & b[199])^(a[28] & b[200])^(a[27] & b[201])^(a[26] & b[202])^(a[25] & b[203])^(a[24] & b[204])^(a[23] & b[205])^(a[22] & b[206])^(a[21] & b[207])^(a[20] & b[208])^(a[19] & b[209])^(a[18] & b[210])^(a[17] & b[211])^(a[16] & b[212])^(a[15] & b[213])^(a[14] & b[214])^(a[13] & b[215])^(a[12] & b[216])^(a[11] & b[217])^(a[10] & b[218])^(a[9] & b[219])^(a[8] & b[220])^(a[7] & b[221])^(a[6] & b[222])^(a[5] & b[223])^(a[4] & b[224])^(a[3] & b[225])^(a[2] & b[226])^(a[1] & b[227])^(a[0] & b[228]);
assign y[229] = (a[229] & b[0])^(a[228] & b[1])^(a[227] & b[2])^(a[226] & b[3])^(a[225] & b[4])^(a[224] & b[5])^(a[223] & b[6])^(a[222] & b[7])^(a[221] & b[8])^(a[220] & b[9])^(a[219] & b[10])^(a[218] & b[11])^(a[217] & b[12])^(a[216] & b[13])^(a[215] & b[14])^(a[214] & b[15])^(a[213] & b[16])^(a[212] & b[17])^(a[211] & b[18])^(a[210] & b[19])^(a[209] & b[20])^(a[208] & b[21])^(a[207] & b[22])^(a[206] & b[23])^(a[205] & b[24])^(a[204] & b[25])^(a[203] & b[26])^(a[202] & b[27])^(a[201] & b[28])^(a[200] & b[29])^(a[199] & b[30])^(a[198] & b[31])^(a[197] & b[32])^(a[196] & b[33])^(a[195] & b[34])^(a[194] & b[35])^(a[193] & b[36])^(a[192] & b[37])^(a[191] & b[38])^(a[190] & b[39])^(a[189] & b[40])^(a[188] & b[41])^(a[187] & b[42])^(a[186] & b[43])^(a[185] & b[44])^(a[184] & b[45])^(a[183] & b[46])^(a[182] & b[47])^(a[181] & b[48])^(a[180] & b[49])^(a[179] & b[50])^(a[178] & b[51])^(a[177] & b[52])^(a[176] & b[53])^(a[175] & b[54])^(a[174] & b[55])^(a[173] & b[56])^(a[172] & b[57])^(a[171] & b[58])^(a[170] & b[59])^(a[169] & b[60])^(a[168] & b[61])^(a[167] & b[62])^(a[166] & b[63])^(a[165] & b[64])^(a[164] & b[65])^(a[163] & b[66])^(a[162] & b[67])^(a[161] & b[68])^(a[160] & b[69])^(a[159] & b[70])^(a[158] & b[71])^(a[157] & b[72])^(a[156] & b[73])^(a[155] & b[74])^(a[154] & b[75])^(a[153] & b[76])^(a[152] & b[77])^(a[151] & b[78])^(a[150] & b[79])^(a[149] & b[80])^(a[148] & b[81])^(a[147] & b[82])^(a[146] & b[83])^(a[145] & b[84])^(a[144] & b[85])^(a[143] & b[86])^(a[142] & b[87])^(a[141] & b[88])^(a[140] & b[89])^(a[139] & b[90])^(a[138] & b[91])^(a[137] & b[92])^(a[136] & b[93])^(a[135] & b[94])^(a[134] & b[95])^(a[133] & b[96])^(a[132] & b[97])^(a[131] & b[98])^(a[130] & b[99])^(a[129] & b[100])^(a[128] & b[101])^(a[127] & b[102])^(a[126] & b[103])^(a[125] & b[104])^(a[124] & b[105])^(a[123] & b[106])^(a[122] & b[107])^(a[121] & b[108])^(a[120] & b[109])^(a[119] & b[110])^(a[118] & b[111])^(a[117] & b[112])^(a[116] & b[113])^(a[115] & b[114])^(a[114] & b[115])^(a[113] & b[116])^(a[112] & b[117])^(a[111] & b[118])^(a[110] & b[119])^(a[109] & b[120])^(a[108] & b[121])^(a[107] & b[122])^(a[106] & b[123])^(a[105] & b[124])^(a[104] & b[125])^(a[103] & b[126])^(a[102] & b[127])^(a[101] & b[128])^(a[100] & b[129])^(a[99] & b[130])^(a[98] & b[131])^(a[97] & b[132])^(a[96] & b[133])^(a[95] & b[134])^(a[94] & b[135])^(a[93] & b[136])^(a[92] & b[137])^(a[91] & b[138])^(a[90] & b[139])^(a[89] & b[140])^(a[88] & b[141])^(a[87] & b[142])^(a[86] & b[143])^(a[85] & b[144])^(a[84] & b[145])^(a[83] & b[146])^(a[82] & b[147])^(a[81] & b[148])^(a[80] & b[149])^(a[79] & b[150])^(a[78] & b[151])^(a[77] & b[152])^(a[76] & b[153])^(a[75] & b[154])^(a[74] & b[155])^(a[73] & b[156])^(a[72] & b[157])^(a[71] & b[158])^(a[70] & b[159])^(a[69] & b[160])^(a[68] & b[161])^(a[67] & b[162])^(a[66] & b[163])^(a[65] & b[164])^(a[64] & b[165])^(a[63] & b[166])^(a[62] & b[167])^(a[61] & b[168])^(a[60] & b[169])^(a[59] & b[170])^(a[58] & b[171])^(a[57] & b[172])^(a[56] & b[173])^(a[55] & b[174])^(a[54] & b[175])^(a[53] & b[176])^(a[52] & b[177])^(a[51] & b[178])^(a[50] & b[179])^(a[49] & b[180])^(a[48] & b[181])^(a[47] & b[182])^(a[46] & b[183])^(a[45] & b[184])^(a[44] & b[185])^(a[43] & b[186])^(a[42] & b[187])^(a[41] & b[188])^(a[40] & b[189])^(a[39] & b[190])^(a[38] & b[191])^(a[37] & b[192])^(a[36] & b[193])^(a[35] & b[194])^(a[34] & b[195])^(a[33] & b[196])^(a[32] & b[197])^(a[31] & b[198])^(a[30] & b[199])^(a[29] & b[200])^(a[28] & b[201])^(a[27] & b[202])^(a[26] & b[203])^(a[25] & b[204])^(a[24] & b[205])^(a[23] & b[206])^(a[22] & b[207])^(a[21] & b[208])^(a[20] & b[209])^(a[19] & b[210])^(a[18] & b[211])^(a[17] & b[212])^(a[16] & b[213])^(a[15] & b[214])^(a[14] & b[215])^(a[13] & b[216])^(a[12] & b[217])^(a[11] & b[218])^(a[10] & b[219])^(a[9] & b[220])^(a[8] & b[221])^(a[7] & b[222])^(a[6] & b[223])^(a[5] & b[224])^(a[4] & b[225])^(a[3] & b[226])^(a[2] & b[227])^(a[1] & b[228])^(a[0] & b[229]);
assign y[230] = (a[230] & b[0])^(a[229] & b[1])^(a[228] & b[2])^(a[227] & b[3])^(a[226] & b[4])^(a[225] & b[5])^(a[224] & b[6])^(a[223] & b[7])^(a[222] & b[8])^(a[221] & b[9])^(a[220] & b[10])^(a[219] & b[11])^(a[218] & b[12])^(a[217] & b[13])^(a[216] & b[14])^(a[215] & b[15])^(a[214] & b[16])^(a[213] & b[17])^(a[212] & b[18])^(a[211] & b[19])^(a[210] & b[20])^(a[209] & b[21])^(a[208] & b[22])^(a[207] & b[23])^(a[206] & b[24])^(a[205] & b[25])^(a[204] & b[26])^(a[203] & b[27])^(a[202] & b[28])^(a[201] & b[29])^(a[200] & b[30])^(a[199] & b[31])^(a[198] & b[32])^(a[197] & b[33])^(a[196] & b[34])^(a[195] & b[35])^(a[194] & b[36])^(a[193] & b[37])^(a[192] & b[38])^(a[191] & b[39])^(a[190] & b[40])^(a[189] & b[41])^(a[188] & b[42])^(a[187] & b[43])^(a[186] & b[44])^(a[185] & b[45])^(a[184] & b[46])^(a[183] & b[47])^(a[182] & b[48])^(a[181] & b[49])^(a[180] & b[50])^(a[179] & b[51])^(a[178] & b[52])^(a[177] & b[53])^(a[176] & b[54])^(a[175] & b[55])^(a[174] & b[56])^(a[173] & b[57])^(a[172] & b[58])^(a[171] & b[59])^(a[170] & b[60])^(a[169] & b[61])^(a[168] & b[62])^(a[167] & b[63])^(a[166] & b[64])^(a[165] & b[65])^(a[164] & b[66])^(a[163] & b[67])^(a[162] & b[68])^(a[161] & b[69])^(a[160] & b[70])^(a[159] & b[71])^(a[158] & b[72])^(a[157] & b[73])^(a[156] & b[74])^(a[155] & b[75])^(a[154] & b[76])^(a[153] & b[77])^(a[152] & b[78])^(a[151] & b[79])^(a[150] & b[80])^(a[149] & b[81])^(a[148] & b[82])^(a[147] & b[83])^(a[146] & b[84])^(a[145] & b[85])^(a[144] & b[86])^(a[143] & b[87])^(a[142] & b[88])^(a[141] & b[89])^(a[140] & b[90])^(a[139] & b[91])^(a[138] & b[92])^(a[137] & b[93])^(a[136] & b[94])^(a[135] & b[95])^(a[134] & b[96])^(a[133] & b[97])^(a[132] & b[98])^(a[131] & b[99])^(a[130] & b[100])^(a[129] & b[101])^(a[128] & b[102])^(a[127] & b[103])^(a[126] & b[104])^(a[125] & b[105])^(a[124] & b[106])^(a[123] & b[107])^(a[122] & b[108])^(a[121] & b[109])^(a[120] & b[110])^(a[119] & b[111])^(a[118] & b[112])^(a[117] & b[113])^(a[116] & b[114])^(a[115] & b[115])^(a[114] & b[116])^(a[113] & b[117])^(a[112] & b[118])^(a[111] & b[119])^(a[110] & b[120])^(a[109] & b[121])^(a[108] & b[122])^(a[107] & b[123])^(a[106] & b[124])^(a[105] & b[125])^(a[104] & b[126])^(a[103] & b[127])^(a[102] & b[128])^(a[101] & b[129])^(a[100] & b[130])^(a[99] & b[131])^(a[98] & b[132])^(a[97] & b[133])^(a[96] & b[134])^(a[95] & b[135])^(a[94] & b[136])^(a[93] & b[137])^(a[92] & b[138])^(a[91] & b[139])^(a[90] & b[140])^(a[89] & b[141])^(a[88] & b[142])^(a[87] & b[143])^(a[86] & b[144])^(a[85] & b[145])^(a[84] & b[146])^(a[83] & b[147])^(a[82] & b[148])^(a[81] & b[149])^(a[80] & b[150])^(a[79] & b[151])^(a[78] & b[152])^(a[77] & b[153])^(a[76] & b[154])^(a[75] & b[155])^(a[74] & b[156])^(a[73] & b[157])^(a[72] & b[158])^(a[71] & b[159])^(a[70] & b[160])^(a[69] & b[161])^(a[68] & b[162])^(a[67] & b[163])^(a[66] & b[164])^(a[65] & b[165])^(a[64] & b[166])^(a[63] & b[167])^(a[62] & b[168])^(a[61] & b[169])^(a[60] & b[170])^(a[59] & b[171])^(a[58] & b[172])^(a[57] & b[173])^(a[56] & b[174])^(a[55] & b[175])^(a[54] & b[176])^(a[53] & b[177])^(a[52] & b[178])^(a[51] & b[179])^(a[50] & b[180])^(a[49] & b[181])^(a[48] & b[182])^(a[47] & b[183])^(a[46] & b[184])^(a[45] & b[185])^(a[44] & b[186])^(a[43] & b[187])^(a[42] & b[188])^(a[41] & b[189])^(a[40] & b[190])^(a[39] & b[191])^(a[38] & b[192])^(a[37] & b[193])^(a[36] & b[194])^(a[35] & b[195])^(a[34] & b[196])^(a[33] & b[197])^(a[32] & b[198])^(a[31] & b[199])^(a[30] & b[200])^(a[29] & b[201])^(a[28] & b[202])^(a[27] & b[203])^(a[26] & b[204])^(a[25] & b[205])^(a[24] & b[206])^(a[23] & b[207])^(a[22] & b[208])^(a[21] & b[209])^(a[20] & b[210])^(a[19] & b[211])^(a[18] & b[212])^(a[17] & b[213])^(a[16] & b[214])^(a[15] & b[215])^(a[14] & b[216])^(a[13] & b[217])^(a[12] & b[218])^(a[11] & b[219])^(a[10] & b[220])^(a[9] & b[221])^(a[8] & b[222])^(a[7] & b[223])^(a[6] & b[224])^(a[5] & b[225])^(a[4] & b[226])^(a[3] & b[227])^(a[2] & b[228])^(a[1] & b[229])^(a[0] & b[230]);
assign y[231] = (a[231] & b[0])^(a[230] & b[1])^(a[229] & b[2])^(a[228] & b[3])^(a[227] & b[4])^(a[226] & b[5])^(a[225] & b[6])^(a[224] & b[7])^(a[223] & b[8])^(a[222] & b[9])^(a[221] & b[10])^(a[220] & b[11])^(a[219] & b[12])^(a[218] & b[13])^(a[217] & b[14])^(a[216] & b[15])^(a[215] & b[16])^(a[214] & b[17])^(a[213] & b[18])^(a[212] & b[19])^(a[211] & b[20])^(a[210] & b[21])^(a[209] & b[22])^(a[208] & b[23])^(a[207] & b[24])^(a[206] & b[25])^(a[205] & b[26])^(a[204] & b[27])^(a[203] & b[28])^(a[202] & b[29])^(a[201] & b[30])^(a[200] & b[31])^(a[199] & b[32])^(a[198] & b[33])^(a[197] & b[34])^(a[196] & b[35])^(a[195] & b[36])^(a[194] & b[37])^(a[193] & b[38])^(a[192] & b[39])^(a[191] & b[40])^(a[190] & b[41])^(a[189] & b[42])^(a[188] & b[43])^(a[187] & b[44])^(a[186] & b[45])^(a[185] & b[46])^(a[184] & b[47])^(a[183] & b[48])^(a[182] & b[49])^(a[181] & b[50])^(a[180] & b[51])^(a[179] & b[52])^(a[178] & b[53])^(a[177] & b[54])^(a[176] & b[55])^(a[175] & b[56])^(a[174] & b[57])^(a[173] & b[58])^(a[172] & b[59])^(a[171] & b[60])^(a[170] & b[61])^(a[169] & b[62])^(a[168] & b[63])^(a[167] & b[64])^(a[166] & b[65])^(a[165] & b[66])^(a[164] & b[67])^(a[163] & b[68])^(a[162] & b[69])^(a[161] & b[70])^(a[160] & b[71])^(a[159] & b[72])^(a[158] & b[73])^(a[157] & b[74])^(a[156] & b[75])^(a[155] & b[76])^(a[154] & b[77])^(a[153] & b[78])^(a[152] & b[79])^(a[151] & b[80])^(a[150] & b[81])^(a[149] & b[82])^(a[148] & b[83])^(a[147] & b[84])^(a[146] & b[85])^(a[145] & b[86])^(a[144] & b[87])^(a[143] & b[88])^(a[142] & b[89])^(a[141] & b[90])^(a[140] & b[91])^(a[139] & b[92])^(a[138] & b[93])^(a[137] & b[94])^(a[136] & b[95])^(a[135] & b[96])^(a[134] & b[97])^(a[133] & b[98])^(a[132] & b[99])^(a[131] & b[100])^(a[130] & b[101])^(a[129] & b[102])^(a[128] & b[103])^(a[127] & b[104])^(a[126] & b[105])^(a[125] & b[106])^(a[124] & b[107])^(a[123] & b[108])^(a[122] & b[109])^(a[121] & b[110])^(a[120] & b[111])^(a[119] & b[112])^(a[118] & b[113])^(a[117] & b[114])^(a[116] & b[115])^(a[115] & b[116])^(a[114] & b[117])^(a[113] & b[118])^(a[112] & b[119])^(a[111] & b[120])^(a[110] & b[121])^(a[109] & b[122])^(a[108] & b[123])^(a[107] & b[124])^(a[106] & b[125])^(a[105] & b[126])^(a[104] & b[127])^(a[103] & b[128])^(a[102] & b[129])^(a[101] & b[130])^(a[100] & b[131])^(a[99] & b[132])^(a[98] & b[133])^(a[97] & b[134])^(a[96] & b[135])^(a[95] & b[136])^(a[94] & b[137])^(a[93] & b[138])^(a[92] & b[139])^(a[91] & b[140])^(a[90] & b[141])^(a[89] & b[142])^(a[88] & b[143])^(a[87] & b[144])^(a[86] & b[145])^(a[85] & b[146])^(a[84] & b[147])^(a[83] & b[148])^(a[82] & b[149])^(a[81] & b[150])^(a[80] & b[151])^(a[79] & b[152])^(a[78] & b[153])^(a[77] & b[154])^(a[76] & b[155])^(a[75] & b[156])^(a[74] & b[157])^(a[73] & b[158])^(a[72] & b[159])^(a[71] & b[160])^(a[70] & b[161])^(a[69] & b[162])^(a[68] & b[163])^(a[67] & b[164])^(a[66] & b[165])^(a[65] & b[166])^(a[64] & b[167])^(a[63] & b[168])^(a[62] & b[169])^(a[61] & b[170])^(a[60] & b[171])^(a[59] & b[172])^(a[58] & b[173])^(a[57] & b[174])^(a[56] & b[175])^(a[55] & b[176])^(a[54] & b[177])^(a[53] & b[178])^(a[52] & b[179])^(a[51] & b[180])^(a[50] & b[181])^(a[49] & b[182])^(a[48] & b[183])^(a[47] & b[184])^(a[46] & b[185])^(a[45] & b[186])^(a[44] & b[187])^(a[43] & b[188])^(a[42] & b[189])^(a[41] & b[190])^(a[40] & b[191])^(a[39] & b[192])^(a[38] & b[193])^(a[37] & b[194])^(a[36] & b[195])^(a[35] & b[196])^(a[34] & b[197])^(a[33] & b[198])^(a[32] & b[199])^(a[31] & b[200])^(a[30] & b[201])^(a[29] & b[202])^(a[28] & b[203])^(a[27] & b[204])^(a[26] & b[205])^(a[25] & b[206])^(a[24] & b[207])^(a[23] & b[208])^(a[22] & b[209])^(a[21] & b[210])^(a[20] & b[211])^(a[19] & b[212])^(a[18] & b[213])^(a[17] & b[214])^(a[16] & b[215])^(a[15] & b[216])^(a[14] & b[217])^(a[13] & b[218])^(a[12] & b[219])^(a[11] & b[220])^(a[10] & b[221])^(a[9] & b[222])^(a[8] & b[223])^(a[7] & b[224])^(a[6] & b[225])^(a[5] & b[226])^(a[4] & b[227])^(a[3] & b[228])^(a[2] & b[229])^(a[1] & b[230])^(a[0] & b[231]);
assign y[232] = (a[232] & b[0])^(a[231] & b[1])^(a[230] & b[2])^(a[229] & b[3])^(a[228] & b[4])^(a[227] & b[5])^(a[226] & b[6])^(a[225] & b[7])^(a[224] & b[8])^(a[223] & b[9])^(a[222] & b[10])^(a[221] & b[11])^(a[220] & b[12])^(a[219] & b[13])^(a[218] & b[14])^(a[217] & b[15])^(a[216] & b[16])^(a[215] & b[17])^(a[214] & b[18])^(a[213] & b[19])^(a[212] & b[20])^(a[211] & b[21])^(a[210] & b[22])^(a[209] & b[23])^(a[208] & b[24])^(a[207] & b[25])^(a[206] & b[26])^(a[205] & b[27])^(a[204] & b[28])^(a[203] & b[29])^(a[202] & b[30])^(a[201] & b[31])^(a[200] & b[32])^(a[199] & b[33])^(a[198] & b[34])^(a[197] & b[35])^(a[196] & b[36])^(a[195] & b[37])^(a[194] & b[38])^(a[193] & b[39])^(a[192] & b[40])^(a[191] & b[41])^(a[190] & b[42])^(a[189] & b[43])^(a[188] & b[44])^(a[187] & b[45])^(a[186] & b[46])^(a[185] & b[47])^(a[184] & b[48])^(a[183] & b[49])^(a[182] & b[50])^(a[181] & b[51])^(a[180] & b[52])^(a[179] & b[53])^(a[178] & b[54])^(a[177] & b[55])^(a[176] & b[56])^(a[175] & b[57])^(a[174] & b[58])^(a[173] & b[59])^(a[172] & b[60])^(a[171] & b[61])^(a[170] & b[62])^(a[169] & b[63])^(a[168] & b[64])^(a[167] & b[65])^(a[166] & b[66])^(a[165] & b[67])^(a[164] & b[68])^(a[163] & b[69])^(a[162] & b[70])^(a[161] & b[71])^(a[160] & b[72])^(a[159] & b[73])^(a[158] & b[74])^(a[157] & b[75])^(a[156] & b[76])^(a[155] & b[77])^(a[154] & b[78])^(a[153] & b[79])^(a[152] & b[80])^(a[151] & b[81])^(a[150] & b[82])^(a[149] & b[83])^(a[148] & b[84])^(a[147] & b[85])^(a[146] & b[86])^(a[145] & b[87])^(a[144] & b[88])^(a[143] & b[89])^(a[142] & b[90])^(a[141] & b[91])^(a[140] & b[92])^(a[139] & b[93])^(a[138] & b[94])^(a[137] & b[95])^(a[136] & b[96])^(a[135] & b[97])^(a[134] & b[98])^(a[133] & b[99])^(a[132] & b[100])^(a[131] & b[101])^(a[130] & b[102])^(a[129] & b[103])^(a[128] & b[104])^(a[127] & b[105])^(a[126] & b[106])^(a[125] & b[107])^(a[124] & b[108])^(a[123] & b[109])^(a[122] & b[110])^(a[121] & b[111])^(a[120] & b[112])^(a[119] & b[113])^(a[118] & b[114])^(a[117] & b[115])^(a[116] & b[116])^(a[115] & b[117])^(a[114] & b[118])^(a[113] & b[119])^(a[112] & b[120])^(a[111] & b[121])^(a[110] & b[122])^(a[109] & b[123])^(a[108] & b[124])^(a[107] & b[125])^(a[106] & b[126])^(a[105] & b[127])^(a[104] & b[128])^(a[103] & b[129])^(a[102] & b[130])^(a[101] & b[131])^(a[100] & b[132])^(a[99] & b[133])^(a[98] & b[134])^(a[97] & b[135])^(a[96] & b[136])^(a[95] & b[137])^(a[94] & b[138])^(a[93] & b[139])^(a[92] & b[140])^(a[91] & b[141])^(a[90] & b[142])^(a[89] & b[143])^(a[88] & b[144])^(a[87] & b[145])^(a[86] & b[146])^(a[85] & b[147])^(a[84] & b[148])^(a[83] & b[149])^(a[82] & b[150])^(a[81] & b[151])^(a[80] & b[152])^(a[79] & b[153])^(a[78] & b[154])^(a[77] & b[155])^(a[76] & b[156])^(a[75] & b[157])^(a[74] & b[158])^(a[73] & b[159])^(a[72] & b[160])^(a[71] & b[161])^(a[70] & b[162])^(a[69] & b[163])^(a[68] & b[164])^(a[67] & b[165])^(a[66] & b[166])^(a[65] & b[167])^(a[64] & b[168])^(a[63] & b[169])^(a[62] & b[170])^(a[61] & b[171])^(a[60] & b[172])^(a[59] & b[173])^(a[58] & b[174])^(a[57] & b[175])^(a[56] & b[176])^(a[55] & b[177])^(a[54] & b[178])^(a[53] & b[179])^(a[52] & b[180])^(a[51] & b[181])^(a[50] & b[182])^(a[49] & b[183])^(a[48] & b[184])^(a[47] & b[185])^(a[46] & b[186])^(a[45] & b[187])^(a[44] & b[188])^(a[43] & b[189])^(a[42] & b[190])^(a[41] & b[191])^(a[40] & b[192])^(a[39] & b[193])^(a[38] & b[194])^(a[37] & b[195])^(a[36] & b[196])^(a[35] & b[197])^(a[34] & b[198])^(a[33] & b[199])^(a[32] & b[200])^(a[31] & b[201])^(a[30] & b[202])^(a[29] & b[203])^(a[28] & b[204])^(a[27] & b[205])^(a[26] & b[206])^(a[25] & b[207])^(a[24] & b[208])^(a[23] & b[209])^(a[22] & b[210])^(a[21] & b[211])^(a[20] & b[212])^(a[19] & b[213])^(a[18] & b[214])^(a[17] & b[215])^(a[16] & b[216])^(a[15] & b[217])^(a[14] & b[218])^(a[13] & b[219])^(a[12] & b[220])^(a[11] & b[221])^(a[10] & b[222])^(a[9] & b[223])^(a[8] & b[224])^(a[7] & b[225])^(a[6] & b[226])^(a[5] & b[227])^(a[4] & b[228])^(a[3] & b[229])^(a[2] & b[230])^(a[1] & b[231])^(a[0] & b[232]);
assign y[233] = (a[233] & b[0])^(a[232] & b[1])^(a[231] & b[2])^(a[230] & b[3])^(a[229] & b[4])^(a[228] & b[5])^(a[227] & b[6])^(a[226] & b[7])^(a[225] & b[8])^(a[224] & b[9])^(a[223] & b[10])^(a[222] & b[11])^(a[221] & b[12])^(a[220] & b[13])^(a[219] & b[14])^(a[218] & b[15])^(a[217] & b[16])^(a[216] & b[17])^(a[215] & b[18])^(a[214] & b[19])^(a[213] & b[20])^(a[212] & b[21])^(a[211] & b[22])^(a[210] & b[23])^(a[209] & b[24])^(a[208] & b[25])^(a[207] & b[26])^(a[206] & b[27])^(a[205] & b[28])^(a[204] & b[29])^(a[203] & b[30])^(a[202] & b[31])^(a[201] & b[32])^(a[200] & b[33])^(a[199] & b[34])^(a[198] & b[35])^(a[197] & b[36])^(a[196] & b[37])^(a[195] & b[38])^(a[194] & b[39])^(a[193] & b[40])^(a[192] & b[41])^(a[191] & b[42])^(a[190] & b[43])^(a[189] & b[44])^(a[188] & b[45])^(a[187] & b[46])^(a[186] & b[47])^(a[185] & b[48])^(a[184] & b[49])^(a[183] & b[50])^(a[182] & b[51])^(a[181] & b[52])^(a[180] & b[53])^(a[179] & b[54])^(a[178] & b[55])^(a[177] & b[56])^(a[176] & b[57])^(a[175] & b[58])^(a[174] & b[59])^(a[173] & b[60])^(a[172] & b[61])^(a[171] & b[62])^(a[170] & b[63])^(a[169] & b[64])^(a[168] & b[65])^(a[167] & b[66])^(a[166] & b[67])^(a[165] & b[68])^(a[164] & b[69])^(a[163] & b[70])^(a[162] & b[71])^(a[161] & b[72])^(a[160] & b[73])^(a[159] & b[74])^(a[158] & b[75])^(a[157] & b[76])^(a[156] & b[77])^(a[155] & b[78])^(a[154] & b[79])^(a[153] & b[80])^(a[152] & b[81])^(a[151] & b[82])^(a[150] & b[83])^(a[149] & b[84])^(a[148] & b[85])^(a[147] & b[86])^(a[146] & b[87])^(a[145] & b[88])^(a[144] & b[89])^(a[143] & b[90])^(a[142] & b[91])^(a[141] & b[92])^(a[140] & b[93])^(a[139] & b[94])^(a[138] & b[95])^(a[137] & b[96])^(a[136] & b[97])^(a[135] & b[98])^(a[134] & b[99])^(a[133] & b[100])^(a[132] & b[101])^(a[131] & b[102])^(a[130] & b[103])^(a[129] & b[104])^(a[128] & b[105])^(a[127] & b[106])^(a[126] & b[107])^(a[125] & b[108])^(a[124] & b[109])^(a[123] & b[110])^(a[122] & b[111])^(a[121] & b[112])^(a[120] & b[113])^(a[119] & b[114])^(a[118] & b[115])^(a[117] & b[116])^(a[116] & b[117])^(a[115] & b[118])^(a[114] & b[119])^(a[113] & b[120])^(a[112] & b[121])^(a[111] & b[122])^(a[110] & b[123])^(a[109] & b[124])^(a[108] & b[125])^(a[107] & b[126])^(a[106] & b[127])^(a[105] & b[128])^(a[104] & b[129])^(a[103] & b[130])^(a[102] & b[131])^(a[101] & b[132])^(a[100] & b[133])^(a[99] & b[134])^(a[98] & b[135])^(a[97] & b[136])^(a[96] & b[137])^(a[95] & b[138])^(a[94] & b[139])^(a[93] & b[140])^(a[92] & b[141])^(a[91] & b[142])^(a[90] & b[143])^(a[89] & b[144])^(a[88] & b[145])^(a[87] & b[146])^(a[86] & b[147])^(a[85] & b[148])^(a[84] & b[149])^(a[83] & b[150])^(a[82] & b[151])^(a[81] & b[152])^(a[80] & b[153])^(a[79] & b[154])^(a[78] & b[155])^(a[77] & b[156])^(a[76] & b[157])^(a[75] & b[158])^(a[74] & b[159])^(a[73] & b[160])^(a[72] & b[161])^(a[71] & b[162])^(a[70] & b[163])^(a[69] & b[164])^(a[68] & b[165])^(a[67] & b[166])^(a[66] & b[167])^(a[65] & b[168])^(a[64] & b[169])^(a[63] & b[170])^(a[62] & b[171])^(a[61] & b[172])^(a[60] & b[173])^(a[59] & b[174])^(a[58] & b[175])^(a[57] & b[176])^(a[56] & b[177])^(a[55] & b[178])^(a[54] & b[179])^(a[53] & b[180])^(a[52] & b[181])^(a[51] & b[182])^(a[50] & b[183])^(a[49] & b[184])^(a[48] & b[185])^(a[47] & b[186])^(a[46] & b[187])^(a[45] & b[188])^(a[44] & b[189])^(a[43] & b[190])^(a[42] & b[191])^(a[41] & b[192])^(a[40] & b[193])^(a[39] & b[194])^(a[38] & b[195])^(a[37] & b[196])^(a[36] & b[197])^(a[35] & b[198])^(a[34] & b[199])^(a[33] & b[200])^(a[32] & b[201])^(a[31] & b[202])^(a[30] & b[203])^(a[29] & b[204])^(a[28] & b[205])^(a[27] & b[206])^(a[26] & b[207])^(a[25] & b[208])^(a[24] & b[209])^(a[23] & b[210])^(a[22] & b[211])^(a[21] & b[212])^(a[20] & b[213])^(a[19] & b[214])^(a[18] & b[215])^(a[17] & b[216])^(a[16] & b[217])^(a[15] & b[218])^(a[14] & b[219])^(a[13] & b[220])^(a[12] & b[221])^(a[11] & b[222])^(a[10] & b[223])^(a[9] & b[224])^(a[8] & b[225])^(a[7] & b[226])^(a[6] & b[227])^(a[5] & b[228])^(a[4] & b[229])^(a[3] & b[230])^(a[2] & b[231])^(a[1] & b[232])^(a[0] & b[233]);
assign y[234] = (a[234] & b[0])^(a[233] & b[1])^(a[232] & b[2])^(a[231] & b[3])^(a[230] & b[4])^(a[229] & b[5])^(a[228] & b[6])^(a[227] & b[7])^(a[226] & b[8])^(a[225] & b[9])^(a[224] & b[10])^(a[223] & b[11])^(a[222] & b[12])^(a[221] & b[13])^(a[220] & b[14])^(a[219] & b[15])^(a[218] & b[16])^(a[217] & b[17])^(a[216] & b[18])^(a[215] & b[19])^(a[214] & b[20])^(a[213] & b[21])^(a[212] & b[22])^(a[211] & b[23])^(a[210] & b[24])^(a[209] & b[25])^(a[208] & b[26])^(a[207] & b[27])^(a[206] & b[28])^(a[205] & b[29])^(a[204] & b[30])^(a[203] & b[31])^(a[202] & b[32])^(a[201] & b[33])^(a[200] & b[34])^(a[199] & b[35])^(a[198] & b[36])^(a[197] & b[37])^(a[196] & b[38])^(a[195] & b[39])^(a[194] & b[40])^(a[193] & b[41])^(a[192] & b[42])^(a[191] & b[43])^(a[190] & b[44])^(a[189] & b[45])^(a[188] & b[46])^(a[187] & b[47])^(a[186] & b[48])^(a[185] & b[49])^(a[184] & b[50])^(a[183] & b[51])^(a[182] & b[52])^(a[181] & b[53])^(a[180] & b[54])^(a[179] & b[55])^(a[178] & b[56])^(a[177] & b[57])^(a[176] & b[58])^(a[175] & b[59])^(a[174] & b[60])^(a[173] & b[61])^(a[172] & b[62])^(a[171] & b[63])^(a[170] & b[64])^(a[169] & b[65])^(a[168] & b[66])^(a[167] & b[67])^(a[166] & b[68])^(a[165] & b[69])^(a[164] & b[70])^(a[163] & b[71])^(a[162] & b[72])^(a[161] & b[73])^(a[160] & b[74])^(a[159] & b[75])^(a[158] & b[76])^(a[157] & b[77])^(a[156] & b[78])^(a[155] & b[79])^(a[154] & b[80])^(a[153] & b[81])^(a[152] & b[82])^(a[151] & b[83])^(a[150] & b[84])^(a[149] & b[85])^(a[148] & b[86])^(a[147] & b[87])^(a[146] & b[88])^(a[145] & b[89])^(a[144] & b[90])^(a[143] & b[91])^(a[142] & b[92])^(a[141] & b[93])^(a[140] & b[94])^(a[139] & b[95])^(a[138] & b[96])^(a[137] & b[97])^(a[136] & b[98])^(a[135] & b[99])^(a[134] & b[100])^(a[133] & b[101])^(a[132] & b[102])^(a[131] & b[103])^(a[130] & b[104])^(a[129] & b[105])^(a[128] & b[106])^(a[127] & b[107])^(a[126] & b[108])^(a[125] & b[109])^(a[124] & b[110])^(a[123] & b[111])^(a[122] & b[112])^(a[121] & b[113])^(a[120] & b[114])^(a[119] & b[115])^(a[118] & b[116])^(a[117] & b[117])^(a[116] & b[118])^(a[115] & b[119])^(a[114] & b[120])^(a[113] & b[121])^(a[112] & b[122])^(a[111] & b[123])^(a[110] & b[124])^(a[109] & b[125])^(a[108] & b[126])^(a[107] & b[127])^(a[106] & b[128])^(a[105] & b[129])^(a[104] & b[130])^(a[103] & b[131])^(a[102] & b[132])^(a[101] & b[133])^(a[100] & b[134])^(a[99] & b[135])^(a[98] & b[136])^(a[97] & b[137])^(a[96] & b[138])^(a[95] & b[139])^(a[94] & b[140])^(a[93] & b[141])^(a[92] & b[142])^(a[91] & b[143])^(a[90] & b[144])^(a[89] & b[145])^(a[88] & b[146])^(a[87] & b[147])^(a[86] & b[148])^(a[85] & b[149])^(a[84] & b[150])^(a[83] & b[151])^(a[82] & b[152])^(a[81] & b[153])^(a[80] & b[154])^(a[79] & b[155])^(a[78] & b[156])^(a[77] & b[157])^(a[76] & b[158])^(a[75] & b[159])^(a[74] & b[160])^(a[73] & b[161])^(a[72] & b[162])^(a[71] & b[163])^(a[70] & b[164])^(a[69] & b[165])^(a[68] & b[166])^(a[67] & b[167])^(a[66] & b[168])^(a[65] & b[169])^(a[64] & b[170])^(a[63] & b[171])^(a[62] & b[172])^(a[61] & b[173])^(a[60] & b[174])^(a[59] & b[175])^(a[58] & b[176])^(a[57] & b[177])^(a[56] & b[178])^(a[55] & b[179])^(a[54] & b[180])^(a[53] & b[181])^(a[52] & b[182])^(a[51] & b[183])^(a[50] & b[184])^(a[49] & b[185])^(a[48] & b[186])^(a[47] & b[187])^(a[46] & b[188])^(a[45] & b[189])^(a[44] & b[190])^(a[43] & b[191])^(a[42] & b[192])^(a[41] & b[193])^(a[40] & b[194])^(a[39] & b[195])^(a[38] & b[196])^(a[37] & b[197])^(a[36] & b[198])^(a[35] & b[199])^(a[34] & b[200])^(a[33] & b[201])^(a[32] & b[202])^(a[31] & b[203])^(a[30] & b[204])^(a[29] & b[205])^(a[28] & b[206])^(a[27] & b[207])^(a[26] & b[208])^(a[25] & b[209])^(a[24] & b[210])^(a[23] & b[211])^(a[22] & b[212])^(a[21] & b[213])^(a[20] & b[214])^(a[19] & b[215])^(a[18] & b[216])^(a[17] & b[217])^(a[16] & b[218])^(a[15] & b[219])^(a[14] & b[220])^(a[13] & b[221])^(a[12] & b[222])^(a[11] & b[223])^(a[10] & b[224])^(a[9] & b[225])^(a[8] & b[226])^(a[7] & b[227])^(a[6] & b[228])^(a[5] & b[229])^(a[4] & b[230])^(a[3] & b[231])^(a[2] & b[232])^(a[1] & b[233])^(a[0] & b[234]);
assign y[235] = (a[235] & b[0])^(a[234] & b[1])^(a[233] & b[2])^(a[232] & b[3])^(a[231] & b[4])^(a[230] & b[5])^(a[229] & b[6])^(a[228] & b[7])^(a[227] & b[8])^(a[226] & b[9])^(a[225] & b[10])^(a[224] & b[11])^(a[223] & b[12])^(a[222] & b[13])^(a[221] & b[14])^(a[220] & b[15])^(a[219] & b[16])^(a[218] & b[17])^(a[217] & b[18])^(a[216] & b[19])^(a[215] & b[20])^(a[214] & b[21])^(a[213] & b[22])^(a[212] & b[23])^(a[211] & b[24])^(a[210] & b[25])^(a[209] & b[26])^(a[208] & b[27])^(a[207] & b[28])^(a[206] & b[29])^(a[205] & b[30])^(a[204] & b[31])^(a[203] & b[32])^(a[202] & b[33])^(a[201] & b[34])^(a[200] & b[35])^(a[199] & b[36])^(a[198] & b[37])^(a[197] & b[38])^(a[196] & b[39])^(a[195] & b[40])^(a[194] & b[41])^(a[193] & b[42])^(a[192] & b[43])^(a[191] & b[44])^(a[190] & b[45])^(a[189] & b[46])^(a[188] & b[47])^(a[187] & b[48])^(a[186] & b[49])^(a[185] & b[50])^(a[184] & b[51])^(a[183] & b[52])^(a[182] & b[53])^(a[181] & b[54])^(a[180] & b[55])^(a[179] & b[56])^(a[178] & b[57])^(a[177] & b[58])^(a[176] & b[59])^(a[175] & b[60])^(a[174] & b[61])^(a[173] & b[62])^(a[172] & b[63])^(a[171] & b[64])^(a[170] & b[65])^(a[169] & b[66])^(a[168] & b[67])^(a[167] & b[68])^(a[166] & b[69])^(a[165] & b[70])^(a[164] & b[71])^(a[163] & b[72])^(a[162] & b[73])^(a[161] & b[74])^(a[160] & b[75])^(a[159] & b[76])^(a[158] & b[77])^(a[157] & b[78])^(a[156] & b[79])^(a[155] & b[80])^(a[154] & b[81])^(a[153] & b[82])^(a[152] & b[83])^(a[151] & b[84])^(a[150] & b[85])^(a[149] & b[86])^(a[148] & b[87])^(a[147] & b[88])^(a[146] & b[89])^(a[145] & b[90])^(a[144] & b[91])^(a[143] & b[92])^(a[142] & b[93])^(a[141] & b[94])^(a[140] & b[95])^(a[139] & b[96])^(a[138] & b[97])^(a[137] & b[98])^(a[136] & b[99])^(a[135] & b[100])^(a[134] & b[101])^(a[133] & b[102])^(a[132] & b[103])^(a[131] & b[104])^(a[130] & b[105])^(a[129] & b[106])^(a[128] & b[107])^(a[127] & b[108])^(a[126] & b[109])^(a[125] & b[110])^(a[124] & b[111])^(a[123] & b[112])^(a[122] & b[113])^(a[121] & b[114])^(a[120] & b[115])^(a[119] & b[116])^(a[118] & b[117])^(a[117] & b[118])^(a[116] & b[119])^(a[115] & b[120])^(a[114] & b[121])^(a[113] & b[122])^(a[112] & b[123])^(a[111] & b[124])^(a[110] & b[125])^(a[109] & b[126])^(a[108] & b[127])^(a[107] & b[128])^(a[106] & b[129])^(a[105] & b[130])^(a[104] & b[131])^(a[103] & b[132])^(a[102] & b[133])^(a[101] & b[134])^(a[100] & b[135])^(a[99] & b[136])^(a[98] & b[137])^(a[97] & b[138])^(a[96] & b[139])^(a[95] & b[140])^(a[94] & b[141])^(a[93] & b[142])^(a[92] & b[143])^(a[91] & b[144])^(a[90] & b[145])^(a[89] & b[146])^(a[88] & b[147])^(a[87] & b[148])^(a[86] & b[149])^(a[85] & b[150])^(a[84] & b[151])^(a[83] & b[152])^(a[82] & b[153])^(a[81] & b[154])^(a[80] & b[155])^(a[79] & b[156])^(a[78] & b[157])^(a[77] & b[158])^(a[76] & b[159])^(a[75] & b[160])^(a[74] & b[161])^(a[73] & b[162])^(a[72] & b[163])^(a[71] & b[164])^(a[70] & b[165])^(a[69] & b[166])^(a[68] & b[167])^(a[67] & b[168])^(a[66] & b[169])^(a[65] & b[170])^(a[64] & b[171])^(a[63] & b[172])^(a[62] & b[173])^(a[61] & b[174])^(a[60] & b[175])^(a[59] & b[176])^(a[58] & b[177])^(a[57] & b[178])^(a[56] & b[179])^(a[55] & b[180])^(a[54] & b[181])^(a[53] & b[182])^(a[52] & b[183])^(a[51] & b[184])^(a[50] & b[185])^(a[49] & b[186])^(a[48] & b[187])^(a[47] & b[188])^(a[46] & b[189])^(a[45] & b[190])^(a[44] & b[191])^(a[43] & b[192])^(a[42] & b[193])^(a[41] & b[194])^(a[40] & b[195])^(a[39] & b[196])^(a[38] & b[197])^(a[37] & b[198])^(a[36] & b[199])^(a[35] & b[200])^(a[34] & b[201])^(a[33] & b[202])^(a[32] & b[203])^(a[31] & b[204])^(a[30] & b[205])^(a[29] & b[206])^(a[28] & b[207])^(a[27] & b[208])^(a[26] & b[209])^(a[25] & b[210])^(a[24] & b[211])^(a[23] & b[212])^(a[22] & b[213])^(a[21] & b[214])^(a[20] & b[215])^(a[19] & b[216])^(a[18] & b[217])^(a[17] & b[218])^(a[16] & b[219])^(a[15] & b[220])^(a[14] & b[221])^(a[13] & b[222])^(a[12] & b[223])^(a[11] & b[224])^(a[10] & b[225])^(a[9] & b[226])^(a[8] & b[227])^(a[7] & b[228])^(a[6] & b[229])^(a[5] & b[230])^(a[4] & b[231])^(a[3] & b[232])^(a[2] & b[233])^(a[1] & b[234])^(a[0] & b[235]);
assign y[236] = (a[236] & b[0])^(a[235] & b[1])^(a[234] & b[2])^(a[233] & b[3])^(a[232] & b[4])^(a[231] & b[5])^(a[230] & b[6])^(a[229] & b[7])^(a[228] & b[8])^(a[227] & b[9])^(a[226] & b[10])^(a[225] & b[11])^(a[224] & b[12])^(a[223] & b[13])^(a[222] & b[14])^(a[221] & b[15])^(a[220] & b[16])^(a[219] & b[17])^(a[218] & b[18])^(a[217] & b[19])^(a[216] & b[20])^(a[215] & b[21])^(a[214] & b[22])^(a[213] & b[23])^(a[212] & b[24])^(a[211] & b[25])^(a[210] & b[26])^(a[209] & b[27])^(a[208] & b[28])^(a[207] & b[29])^(a[206] & b[30])^(a[205] & b[31])^(a[204] & b[32])^(a[203] & b[33])^(a[202] & b[34])^(a[201] & b[35])^(a[200] & b[36])^(a[199] & b[37])^(a[198] & b[38])^(a[197] & b[39])^(a[196] & b[40])^(a[195] & b[41])^(a[194] & b[42])^(a[193] & b[43])^(a[192] & b[44])^(a[191] & b[45])^(a[190] & b[46])^(a[189] & b[47])^(a[188] & b[48])^(a[187] & b[49])^(a[186] & b[50])^(a[185] & b[51])^(a[184] & b[52])^(a[183] & b[53])^(a[182] & b[54])^(a[181] & b[55])^(a[180] & b[56])^(a[179] & b[57])^(a[178] & b[58])^(a[177] & b[59])^(a[176] & b[60])^(a[175] & b[61])^(a[174] & b[62])^(a[173] & b[63])^(a[172] & b[64])^(a[171] & b[65])^(a[170] & b[66])^(a[169] & b[67])^(a[168] & b[68])^(a[167] & b[69])^(a[166] & b[70])^(a[165] & b[71])^(a[164] & b[72])^(a[163] & b[73])^(a[162] & b[74])^(a[161] & b[75])^(a[160] & b[76])^(a[159] & b[77])^(a[158] & b[78])^(a[157] & b[79])^(a[156] & b[80])^(a[155] & b[81])^(a[154] & b[82])^(a[153] & b[83])^(a[152] & b[84])^(a[151] & b[85])^(a[150] & b[86])^(a[149] & b[87])^(a[148] & b[88])^(a[147] & b[89])^(a[146] & b[90])^(a[145] & b[91])^(a[144] & b[92])^(a[143] & b[93])^(a[142] & b[94])^(a[141] & b[95])^(a[140] & b[96])^(a[139] & b[97])^(a[138] & b[98])^(a[137] & b[99])^(a[136] & b[100])^(a[135] & b[101])^(a[134] & b[102])^(a[133] & b[103])^(a[132] & b[104])^(a[131] & b[105])^(a[130] & b[106])^(a[129] & b[107])^(a[128] & b[108])^(a[127] & b[109])^(a[126] & b[110])^(a[125] & b[111])^(a[124] & b[112])^(a[123] & b[113])^(a[122] & b[114])^(a[121] & b[115])^(a[120] & b[116])^(a[119] & b[117])^(a[118] & b[118])^(a[117] & b[119])^(a[116] & b[120])^(a[115] & b[121])^(a[114] & b[122])^(a[113] & b[123])^(a[112] & b[124])^(a[111] & b[125])^(a[110] & b[126])^(a[109] & b[127])^(a[108] & b[128])^(a[107] & b[129])^(a[106] & b[130])^(a[105] & b[131])^(a[104] & b[132])^(a[103] & b[133])^(a[102] & b[134])^(a[101] & b[135])^(a[100] & b[136])^(a[99] & b[137])^(a[98] & b[138])^(a[97] & b[139])^(a[96] & b[140])^(a[95] & b[141])^(a[94] & b[142])^(a[93] & b[143])^(a[92] & b[144])^(a[91] & b[145])^(a[90] & b[146])^(a[89] & b[147])^(a[88] & b[148])^(a[87] & b[149])^(a[86] & b[150])^(a[85] & b[151])^(a[84] & b[152])^(a[83] & b[153])^(a[82] & b[154])^(a[81] & b[155])^(a[80] & b[156])^(a[79] & b[157])^(a[78] & b[158])^(a[77] & b[159])^(a[76] & b[160])^(a[75] & b[161])^(a[74] & b[162])^(a[73] & b[163])^(a[72] & b[164])^(a[71] & b[165])^(a[70] & b[166])^(a[69] & b[167])^(a[68] & b[168])^(a[67] & b[169])^(a[66] & b[170])^(a[65] & b[171])^(a[64] & b[172])^(a[63] & b[173])^(a[62] & b[174])^(a[61] & b[175])^(a[60] & b[176])^(a[59] & b[177])^(a[58] & b[178])^(a[57] & b[179])^(a[56] & b[180])^(a[55] & b[181])^(a[54] & b[182])^(a[53] & b[183])^(a[52] & b[184])^(a[51] & b[185])^(a[50] & b[186])^(a[49] & b[187])^(a[48] & b[188])^(a[47] & b[189])^(a[46] & b[190])^(a[45] & b[191])^(a[44] & b[192])^(a[43] & b[193])^(a[42] & b[194])^(a[41] & b[195])^(a[40] & b[196])^(a[39] & b[197])^(a[38] & b[198])^(a[37] & b[199])^(a[36] & b[200])^(a[35] & b[201])^(a[34] & b[202])^(a[33] & b[203])^(a[32] & b[204])^(a[31] & b[205])^(a[30] & b[206])^(a[29] & b[207])^(a[28] & b[208])^(a[27] & b[209])^(a[26] & b[210])^(a[25] & b[211])^(a[24] & b[212])^(a[23] & b[213])^(a[22] & b[214])^(a[21] & b[215])^(a[20] & b[216])^(a[19] & b[217])^(a[18] & b[218])^(a[17] & b[219])^(a[16] & b[220])^(a[15] & b[221])^(a[14] & b[222])^(a[13] & b[223])^(a[12] & b[224])^(a[11] & b[225])^(a[10] & b[226])^(a[9] & b[227])^(a[8] & b[228])^(a[7] & b[229])^(a[6] & b[230])^(a[5] & b[231])^(a[4] & b[232])^(a[3] & b[233])^(a[2] & b[234])^(a[1] & b[235])^(a[0] & b[236]);
assign y[237] = (a[237] & b[0])^(a[236] & b[1])^(a[235] & b[2])^(a[234] & b[3])^(a[233] & b[4])^(a[232] & b[5])^(a[231] & b[6])^(a[230] & b[7])^(a[229] & b[8])^(a[228] & b[9])^(a[227] & b[10])^(a[226] & b[11])^(a[225] & b[12])^(a[224] & b[13])^(a[223] & b[14])^(a[222] & b[15])^(a[221] & b[16])^(a[220] & b[17])^(a[219] & b[18])^(a[218] & b[19])^(a[217] & b[20])^(a[216] & b[21])^(a[215] & b[22])^(a[214] & b[23])^(a[213] & b[24])^(a[212] & b[25])^(a[211] & b[26])^(a[210] & b[27])^(a[209] & b[28])^(a[208] & b[29])^(a[207] & b[30])^(a[206] & b[31])^(a[205] & b[32])^(a[204] & b[33])^(a[203] & b[34])^(a[202] & b[35])^(a[201] & b[36])^(a[200] & b[37])^(a[199] & b[38])^(a[198] & b[39])^(a[197] & b[40])^(a[196] & b[41])^(a[195] & b[42])^(a[194] & b[43])^(a[193] & b[44])^(a[192] & b[45])^(a[191] & b[46])^(a[190] & b[47])^(a[189] & b[48])^(a[188] & b[49])^(a[187] & b[50])^(a[186] & b[51])^(a[185] & b[52])^(a[184] & b[53])^(a[183] & b[54])^(a[182] & b[55])^(a[181] & b[56])^(a[180] & b[57])^(a[179] & b[58])^(a[178] & b[59])^(a[177] & b[60])^(a[176] & b[61])^(a[175] & b[62])^(a[174] & b[63])^(a[173] & b[64])^(a[172] & b[65])^(a[171] & b[66])^(a[170] & b[67])^(a[169] & b[68])^(a[168] & b[69])^(a[167] & b[70])^(a[166] & b[71])^(a[165] & b[72])^(a[164] & b[73])^(a[163] & b[74])^(a[162] & b[75])^(a[161] & b[76])^(a[160] & b[77])^(a[159] & b[78])^(a[158] & b[79])^(a[157] & b[80])^(a[156] & b[81])^(a[155] & b[82])^(a[154] & b[83])^(a[153] & b[84])^(a[152] & b[85])^(a[151] & b[86])^(a[150] & b[87])^(a[149] & b[88])^(a[148] & b[89])^(a[147] & b[90])^(a[146] & b[91])^(a[145] & b[92])^(a[144] & b[93])^(a[143] & b[94])^(a[142] & b[95])^(a[141] & b[96])^(a[140] & b[97])^(a[139] & b[98])^(a[138] & b[99])^(a[137] & b[100])^(a[136] & b[101])^(a[135] & b[102])^(a[134] & b[103])^(a[133] & b[104])^(a[132] & b[105])^(a[131] & b[106])^(a[130] & b[107])^(a[129] & b[108])^(a[128] & b[109])^(a[127] & b[110])^(a[126] & b[111])^(a[125] & b[112])^(a[124] & b[113])^(a[123] & b[114])^(a[122] & b[115])^(a[121] & b[116])^(a[120] & b[117])^(a[119] & b[118])^(a[118] & b[119])^(a[117] & b[120])^(a[116] & b[121])^(a[115] & b[122])^(a[114] & b[123])^(a[113] & b[124])^(a[112] & b[125])^(a[111] & b[126])^(a[110] & b[127])^(a[109] & b[128])^(a[108] & b[129])^(a[107] & b[130])^(a[106] & b[131])^(a[105] & b[132])^(a[104] & b[133])^(a[103] & b[134])^(a[102] & b[135])^(a[101] & b[136])^(a[100] & b[137])^(a[99] & b[138])^(a[98] & b[139])^(a[97] & b[140])^(a[96] & b[141])^(a[95] & b[142])^(a[94] & b[143])^(a[93] & b[144])^(a[92] & b[145])^(a[91] & b[146])^(a[90] & b[147])^(a[89] & b[148])^(a[88] & b[149])^(a[87] & b[150])^(a[86] & b[151])^(a[85] & b[152])^(a[84] & b[153])^(a[83] & b[154])^(a[82] & b[155])^(a[81] & b[156])^(a[80] & b[157])^(a[79] & b[158])^(a[78] & b[159])^(a[77] & b[160])^(a[76] & b[161])^(a[75] & b[162])^(a[74] & b[163])^(a[73] & b[164])^(a[72] & b[165])^(a[71] & b[166])^(a[70] & b[167])^(a[69] & b[168])^(a[68] & b[169])^(a[67] & b[170])^(a[66] & b[171])^(a[65] & b[172])^(a[64] & b[173])^(a[63] & b[174])^(a[62] & b[175])^(a[61] & b[176])^(a[60] & b[177])^(a[59] & b[178])^(a[58] & b[179])^(a[57] & b[180])^(a[56] & b[181])^(a[55] & b[182])^(a[54] & b[183])^(a[53] & b[184])^(a[52] & b[185])^(a[51] & b[186])^(a[50] & b[187])^(a[49] & b[188])^(a[48] & b[189])^(a[47] & b[190])^(a[46] & b[191])^(a[45] & b[192])^(a[44] & b[193])^(a[43] & b[194])^(a[42] & b[195])^(a[41] & b[196])^(a[40] & b[197])^(a[39] & b[198])^(a[38] & b[199])^(a[37] & b[200])^(a[36] & b[201])^(a[35] & b[202])^(a[34] & b[203])^(a[33] & b[204])^(a[32] & b[205])^(a[31] & b[206])^(a[30] & b[207])^(a[29] & b[208])^(a[28] & b[209])^(a[27] & b[210])^(a[26] & b[211])^(a[25] & b[212])^(a[24] & b[213])^(a[23] & b[214])^(a[22] & b[215])^(a[21] & b[216])^(a[20] & b[217])^(a[19] & b[218])^(a[18] & b[219])^(a[17] & b[220])^(a[16] & b[221])^(a[15] & b[222])^(a[14] & b[223])^(a[13] & b[224])^(a[12] & b[225])^(a[11] & b[226])^(a[10] & b[227])^(a[9] & b[228])^(a[8] & b[229])^(a[7] & b[230])^(a[6] & b[231])^(a[5] & b[232])^(a[4] & b[233])^(a[3] & b[234])^(a[2] & b[235])^(a[1] & b[236])^(a[0] & b[237]);
assign y[238] = (a[238] & b[0])^(a[237] & b[1])^(a[236] & b[2])^(a[235] & b[3])^(a[234] & b[4])^(a[233] & b[5])^(a[232] & b[6])^(a[231] & b[7])^(a[230] & b[8])^(a[229] & b[9])^(a[228] & b[10])^(a[227] & b[11])^(a[226] & b[12])^(a[225] & b[13])^(a[224] & b[14])^(a[223] & b[15])^(a[222] & b[16])^(a[221] & b[17])^(a[220] & b[18])^(a[219] & b[19])^(a[218] & b[20])^(a[217] & b[21])^(a[216] & b[22])^(a[215] & b[23])^(a[214] & b[24])^(a[213] & b[25])^(a[212] & b[26])^(a[211] & b[27])^(a[210] & b[28])^(a[209] & b[29])^(a[208] & b[30])^(a[207] & b[31])^(a[206] & b[32])^(a[205] & b[33])^(a[204] & b[34])^(a[203] & b[35])^(a[202] & b[36])^(a[201] & b[37])^(a[200] & b[38])^(a[199] & b[39])^(a[198] & b[40])^(a[197] & b[41])^(a[196] & b[42])^(a[195] & b[43])^(a[194] & b[44])^(a[193] & b[45])^(a[192] & b[46])^(a[191] & b[47])^(a[190] & b[48])^(a[189] & b[49])^(a[188] & b[50])^(a[187] & b[51])^(a[186] & b[52])^(a[185] & b[53])^(a[184] & b[54])^(a[183] & b[55])^(a[182] & b[56])^(a[181] & b[57])^(a[180] & b[58])^(a[179] & b[59])^(a[178] & b[60])^(a[177] & b[61])^(a[176] & b[62])^(a[175] & b[63])^(a[174] & b[64])^(a[173] & b[65])^(a[172] & b[66])^(a[171] & b[67])^(a[170] & b[68])^(a[169] & b[69])^(a[168] & b[70])^(a[167] & b[71])^(a[166] & b[72])^(a[165] & b[73])^(a[164] & b[74])^(a[163] & b[75])^(a[162] & b[76])^(a[161] & b[77])^(a[160] & b[78])^(a[159] & b[79])^(a[158] & b[80])^(a[157] & b[81])^(a[156] & b[82])^(a[155] & b[83])^(a[154] & b[84])^(a[153] & b[85])^(a[152] & b[86])^(a[151] & b[87])^(a[150] & b[88])^(a[149] & b[89])^(a[148] & b[90])^(a[147] & b[91])^(a[146] & b[92])^(a[145] & b[93])^(a[144] & b[94])^(a[143] & b[95])^(a[142] & b[96])^(a[141] & b[97])^(a[140] & b[98])^(a[139] & b[99])^(a[138] & b[100])^(a[137] & b[101])^(a[136] & b[102])^(a[135] & b[103])^(a[134] & b[104])^(a[133] & b[105])^(a[132] & b[106])^(a[131] & b[107])^(a[130] & b[108])^(a[129] & b[109])^(a[128] & b[110])^(a[127] & b[111])^(a[126] & b[112])^(a[125] & b[113])^(a[124] & b[114])^(a[123] & b[115])^(a[122] & b[116])^(a[121] & b[117])^(a[120] & b[118])^(a[119] & b[119])^(a[118] & b[120])^(a[117] & b[121])^(a[116] & b[122])^(a[115] & b[123])^(a[114] & b[124])^(a[113] & b[125])^(a[112] & b[126])^(a[111] & b[127])^(a[110] & b[128])^(a[109] & b[129])^(a[108] & b[130])^(a[107] & b[131])^(a[106] & b[132])^(a[105] & b[133])^(a[104] & b[134])^(a[103] & b[135])^(a[102] & b[136])^(a[101] & b[137])^(a[100] & b[138])^(a[99] & b[139])^(a[98] & b[140])^(a[97] & b[141])^(a[96] & b[142])^(a[95] & b[143])^(a[94] & b[144])^(a[93] & b[145])^(a[92] & b[146])^(a[91] & b[147])^(a[90] & b[148])^(a[89] & b[149])^(a[88] & b[150])^(a[87] & b[151])^(a[86] & b[152])^(a[85] & b[153])^(a[84] & b[154])^(a[83] & b[155])^(a[82] & b[156])^(a[81] & b[157])^(a[80] & b[158])^(a[79] & b[159])^(a[78] & b[160])^(a[77] & b[161])^(a[76] & b[162])^(a[75] & b[163])^(a[74] & b[164])^(a[73] & b[165])^(a[72] & b[166])^(a[71] & b[167])^(a[70] & b[168])^(a[69] & b[169])^(a[68] & b[170])^(a[67] & b[171])^(a[66] & b[172])^(a[65] & b[173])^(a[64] & b[174])^(a[63] & b[175])^(a[62] & b[176])^(a[61] & b[177])^(a[60] & b[178])^(a[59] & b[179])^(a[58] & b[180])^(a[57] & b[181])^(a[56] & b[182])^(a[55] & b[183])^(a[54] & b[184])^(a[53] & b[185])^(a[52] & b[186])^(a[51] & b[187])^(a[50] & b[188])^(a[49] & b[189])^(a[48] & b[190])^(a[47] & b[191])^(a[46] & b[192])^(a[45] & b[193])^(a[44] & b[194])^(a[43] & b[195])^(a[42] & b[196])^(a[41] & b[197])^(a[40] & b[198])^(a[39] & b[199])^(a[38] & b[200])^(a[37] & b[201])^(a[36] & b[202])^(a[35] & b[203])^(a[34] & b[204])^(a[33] & b[205])^(a[32] & b[206])^(a[31] & b[207])^(a[30] & b[208])^(a[29] & b[209])^(a[28] & b[210])^(a[27] & b[211])^(a[26] & b[212])^(a[25] & b[213])^(a[24] & b[214])^(a[23] & b[215])^(a[22] & b[216])^(a[21] & b[217])^(a[20] & b[218])^(a[19] & b[219])^(a[18] & b[220])^(a[17] & b[221])^(a[16] & b[222])^(a[15] & b[223])^(a[14] & b[224])^(a[13] & b[225])^(a[12] & b[226])^(a[11] & b[227])^(a[10] & b[228])^(a[9] & b[229])^(a[8] & b[230])^(a[7] & b[231])^(a[6] & b[232])^(a[5] & b[233])^(a[4] & b[234])^(a[3] & b[235])^(a[2] & b[236])^(a[1] & b[237])^(a[0] & b[238]);
assign y[239] = (a[239] & b[0])^(a[238] & b[1])^(a[237] & b[2])^(a[236] & b[3])^(a[235] & b[4])^(a[234] & b[5])^(a[233] & b[6])^(a[232] & b[7])^(a[231] & b[8])^(a[230] & b[9])^(a[229] & b[10])^(a[228] & b[11])^(a[227] & b[12])^(a[226] & b[13])^(a[225] & b[14])^(a[224] & b[15])^(a[223] & b[16])^(a[222] & b[17])^(a[221] & b[18])^(a[220] & b[19])^(a[219] & b[20])^(a[218] & b[21])^(a[217] & b[22])^(a[216] & b[23])^(a[215] & b[24])^(a[214] & b[25])^(a[213] & b[26])^(a[212] & b[27])^(a[211] & b[28])^(a[210] & b[29])^(a[209] & b[30])^(a[208] & b[31])^(a[207] & b[32])^(a[206] & b[33])^(a[205] & b[34])^(a[204] & b[35])^(a[203] & b[36])^(a[202] & b[37])^(a[201] & b[38])^(a[200] & b[39])^(a[199] & b[40])^(a[198] & b[41])^(a[197] & b[42])^(a[196] & b[43])^(a[195] & b[44])^(a[194] & b[45])^(a[193] & b[46])^(a[192] & b[47])^(a[191] & b[48])^(a[190] & b[49])^(a[189] & b[50])^(a[188] & b[51])^(a[187] & b[52])^(a[186] & b[53])^(a[185] & b[54])^(a[184] & b[55])^(a[183] & b[56])^(a[182] & b[57])^(a[181] & b[58])^(a[180] & b[59])^(a[179] & b[60])^(a[178] & b[61])^(a[177] & b[62])^(a[176] & b[63])^(a[175] & b[64])^(a[174] & b[65])^(a[173] & b[66])^(a[172] & b[67])^(a[171] & b[68])^(a[170] & b[69])^(a[169] & b[70])^(a[168] & b[71])^(a[167] & b[72])^(a[166] & b[73])^(a[165] & b[74])^(a[164] & b[75])^(a[163] & b[76])^(a[162] & b[77])^(a[161] & b[78])^(a[160] & b[79])^(a[159] & b[80])^(a[158] & b[81])^(a[157] & b[82])^(a[156] & b[83])^(a[155] & b[84])^(a[154] & b[85])^(a[153] & b[86])^(a[152] & b[87])^(a[151] & b[88])^(a[150] & b[89])^(a[149] & b[90])^(a[148] & b[91])^(a[147] & b[92])^(a[146] & b[93])^(a[145] & b[94])^(a[144] & b[95])^(a[143] & b[96])^(a[142] & b[97])^(a[141] & b[98])^(a[140] & b[99])^(a[139] & b[100])^(a[138] & b[101])^(a[137] & b[102])^(a[136] & b[103])^(a[135] & b[104])^(a[134] & b[105])^(a[133] & b[106])^(a[132] & b[107])^(a[131] & b[108])^(a[130] & b[109])^(a[129] & b[110])^(a[128] & b[111])^(a[127] & b[112])^(a[126] & b[113])^(a[125] & b[114])^(a[124] & b[115])^(a[123] & b[116])^(a[122] & b[117])^(a[121] & b[118])^(a[120] & b[119])^(a[119] & b[120])^(a[118] & b[121])^(a[117] & b[122])^(a[116] & b[123])^(a[115] & b[124])^(a[114] & b[125])^(a[113] & b[126])^(a[112] & b[127])^(a[111] & b[128])^(a[110] & b[129])^(a[109] & b[130])^(a[108] & b[131])^(a[107] & b[132])^(a[106] & b[133])^(a[105] & b[134])^(a[104] & b[135])^(a[103] & b[136])^(a[102] & b[137])^(a[101] & b[138])^(a[100] & b[139])^(a[99] & b[140])^(a[98] & b[141])^(a[97] & b[142])^(a[96] & b[143])^(a[95] & b[144])^(a[94] & b[145])^(a[93] & b[146])^(a[92] & b[147])^(a[91] & b[148])^(a[90] & b[149])^(a[89] & b[150])^(a[88] & b[151])^(a[87] & b[152])^(a[86] & b[153])^(a[85] & b[154])^(a[84] & b[155])^(a[83] & b[156])^(a[82] & b[157])^(a[81] & b[158])^(a[80] & b[159])^(a[79] & b[160])^(a[78] & b[161])^(a[77] & b[162])^(a[76] & b[163])^(a[75] & b[164])^(a[74] & b[165])^(a[73] & b[166])^(a[72] & b[167])^(a[71] & b[168])^(a[70] & b[169])^(a[69] & b[170])^(a[68] & b[171])^(a[67] & b[172])^(a[66] & b[173])^(a[65] & b[174])^(a[64] & b[175])^(a[63] & b[176])^(a[62] & b[177])^(a[61] & b[178])^(a[60] & b[179])^(a[59] & b[180])^(a[58] & b[181])^(a[57] & b[182])^(a[56] & b[183])^(a[55] & b[184])^(a[54] & b[185])^(a[53] & b[186])^(a[52] & b[187])^(a[51] & b[188])^(a[50] & b[189])^(a[49] & b[190])^(a[48] & b[191])^(a[47] & b[192])^(a[46] & b[193])^(a[45] & b[194])^(a[44] & b[195])^(a[43] & b[196])^(a[42] & b[197])^(a[41] & b[198])^(a[40] & b[199])^(a[39] & b[200])^(a[38] & b[201])^(a[37] & b[202])^(a[36] & b[203])^(a[35] & b[204])^(a[34] & b[205])^(a[33] & b[206])^(a[32] & b[207])^(a[31] & b[208])^(a[30] & b[209])^(a[29] & b[210])^(a[28] & b[211])^(a[27] & b[212])^(a[26] & b[213])^(a[25] & b[214])^(a[24] & b[215])^(a[23] & b[216])^(a[22] & b[217])^(a[21] & b[218])^(a[20] & b[219])^(a[19] & b[220])^(a[18] & b[221])^(a[17] & b[222])^(a[16] & b[223])^(a[15] & b[224])^(a[14] & b[225])^(a[13] & b[226])^(a[12] & b[227])^(a[11] & b[228])^(a[10] & b[229])^(a[9] & b[230])^(a[8] & b[231])^(a[7] & b[232])^(a[6] & b[233])^(a[5] & b[234])^(a[4] & b[235])^(a[3] & b[236])^(a[2] & b[237])^(a[1] & b[238])^(a[0] & b[239]);
assign y[240] = (a[240] & b[0])^(a[239] & b[1])^(a[238] & b[2])^(a[237] & b[3])^(a[236] & b[4])^(a[235] & b[5])^(a[234] & b[6])^(a[233] & b[7])^(a[232] & b[8])^(a[231] & b[9])^(a[230] & b[10])^(a[229] & b[11])^(a[228] & b[12])^(a[227] & b[13])^(a[226] & b[14])^(a[225] & b[15])^(a[224] & b[16])^(a[223] & b[17])^(a[222] & b[18])^(a[221] & b[19])^(a[220] & b[20])^(a[219] & b[21])^(a[218] & b[22])^(a[217] & b[23])^(a[216] & b[24])^(a[215] & b[25])^(a[214] & b[26])^(a[213] & b[27])^(a[212] & b[28])^(a[211] & b[29])^(a[210] & b[30])^(a[209] & b[31])^(a[208] & b[32])^(a[207] & b[33])^(a[206] & b[34])^(a[205] & b[35])^(a[204] & b[36])^(a[203] & b[37])^(a[202] & b[38])^(a[201] & b[39])^(a[200] & b[40])^(a[199] & b[41])^(a[198] & b[42])^(a[197] & b[43])^(a[196] & b[44])^(a[195] & b[45])^(a[194] & b[46])^(a[193] & b[47])^(a[192] & b[48])^(a[191] & b[49])^(a[190] & b[50])^(a[189] & b[51])^(a[188] & b[52])^(a[187] & b[53])^(a[186] & b[54])^(a[185] & b[55])^(a[184] & b[56])^(a[183] & b[57])^(a[182] & b[58])^(a[181] & b[59])^(a[180] & b[60])^(a[179] & b[61])^(a[178] & b[62])^(a[177] & b[63])^(a[176] & b[64])^(a[175] & b[65])^(a[174] & b[66])^(a[173] & b[67])^(a[172] & b[68])^(a[171] & b[69])^(a[170] & b[70])^(a[169] & b[71])^(a[168] & b[72])^(a[167] & b[73])^(a[166] & b[74])^(a[165] & b[75])^(a[164] & b[76])^(a[163] & b[77])^(a[162] & b[78])^(a[161] & b[79])^(a[160] & b[80])^(a[159] & b[81])^(a[158] & b[82])^(a[157] & b[83])^(a[156] & b[84])^(a[155] & b[85])^(a[154] & b[86])^(a[153] & b[87])^(a[152] & b[88])^(a[151] & b[89])^(a[150] & b[90])^(a[149] & b[91])^(a[148] & b[92])^(a[147] & b[93])^(a[146] & b[94])^(a[145] & b[95])^(a[144] & b[96])^(a[143] & b[97])^(a[142] & b[98])^(a[141] & b[99])^(a[140] & b[100])^(a[139] & b[101])^(a[138] & b[102])^(a[137] & b[103])^(a[136] & b[104])^(a[135] & b[105])^(a[134] & b[106])^(a[133] & b[107])^(a[132] & b[108])^(a[131] & b[109])^(a[130] & b[110])^(a[129] & b[111])^(a[128] & b[112])^(a[127] & b[113])^(a[126] & b[114])^(a[125] & b[115])^(a[124] & b[116])^(a[123] & b[117])^(a[122] & b[118])^(a[121] & b[119])^(a[120] & b[120])^(a[119] & b[121])^(a[118] & b[122])^(a[117] & b[123])^(a[116] & b[124])^(a[115] & b[125])^(a[114] & b[126])^(a[113] & b[127])^(a[112] & b[128])^(a[111] & b[129])^(a[110] & b[130])^(a[109] & b[131])^(a[108] & b[132])^(a[107] & b[133])^(a[106] & b[134])^(a[105] & b[135])^(a[104] & b[136])^(a[103] & b[137])^(a[102] & b[138])^(a[101] & b[139])^(a[100] & b[140])^(a[99] & b[141])^(a[98] & b[142])^(a[97] & b[143])^(a[96] & b[144])^(a[95] & b[145])^(a[94] & b[146])^(a[93] & b[147])^(a[92] & b[148])^(a[91] & b[149])^(a[90] & b[150])^(a[89] & b[151])^(a[88] & b[152])^(a[87] & b[153])^(a[86] & b[154])^(a[85] & b[155])^(a[84] & b[156])^(a[83] & b[157])^(a[82] & b[158])^(a[81] & b[159])^(a[80] & b[160])^(a[79] & b[161])^(a[78] & b[162])^(a[77] & b[163])^(a[76] & b[164])^(a[75] & b[165])^(a[74] & b[166])^(a[73] & b[167])^(a[72] & b[168])^(a[71] & b[169])^(a[70] & b[170])^(a[69] & b[171])^(a[68] & b[172])^(a[67] & b[173])^(a[66] & b[174])^(a[65] & b[175])^(a[64] & b[176])^(a[63] & b[177])^(a[62] & b[178])^(a[61] & b[179])^(a[60] & b[180])^(a[59] & b[181])^(a[58] & b[182])^(a[57] & b[183])^(a[56] & b[184])^(a[55] & b[185])^(a[54] & b[186])^(a[53] & b[187])^(a[52] & b[188])^(a[51] & b[189])^(a[50] & b[190])^(a[49] & b[191])^(a[48] & b[192])^(a[47] & b[193])^(a[46] & b[194])^(a[45] & b[195])^(a[44] & b[196])^(a[43] & b[197])^(a[42] & b[198])^(a[41] & b[199])^(a[40] & b[200])^(a[39] & b[201])^(a[38] & b[202])^(a[37] & b[203])^(a[36] & b[204])^(a[35] & b[205])^(a[34] & b[206])^(a[33] & b[207])^(a[32] & b[208])^(a[31] & b[209])^(a[30] & b[210])^(a[29] & b[211])^(a[28] & b[212])^(a[27] & b[213])^(a[26] & b[214])^(a[25] & b[215])^(a[24] & b[216])^(a[23] & b[217])^(a[22] & b[218])^(a[21] & b[219])^(a[20] & b[220])^(a[19] & b[221])^(a[18] & b[222])^(a[17] & b[223])^(a[16] & b[224])^(a[15] & b[225])^(a[14] & b[226])^(a[13] & b[227])^(a[12] & b[228])^(a[11] & b[229])^(a[10] & b[230])^(a[9] & b[231])^(a[8] & b[232])^(a[7] & b[233])^(a[6] & b[234])^(a[5] & b[235])^(a[4] & b[236])^(a[3] & b[237])^(a[2] & b[238])^(a[1] & b[239])^(a[0] & b[240]);
assign y[241] = (a[241] & b[0])^(a[240] & b[1])^(a[239] & b[2])^(a[238] & b[3])^(a[237] & b[4])^(a[236] & b[5])^(a[235] & b[6])^(a[234] & b[7])^(a[233] & b[8])^(a[232] & b[9])^(a[231] & b[10])^(a[230] & b[11])^(a[229] & b[12])^(a[228] & b[13])^(a[227] & b[14])^(a[226] & b[15])^(a[225] & b[16])^(a[224] & b[17])^(a[223] & b[18])^(a[222] & b[19])^(a[221] & b[20])^(a[220] & b[21])^(a[219] & b[22])^(a[218] & b[23])^(a[217] & b[24])^(a[216] & b[25])^(a[215] & b[26])^(a[214] & b[27])^(a[213] & b[28])^(a[212] & b[29])^(a[211] & b[30])^(a[210] & b[31])^(a[209] & b[32])^(a[208] & b[33])^(a[207] & b[34])^(a[206] & b[35])^(a[205] & b[36])^(a[204] & b[37])^(a[203] & b[38])^(a[202] & b[39])^(a[201] & b[40])^(a[200] & b[41])^(a[199] & b[42])^(a[198] & b[43])^(a[197] & b[44])^(a[196] & b[45])^(a[195] & b[46])^(a[194] & b[47])^(a[193] & b[48])^(a[192] & b[49])^(a[191] & b[50])^(a[190] & b[51])^(a[189] & b[52])^(a[188] & b[53])^(a[187] & b[54])^(a[186] & b[55])^(a[185] & b[56])^(a[184] & b[57])^(a[183] & b[58])^(a[182] & b[59])^(a[181] & b[60])^(a[180] & b[61])^(a[179] & b[62])^(a[178] & b[63])^(a[177] & b[64])^(a[176] & b[65])^(a[175] & b[66])^(a[174] & b[67])^(a[173] & b[68])^(a[172] & b[69])^(a[171] & b[70])^(a[170] & b[71])^(a[169] & b[72])^(a[168] & b[73])^(a[167] & b[74])^(a[166] & b[75])^(a[165] & b[76])^(a[164] & b[77])^(a[163] & b[78])^(a[162] & b[79])^(a[161] & b[80])^(a[160] & b[81])^(a[159] & b[82])^(a[158] & b[83])^(a[157] & b[84])^(a[156] & b[85])^(a[155] & b[86])^(a[154] & b[87])^(a[153] & b[88])^(a[152] & b[89])^(a[151] & b[90])^(a[150] & b[91])^(a[149] & b[92])^(a[148] & b[93])^(a[147] & b[94])^(a[146] & b[95])^(a[145] & b[96])^(a[144] & b[97])^(a[143] & b[98])^(a[142] & b[99])^(a[141] & b[100])^(a[140] & b[101])^(a[139] & b[102])^(a[138] & b[103])^(a[137] & b[104])^(a[136] & b[105])^(a[135] & b[106])^(a[134] & b[107])^(a[133] & b[108])^(a[132] & b[109])^(a[131] & b[110])^(a[130] & b[111])^(a[129] & b[112])^(a[128] & b[113])^(a[127] & b[114])^(a[126] & b[115])^(a[125] & b[116])^(a[124] & b[117])^(a[123] & b[118])^(a[122] & b[119])^(a[121] & b[120])^(a[120] & b[121])^(a[119] & b[122])^(a[118] & b[123])^(a[117] & b[124])^(a[116] & b[125])^(a[115] & b[126])^(a[114] & b[127])^(a[113] & b[128])^(a[112] & b[129])^(a[111] & b[130])^(a[110] & b[131])^(a[109] & b[132])^(a[108] & b[133])^(a[107] & b[134])^(a[106] & b[135])^(a[105] & b[136])^(a[104] & b[137])^(a[103] & b[138])^(a[102] & b[139])^(a[101] & b[140])^(a[100] & b[141])^(a[99] & b[142])^(a[98] & b[143])^(a[97] & b[144])^(a[96] & b[145])^(a[95] & b[146])^(a[94] & b[147])^(a[93] & b[148])^(a[92] & b[149])^(a[91] & b[150])^(a[90] & b[151])^(a[89] & b[152])^(a[88] & b[153])^(a[87] & b[154])^(a[86] & b[155])^(a[85] & b[156])^(a[84] & b[157])^(a[83] & b[158])^(a[82] & b[159])^(a[81] & b[160])^(a[80] & b[161])^(a[79] & b[162])^(a[78] & b[163])^(a[77] & b[164])^(a[76] & b[165])^(a[75] & b[166])^(a[74] & b[167])^(a[73] & b[168])^(a[72] & b[169])^(a[71] & b[170])^(a[70] & b[171])^(a[69] & b[172])^(a[68] & b[173])^(a[67] & b[174])^(a[66] & b[175])^(a[65] & b[176])^(a[64] & b[177])^(a[63] & b[178])^(a[62] & b[179])^(a[61] & b[180])^(a[60] & b[181])^(a[59] & b[182])^(a[58] & b[183])^(a[57] & b[184])^(a[56] & b[185])^(a[55] & b[186])^(a[54] & b[187])^(a[53] & b[188])^(a[52] & b[189])^(a[51] & b[190])^(a[50] & b[191])^(a[49] & b[192])^(a[48] & b[193])^(a[47] & b[194])^(a[46] & b[195])^(a[45] & b[196])^(a[44] & b[197])^(a[43] & b[198])^(a[42] & b[199])^(a[41] & b[200])^(a[40] & b[201])^(a[39] & b[202])^(a[38] & b[203])^(a[37] & b[204])^(a[36] & b[205])^(a[35] & b[206])^(a[34] & b[207])^(a[33] & b[208])^(a[32] & b[209])^(a[31] & b[210])^(a[30] & b[211])^(a[29] & b[212])^(a[28] & b[213])^(a[27] & b[214])^(a[26] & b[215])^(a[25] & b[216])^(a[24] & b[217])^(a[23] & b[218])^(a[22] & b[219])^(a[21] & b[220])^(a[20] & b[221])^(a[19] & b[222])^(a[18] & b[223])^(a[17] & b[224])^(a[16] & b[225])^(a[15] & b[226])^(a[14] & b[227])^(a[13] & b[228])^(a[12] & b[229])^(a[11] & b[230])^(a[10] & b[231])^(a[9] & b[232])^(a[8] & b[233])^(a[7] & b[234])^(a[6] & b[235])^(a[5] & b[236])^(a[4] & b[237])^(a[3] & b[238])^(a[2] & b[239])^(a[1] & b[240])^(a[0] & b[241]);
assign y[242] = (a[242] & b[0])^(a[241] & b[1])^(a[240] & b[2])^(a[239] & b[3])^(a[238] & b[4])^(a[237] & b[5])^(a[236] & b[6])^(a[235] & b[7])^(a[234] & b[8])^(a[233] & b[9])^(a[232] & b[10])^(a[231] & b[11])^(a[230] & b[12])^(a[229] & b[13])^(a[228] & b[14])^(a[227] & b[15])^(a[226] & b[16])^(a[225] & b[17])^(a[224] & b[18])^(a[223] & b[19])^(a[222] & b[20])^(a[221] & b[21])^(a[220] & b[22])^(a[219] & b[23])^(a[218] & b[24])^(a[217] & b[25])^(a[216] & b[26])^(a[215] & b[27])^(a[214] & b[28])^(a[213] & b[29])^(a[212] & b[30])^(a[211] & b[31])^(a[210] & b[32])^(a[209] & b[33])^(a[208] & b[34])^(a[207] & b[35])^(a[206] & b[36])^(a[205] & b[37])^(a[204] & b[38])^(a[203] & b[39])^(a[202] & b[40])^(a[201] & b[41])^(a[200] & b[42])^(a[199] & b[43])^(a[198] & b[44])^(a[197] & b[45])^(a[196] & b[46])^(a[195] & b[47])^(a[194] & b[48])^(a[193] & b[49])^(a[192] & b[50])^(a[191] & b[51])^(a[190] & b[52])^(a[189] & b[53])^(a[188] & b[54])^(a[187] & b[55])^(a[186] & b[56])^(a[185] & b[57])^(a[184] & b[58])^(a[183] & b[59])^(a[182] & b[60])^(a[181] & b[61])^(a[180] & b[62])^(a[179] & b[63])^(a[178] & b[64])^(a[177] & b[65])^(a[176] & b[66])^(a[175] & b[67])^(a[174] & b[68])^(a[173] & b[69])^(a[172] & b[70])^(a[171] & b[71])^(a[170] & b[72])^(a[169] & b[73])^(a[168] & b[74])^(a[167] & b[75])^(a[166] & b[76])^(a[165] & b[77])^(a[164] & b[78])^(a[163] & b[79])^(a[162] & b[80])^(a[161] & b[81])^(a[160] & b[82])^(a[159] & b[83])^(a[158] & b[84])^(a[157] & b[85])^(a[156] & b[86])^(a[155] & b[87])^(a[154] & b[88])^(a[153] & b[89])^(a[152] & b[90])^(a[151] & b[91])^(a[150] & b[92])^(a[149] & b[93])^(a[148] & b[94])^(a[147] & b[95])^(a[146] & b[96])^(a[145] & b[97])^(a[144] & b[98])^(a[143] & b[99])^(a[142] & b[100])^(a[141] & b[101])^(a[140] & b[102])^(a[139] & b[103])^(a[138] & b[104])^(a[137] & b[105])^(a[136] & b[106])^(a[135] & b[107])^(a[134] & b[108])^(a[133] & b[109])^(a[132] & b[110])^(a[131] & b[111])^(a[130] & b[112])^(a[129] & b[113])^(a[128] & b[114])^(a[127] & b[115])^(a[126] & b[116])^(a[125] & b[117])^(a[124] & b[118])^(a[123] & b[119])^(a[122] & b[120])^(a[121] & b[121])^(a[120] & b[122])^(a[119] & b[123])^(a[118] & b[124])^(a[117] & b[125])^(a[116] & b[126])^(a[115] & b[127])^(a[114] & b[128])^(a[113] & b[129])^(a[112] & b[130])^(a[111] & b[131])^(a[110] & b[132])^(a[109] & b[133])^(a[108] & b[134])^(a[107] & b[135])^(a[106] & b[136])^(a[105] & b[137])^(a[104] & b[138])^(a[103] & b[139])^(a[102] & b[140])^(a[101] & b[141])^(a[100] & b[142])^(a[99] & b[143])^(a[98] & b[144])^(a[97] & b[145])^(a[96] & b[146])^(a[95] & b[147])^(a[94] & b[148])^(a[93] & b[149])^(a[92] & b[150])^(a[91] & b[151])^(a[90] & b[152])^(a[89] & b[153])^(a[88] & b[154])^(a[87] & b[155])^(a[86] & b[156])^(a[85] & b[157])^(a[84] & b[158])^(a[83] & b[159])^(a[82] & b[160])^(a[81] & b[161])^(a[80] & b[162])^(a[79] & b[163])^(a[78] & b[164])^(a[77] & b[165])^(a[76] & b[166])^(a[75] & b[167])^(a[74] & b[168])^(a[73] & b[169])^(a[72] & b[170])^(a[71] & b[171])^(a[70] & b[172])^(a[69] & b[173])^(a[68] & b[174])^(a[67] & b[175])^(a[66] & b[176])^(a[65] & b[177])^(a[64] & b[178])^(a[63] & b[179])^(a[62] & b[180])^(a[61] & b[181])^(a[60] & b[182])^(a[59] & b[183])^(a[58] & b[184])^(a[57] & b[185])^(a[56] & b[186])^(a[55] & b[187])^(a[54] & b[188])^(a[53] & b[189])^(a[52] & b[190])^(a[51] & b[191])^(a[50] & b[192])^(a[49] & b[193])^(a[48] & b[194])^(a[47] & b[195])^(a[46] & b[196])^(a[45] & b[197])^(a[44] & b[198])^(a[43] & b[199])^(a[42] & b[200])^(a[41] & b[201])^(a[40] & b[202])^(a[39] & b[203])^(a[38] & b[204])^(a[37] & b[205])^(a[36] & b[206])^(a[35] & b[207])^(a[34] & b[208])^(a[33] & b[209])^(a[32] & b[210])^(a[31] & b[211])^(a[30] & b[212])^(a[29] & b[213])^(a[28] & b[214])^(a[27] & b[215])^(a[26] & b[216])^(a[25] & b[217])^(a[24] & b[218])^(a[23] & b[219])^(a[22] & b[220])^(a[21] & b[221])^(a[20] & b[222])^(a[19] & b[223])^(a[18] & b[224])^(a[17] & b[225])^(a[16] & b[226])^(a[15] & b[227])^(a[14] & b[228])^(a[13] & b[229])^(a[12] & b[230])^(a[11] & b[231])^(a[10] & b[232])^(a[9] & b[233])^(a[8] & b[234])^(a[7] & b[235])^(a[6] & b[236])^(a[5] & b[237])^(a[4] & b[238])^(a[3] & b[239])^(a[2] & b[240])^(a[1] & b[241])^(a[0] & b[242]);
assign y[243] = (a[243] & b[0])^(a[242] & b[1])^(a[241] & b[2])^(a[240] & b[3])^(a[239] & b[4])^(a[238] & b[5])^(a[237] & b[6])^(a[236] & b[7])^(a[235] & b[8])^(a[234] & b[9])^(a[233] & b[10])^(a[232] & b[11])^(a[231] & b[12])^(a[230] & b[13])^(a[229] & b[14])^(a[228] & b[15])^(a[227] & b[16])^(a[226] & b[17])^(a[225] & b[18])^(a[224] & b[19])^(a[223] & b[20])^(a[222] & b[21])^(a[221] & b[22])^(a[220] & b[23])^(a[219] & b[24])^(a[218] & b[25])^(a[217] & b[26])^(a[216] & b[27])^(a[215] & b[28])^(a[214] & b[29])^(a[213] & b[30])^(a[212] & b[31])^(a[211] & b[32])^(a[210] & b[33])^(a[209] & b[34])^(a[208] & b[35])^(a[207] & b[36])^(a[206] & b[37])^(a[205] & b[38])^(a[204] & b[39])^(a[203] & b[40])^(a[202] & b[41])^(a[201] & b[42])^(a[200] & b[43])^(a[199] & b[44])^(a[198] & b[45])^(a[197] & b[46])^(a[196] & b[47])^(a[195] & b[48])^(a[194] & b[49])^(a[193] & b[50])^(a[192] & b[51])^(a[191] & b[52])^(a[190] & b[53])^(a[189] & b[54])^(a[188] & b[55])^(a[187] & b[56])^(a[186] & b[57])^(a[185] & b[58])^(a[184] & b[59])^(a[183] & b[60])^(a[182] & b[61])^(a[181] & b[62])^(a[180] & b[63])^(a[179] & b[64])^(a[178] & b[65])^(a[177] & b[66])^(a[176] & b[67])^(a[175] & b[68])^(a[174] & b[69])^(a[173] & b[70])^(a[172] & b[71])^(a[171] & b[72])^(a[170] & b[73])^(a[169] & b[74])^(a[168] & b[75])^(a[167] & b[76])^(a[166] & b[77])^(a[165] & b[78])^(a[164] & b[79])^(a[163] & b[80])^(a[162] & b[81])^(a[161] & b[82])^(a[160] & b[83])^(a[159] & b[84])^(a[158] & b[85])^(a[157] & b[86])^(a[156] & b[87])^(a[155] & b[88])^(a[154] & b[89])^(a[153] & b[90])^(a[152] & b[91])^(a[151] & b[92])^(a[150] & b[93])^(a[149] & b[94])^(a[148] & b[95])^(a[147] & b[96])^(a[146] & b[97])^(a[145] & b[98])^(a[144] & b[99])^(a[143] & b[100])^(a[142] & b[101])^(a[141] & b[102])^(a[140] & b[103])^(a[139] & b[104])^(a[138] & b[105])^(a[137] & b[106])^(a[136] & b[107])^(a[135] & b[108])^(a[134] & b[109])^(a[133] & b[110])^(a[132] & b[111])^(a[131] & b[112])^(a[130] & b[113])^(a[129] & b[114])^(a[128] & b[115])^(a[127] & b[116])^(a[126] & b[117])^(a[125] & b[118])^(a[124] & b[119])^(a[123] & b[120])^(a[122] & b[121])^(a[121] & b[122])^(a[120] & b[123])^(a[119] & b[124])^(a[118] & b[125])^(a[117] & b[126])^(a[116] & b[127])^(a[115] & b[128])^(a[114] & b[129])^(a[113] & b[130])^(a[112] & b[131])^(a[111] & b[132])^(a[110] & b[133])^(a[109] & b[134])^(a[108] & b[135])^(a[107] & b[136])^(a[106] & b[137])^(a[105] & b[138])^(a[104] & b[139])^(a[103] & b[140])^(a[102] & b[141])^(a[101] & b[142])^(a[100] & b[143])^(a[99] & b[144])^(a[98] & b[145])^(a[97] & b[146])^(a[96] & b[147])^(a[95] & b[148])^(a[94] & b[149])^(a[93] & b[150])^(a[92] & b[151])^(a[91] & b[152])^(a[90] & b[153])^(a[89] & b[154])^(a[88] & b[155])^(a[87] & b[156])^(a[86] & b[157])^(a[85] & b[158])^(a[84] & b[159])^(a[83] & b[160])^(a[82] & b[161])^(a[81] & b[162])^(a[80] & b[163])^(a[79] & b[164])^(a[78] & b[165])^(a[77] & b[166])^(a[76] & b[167])^(a[75] & b[168])^(a[74] & b[169])^(a[73] & b[170])^(a[72] & b[171])^(a[71] & b[172])^(a[70] & b[173])^(a[69] & b[174])^(a[68] & b[175])^(a[67] & b[176])^(a[66] & b[177])^(a[65] & b[178])^(a[64] & b[179])^(a[63] & b[180])^(a[62] & b[181])^(a[61] & b[182])^(a[60] & b[183])^(a[59] & b[184])^(a[58] & b[185])^(a[57] & b[186])^(a[56] & b[187])^(a[55] & b[188])^(a[54] & b[189])^(a[53] & b[190])^(a[52] & b[191])^(a[51] & b[192])^(a[50] & b[193])^(a[49] & b[194])^(a[48] & b[195])^(a[47] & b[196])^(a[46] & b[197])^(a[45] & b[198])^(a[44] & b[199])^(a[43] & b[200])^(a[42] & b[201])^(a[41] & b[202])^(a[40] & b[203])^(a[39] & b[204])^(a[38] & b[205])^(a[37] & b[206])^(a[36] & b[207])^(a[35] & b[208])^(a[34] & b[209])^(a[33] & b[210])^(a[32] & b[211])^(a[31] & b[212])^(a[30] & b[213])^(a[29] & b[214])^(a[28] & b[215])^(a[27] & b[216])^(a[26] & b[217])^(a[25] & b[218])^(a[24] & b[219])^(a[23] & b[220])^(a[22] & b[221])^(a[21] & b[222])^(a[20] & b[223])^(a[19] & b[224])^(a[18] & b[225])^(a[17] & b[226])^(a[16] & b[227])^(a[15] & b[228])^(a[14] & b[229])^(a[13] & b[230])^(a[12] & b[231])^(a[11] & b[232])^(a[10] & b[233])^(a[9] & b[234])^(a[8] & b[235])^(a[7] & b[236])^(a[6] & b[237])^(a[5] & b[238])^(a[4] & b[239])^(a[3] & b[240])^(a[2] & b[241])^(a[1] & b[242])^(a[0] & b[243]);
assign y[244] = (a[244] & b[0])^(a[243] & b[1])^(a[242] & b[2])^(a[241] & b[3])^(a[240] & b[4])^(a[239] & b[5])^(a[238] & b[6])^(a[237] & b[7])^(a[236] & b[8])^(a[235] & b[9])^(a[234] & b[10])^(a[233] & b[11])^(a[232] & b[12])^(a[231] & b[13])^(a[230] & b[14])^(a[229] & b[15])^(a[228] & b[16])^(a[227] & b[17])^(a[226] & b[18])^(a[225] & b[19])^(a[224] & b[20])^(a[223] & b[21])^(a[222] & b[22])^(a[221] & b[23])^(a[220] & b[24])^(a[219] & b[25])^(a[218] & b[26])^(a[217] & b[27])^(a[216] & b[28])^(a[215] & b[29])^(a[214] & b[30])^(a[213] & b[31])^(a[212] & b[32])^(a[211] & b[33])^(a[210] & b[34])^(a[209] & b[35])^(a[208] & b[36])^(a[207] & b[37])^(a[206] & b[38])^(a[205] & b[39])^(a[204] & b[40])^(a[203] & b[41])^(a[202] & b[42])^(a[201] & b[43])^(a[200] & b[44])^(a[199] & b[45])^(a[198] & b[46])^(a[197] & b[47])^(a[196] & b[48])^(a[195] & b[49])^(a[194] & b[50])^(a[193] & b[51])^(a[192] & b[52])^(a[191] & b[53])^(a[190] & b[54])^(a[189] & b[55])^(a[188] & b[56])^(a[187] & b[57])^(a[186] & b[58])^(a[185] & b[59])^(a[184] & b[60])^(a[183] & b[61])^(a[182] & b[62])^(a[181] & b[63])^(a[180] & b[64])^(a[179] & b[65])^(a[178] & b[66])^(a[177] & b[67])^(a[176] & b[68])^(a[175] & b[69])^(a[174] & b[70])^(a[173] & b[71])^(a[172] & b[72])^(a[171] & b[73])^(a[170] & b[74])^(a[169] & b[75])^(a[168] & b[76])^(a[167] & b[77])^(a[166] & b[78])^(a[165] & b[79])^(a[164] & b[80])^(a[163] & b[81])^(a[162] & b[82])^(a[161] & b[83])^(a[160] & b[84])^(a[159] & b[85])^(a[158] & b[86])^(a[157] & b[87])^(a[156] & b[88])^(a[155] & b[89])^(a[154] & b[90])^(a[153] & b[91])^(a[152] & b[92])^(a[151] & b[93])^(a[150] & b[94])^(a[149] & b[95])^(a[148] & b[96])^(a[147] & b[97])^(a[146] & b[98])^(a[145] & b[99])^(a[144] & b[100])^(a[143] & b[101])^(a[142] & b[102])^(a[141] & b[103])^(a[140] & b[104])^(a[139] & b[105])^(a[138] & b[106])^(a[137] & b[107])^(a[136] & b[108])^(a[135] & b[109])^(a[134] & b[110])^(a[133] & b[111])^(a[132] & b[112])^(a[131] & b[113])^(a[130] & b[114])^(a[129] & b[115])^(a[128] & b[116])^(a[127] & b[117])^(a[126] & b[118])^(a[125] & b[119])^(a[124] & b[120])^(a[123] & b[121])^(a[122] & b[122])^(a[121] & b[123])^(a[120] & b[124])^(a[119] & b[125])^(a[118] & b[126])^(a[117] & b[127])^(a[116] & b[128])^(a[115] & b[129])^(a[114] & b[130])^(a[113] & b[131])^(a[112] & b[132])^(a[111] & b[133])^(a[110] & b[134])^(a[109] & b[135])^(a[108] & b[136])^(a[107] & b[137])^(a[106] & b[138])^(a[105] & b[139])^(a[104] & b[140])^(a[103] & b[141])^(a[102] & b[142])^(a[101] & b[143])^(a[100] & b[144])^(a[99] & b[145])^(a[98] & b[146])^(a[97] & b[147])^(a[96] & b[148])^(a[95] & b[149])^(a[94] & b[150])^(a[93] & b[151])^(a[92] & b[152])^(a[91] & b[153])^(a[90] & b[154])^(a[89] & b[155])^(a[88] & b[156])^(a[87] & b[157])^(a[86] & b[158])^(a[85] & b[159])^(a[84] & b[160])^(a[83] & b[161])^(a[82] & b[162])^(a[81] & b[163])^(a[80] & b[164])^(a[79] & b[165])^(a[78] & b[166])^(a[77] & b[167])^(a[76] & b[168])^(a[75] & b[169])^(a[74] & b[170])^(a[73] & b[171])^(a[72] & b[172])^(a[71] & b[173])^(a[70] & b[174])^(a[69] & b[175])^(a[68] & b[176])^(a[67] & b[177])^(a[66] & b[178])^(a[65] & b[179])^(a[64] & b[180])^(a[63] & b[181])^(a[62] & b[182])^(a[61] & b[183])^(a[60] & b[184])^(a[59] & b[185])^(a[58] & b[186])^(a[57] & b[187])^(a[56] & b[188])^(a[55] & b[189])^(a[54] & b[190])^(a[53] & b[191])^(a[52] & b[192])^(a[51] & b[193])^(a[50] & b[194])^(a[49] & b[195])^(a[48] & b[196])^(a[47] & b[197])^(a[46] & b[198])^(a[45] & b[199])^(a[44] & b[200])^(a[43] & b[201])^(a[42] & b[202])^(a[41] & b[203])^(a[40] & b[204])^(a[39] & b[205])^(a[38] & b[206])^(a[37] & b[207])^(a[36] & b[208])^(a[35] & b[209])^(a[34] & b[210])^(a[33] & b[211])^(a[32] & b[212])^(a[31] & b[213])^(a[30] & b[214])^(a[29] & b[215])^(a[28] & b[216])^(a[27] & b[217])^(a[26] & b[218])^(a[25] & b[219])^(a[24] & b[220])^(a[23] & b[221])^(a[22] & b[222])^(a[21] & b[223])^(a[20] & b[224])^(a[19] & b[225])^(a[18] & b[226])^(a[17] & b[227])^(a[16] & b[228])^(a[15] & b[229])^(a[14] & b[230])^(a[13] & b[231])^(a[12] & b[232])^(a[11] & b[233])^(a[10] & b[234])^(a[9] & b[235])^(a[8] & b[236])^(a[7] & b[237])^(a[6] & b[238])^(a[5] & b[239])^(a[4] & b[240])^(a[3] & b[241])^(a[2] & b[242])^(a[1] & b[243])^(a[0] & b[244]);
assign y[245] = (a[245] & b[0])^(a[244] & b[1])^(a[243] & b[2])^(a[242] & b[3])^(a[241] & b[4])^(a[240] & b[5])^(a[239] & b[6])^(a[238] & b[7])^(a[237] & b[8])^(a[236] & b[9])^(a[235] & b[10])^(a[234] & b[11])^(a[233] & b[12])^(a[232] & b[13])^(a[231] & b[14])^(a[230] & b[15])^(a[229] & b[16])^(a[228] & b[17])^(a[227] & b[18])^(a[226] & b[19])^(a[225] & b[20])^(a[224] & b[21])^(a[223] & b[22])^(a[222] & b[23])^(a[221] & b[24])^(a[220] & b[25])^(a[219] & b[26])^(a[218] & b[27])^(a[217] & b[28])^(a[216] & b[29])^(a[215] & b[30])^(a[214] & b[31])^(a[213] & b[32])^(a[212] & b[33])^(a[211] & b[34])^(a[210] & b[35])^(a[209] & b[36])^(a[208] & b[37])^(a[207] & b[38])^(a[206] & b[39])^(a[205] & b[40])^(a[204] & b[41])^(a[203] & b[42])^(a[202] & b[43])^(a[201] & b[44])^(a[200] & b[45])^(a[199] & b[46])^(a[198] & b[47])^(a[197] & b[48])^(a[196] & b[49])^(a[195] & b[50])^(a[194] & b[51])^(a[193] & b[52])^(a[192] & b[53])^(a[191] & b[54])^(a[190] & b[55])^(a[189] & b[56])^(a[188] & b[57])^(a[187] & b[58])^(a[186] & b[59])^(a[185] & b[60])^(a[184] & b[61])^(a[183] & b[62])^(a[182] & b[63])^(a[181] & b[64])^(a[180] & b[65])^(a[179] & b[66])^(a[178] & b[67])^(a[177] & b[68])^(a[176] & b[69])^(a[175] & b[70])^(a[174] & b[71])^(a[173] & b[72])^(a[172] & b[73])^(a[171] & b[74])^(a[170] & b[75])^(a[169] & b[76])^(a[168] & b[77])^(a[167] & b[78])^(a[166] & b[79])^(a[165] & b[80])^(a[164] & b[81])^(a[163] & b[82])^(a[162] & b[83])^(a[161] & b[84])^(a[160] & b[85])^(a[159] & b[86])^(a[158] & b[87])^(a[157] & b[88])^(a[156] & b[89])^(a[155] & b[90])^(a[154] & b[91])^(a[153] & b[92])^(a[152] & b[93])^(a[151] & b[94])^(a[150] & b[95])^(a[149] & b[96])^(a[148] & b[97])^(a[147] & b[98])^(a[146] & b[99])^(a[145] & b[100])^(a[144] & b[101])^(a[143] & b[102])^(a[142] & b[103])^(a[141] & b[104])^(a[140] & b[105])^(a[139] & b[106])^(a[138] & b[107])^(a[137] & b[108])^(a[136] & b[109])^(a[135] & b[110])^(a[134] & b[111])^(a[133] & b[112])^(a[132] & b[113])^(a[131] & b[114])^(a[130] & b[115])^(a[129] & b[116])^(a[128] & b[117])^(a[127] & b[118])^(a[126] & b[119])^(a[125] & b[120])^(a[124] & b[121])^(a[123] & b[122])^(a[122] & b[123])^(a[121] & b[124])^(a[120] & b[125])^(a[119] & b[126])^(a[118] & b[127])^(a[117] & b[128])^(a[116] & b[129])^(a[115] & b[130])^(a[114] & b[131])^(a[113] & b[132])^(a[112] & b[133])^(a[111] & b[134])^(a[110] & b[135])^(a[109] & b[136])^(a[108] & b[137])^(a[107] & b[138])^(a[106] & b[139])^(a[105] & b[140])^(a[104] & b[141])^(a[103] & b[142])^(a[102] & b[143])^(a[101] & b[144])^(a[100] & b[145])^(a[99] & b[146])^(a[98] & b[147])^(a[97] & b[148])^(a[96] & b[149])^(a[95] & b[150])^(a[94] & b[151])^(a[93] & b[152])^(a[92] & b[153])^(a[91] & b[154])^(a[90] & b[155])^(a[89] & b[156])^(a[88] & b[157])^(a[87] & b[158])^(a[86] & b[159])^(a[85] & b[160])^(a[84] & b[161])^(a[83] & b[162])^(a[82] & b[163])^(a[81] & b[164])^(a[80] & b[165])^(a[79] & b[166])^(a[78] & b[167])^(a[77] & b[168])^(a[76] & b[169])^(a[75] & b[170])^(a[74] & b[171])^(a[73] & b[172])^(a[72] & b[173])^(a[71] & b[174])^(a[70] & b[175])^(a[69] & b[176])^(a[68] & b[177])^(a[67] & b[178])^(a[66] & b[179])^(a[65] & b[180])^(a[64] & b[181])^(a[63] & b[182])^(a[62] & b[183])^(a[61] & b[184])^(a[60] & b[185])^(a[59] & b[186])^(a[58] & b[187])^(a[57] & b[188])^(a[56] & b[189])^(a[55] & b[190])^(a[54] & b[191])^(a[53] & b[192])^(a[52] & b[193])^(a[51] & b[194])^(a[50] & b[195])^(a[49] & b[196])^(a[48] & b[197])^(a[47] & b[198])^(a[46] & b[199])^(a[45] & b[200])^(a[44] & b[201])^(a[43] & b[202])^(a[42] & b[203])^(a[41] & b[204])^(a[40] & b[205])^(a[39] & b[206])^(a[38] & b[207])^(a[37] & b[208])^(a[36] & b[209])^(a[35] & b[210])^(a[34] & b[211])^(a[33] & b[212])^(a[32] & b[213])^(a[31] & b[214])^(a[30] & b[215])^(a[29] & b[216])^(a[28] & b[217])^(a[27] & b[218])^(a[26] & b[219])^(a[25] & b[220])^(a[24] & b[221])^(a[23] & b[222])^(a[22] & b[223])^(a[21] & b[224])^(a[20] & b[225])^(a[19] & b[226])^(a[18] & b[227])^(a[17] & b[228])^(a[16] & b[229])^(a[15] & b[230])^(a[14] & b[231])^(a[13] & b[232])^(a[12] & b[233])^(a[11] & b[234])^(a[10] & b[235])^(a[9] & b[236])^(a[8] & b[237])^(a[7] & b[238])^(a[6] & b[239])^(a[5] & b[240])^(a[4] & b[241])^(a[3] & b[242])^(a[2] & b[243])^(a[1] & b[244])^(a[0] & b[245]);
assign y[246] = (a[246] & b[0])^(a[245] & b[1])^(a[244] & b[2])^(a[243] & b[3])^(a[242] & b[4])^(a[241] & b[5])^(a[240] & b[6])^(a[239] & b[7])^(a[238] & b[8])^(a[237] & b[9])^(a[236] & b[10])^(a[235] & b[11])^(a[234] & b[12])^(a[233] & b[13])^(a[232] & b[14])^(a[231] & b[15])^(a[230] & b[16])^(a[229] & b[17])^(a[228] & b[18])^(a[227] & b[19])^(a[226] & b[20])^(a[225] & b[21])^(a[224] & b[22])^(a[223] & b[23])^(a[222] & b[24])^(a[221] & b[25])^(a[220] & b[26])^(a[219] & b[27])^(a[218] & b[28])^(a[217] & b[29])^(a[216] & b[30])^(a[215] & b[31])^(a[214] & b[32])^(a[213] & b[33])^(a[212] & b[34])^(a[211] & b[35])^(a[210] & b[36])^(a[209] & b[37])^(a[208] & b[38])^(a[207] & b[39])^(a[206] & b[40])^(a[205] & b[41])^(a[204] & b[42])^(a[203] & b[43])^(a[202] & b[44])^(a[201] & b[45])^(a[200] & b[46])^(a[199] & b[47])^(a[198] & b[48])^(a[197] & b[49])^(a[196] & b[50])^(a[195] & b[51])^(a[194] & b[52])^(a[193] & b[53])^(a[192] & b[54])^(a[191] & b[55])^(a[190] & b[56])^(a[189] & b[57])^(a[188] & b[58])^(a[187] & b[59])^(a[186] & b[60])^(a[185] & b[61])^(a[184] & b[62])^(a[183] & b[63])^(a[182] & b[64])^(a[181] & b[65])^(a[180] & b[66])^(a[179] & b[67])^(a[178] & b[68])^(a[177] & b[69])^(a[176] & b[70])^(a[175] & b[71])^(a[174] & b[72])^(a[173] & b[73])^(a[172] & b[74])^(a[171] & b[75])^(a[170] & b[76])^(a[169] & b[77])^(a[168] & b[78])^(a[167] & b[79])^(a[166] & b[80])^(a[165] & b[81])^(a[164] & b[82])^(a[163] & b[83])^(a[162] & b[84])^(a[161] & b[85])^(a[160] & b[86])^(a[159] & b[87])^(a[158] & b[88])^(a[157] & b[89])^(a[156] & b[90])^(a[155] & b[91])^(a[154] & b[92])^(a[153] & b[93])^(a[152] & b[94])^(a[151] & b[95])^(a[150] & b[96])^(a[149] & b[97])^(a[148] & b[98])^(a[147] & b[99])^(a[146] & b[100])^(a[145] & b[101])^(a[144] & b[102])^(a[143] & b[103])^(a[142] & b[104])^(a[141] & b[105])^(a[140] & b[106])^(a[139] & b[107])^(a[138] & b[108])^(a[137] & b[109])^(a[136] & b[110])^(a[135] & b[111])^(a[134] & b[112])^(a[133] & b[113])^(a[132] & b[114])^(a[131] & b[115])^(a[130] & b[116])^(a[129] & b[117])^(a[128] & b[118])^(a[127] & b[119])^(a[126] & b[120])^(a[125] & b[121])^(a[124] & b[122])^(a[123] & b[123])^(a[122] & b[124])^(a[121] & b[125])^(a[120] & b[126])^(a[119] & b[127])^(a[118] & b[128])^(a[117] & b[129])^(a[116] & b[130])^(a[115] & b[131])^(a[114] & b[132])^(a[113] & b[133])^(a[112] & b[134])^(a[111] & b[135])^(a[110] & b[136])^(a[109] & b[137])^(a[108] & b[138])^(a[107] & b[139])^(a[106] & b[140])^(a[105] & b[141])^(a[104] & b[142])^(a[103] & b[143])^(a[102] & b[144])^(a[101] & b[145])^(a[100] & b[146])^(a[99] & b[147])^(a[98] & b[148])^(a[97] & b[149])^(a[96] & b[150])^(a[95] & b[151])^(a[94] & b[152])^(a[93] & b[153])^(a[92] & b[154])^(a[91] & b[155])^(a[90] & b[156])^(a[89] & b[157])^(a[88] & b[158])^(a[87] & b[159])^(a[86] & b[160])^(a[85] & b[161])^(a[84] & b[162])^(a[83] & b[163])^(a[82] & b[164])^(a[81] & b[165])^(a[80] & b[166])^(a[79] & b[167])^(a[78] & b[168])^(a[77] & b[169])^(a[76] & b[170])^(a[75] & b[171])^(a[74] & b[172])^(a[73] & b[173])^(a[72] & b[174])^(a[71] & b[175])^(a[70] & b[176])^(a[69] & b[177])^(a[68] & b[178])^(a[67] & b[179])^(a[66] & b[180])^(a[65] & b[181])^(a[64] & b[182])^(a[63] & b[183])^(a[62] & b[184])^(a[61] & b[185])^(a[60] & b[186])^(a[59] & b[187])^(a[58] & b[188])^(a[57] & b[189])^(a[56] & b[190])^(a[55] & b[191])^(a[54] & b[192])^(a[53] & b[193])^(a[52] & b[194])^(a[51] & b[195])^(a[50] & b[196])^(a[49] & b[197])^(a[48] & b[198])^(a[47] & b[199])^(a[46] & b[200])^(a[45] & b[201])^(a[44] & b[202])^(a[43] & b[203])^(a[42] & b[204])^(a[41] & b[205])^(a[40] & b[206])^(a[39] & b[207])^(a[38] & b[208])^(a[37] & b[209])^(a[36] & b[210])^(a[35] & b[211])^(a[34] & b[212])^(a[33] & b[213])^(a[32] & b[214])^(a[31] & b[215])^(a[30] & b[216])^(a[29] & b[217])^(a[28] & b[218])^(a[27] & b[219])^(a[26] & b[220])^(a[25] & b[221])^(a[24] & b[222])^(a[23] & b[223])^(a[22] & b[224])^(a[21] & b[225])^(a[20] & b[226])^(a[19] & b[227])^(a[18] & b[228])^(a[17] & b[229])^(a[16] & b[230])^(a[15] & b[231])^(a[14] & b[232])^(a[13] & b[233])^(a[12] & b[234])^(a[11] & b[235])^(a[10] & b[236])^(a[9] & b[237])^(a[8] & b[238])^(a[7] & b[239])^(a[6] & b[240])^(a[5] & b[241])^(a[4] & b[242])^(a[3] & b[243])^(a[2] & b[244])^(a[1] & b[245])^(a[0] & b[246]);
assign y[247] = (a[247] & b[0])^(a[246] & b[1])^(a[245] & b[2])^(a[244] & b[3])^(a[243] & b[4])^(a[242] & b[5])^(a[241] & b[6])^(a[240] & b[7])^(a[239] & b[8])^(a[238] & b[9])^(a[237] & b[10])^(a[236] & b[11])^(a[235] & b[12])^(a[234] & b[13])^(a[233] & b[14])^(a[232] & b[15])^(a[231] & b[16])^(a[230] & b[17])^(a[229] & b[18])^(a[228] & b[19])^(a[227] & b[20])^(a[226] & b[21])^(a[225] & b[22])^(a[224] & b[23])^(a[223] & b[24])^(a[222] & b[25])^(a[221] & b[26])^(a[220] & b[27])^(a[219] & b[28])^(a[218] & b[29])^(a[217] & b[30])^(a[216] & b[31])^(a[215] & b[32])^(a[214] & b[33])^(a[213] & b[34])^(a[212] & b[35])^(a[211] & b[36])^(a[210] & b[37])^(a[209] & b[38])^(a[208] & b[39])^(a[207] & b[40])^(a[206] & b[41])^(a[205] & b[42])^(a[204] & b[43])^(a[203] & b[44])^(a[202] & b[45])^(a[201] & b[46])^(a[200] & b[47])^(a[199] & b[48])^(a[198] & b[49])^(a[197] & b[50])^(a[196] & b[51])^(a[195] & b[52])^(a[194] & b[53])^(a[193] & b[54])^(a[192] & b[55])^(a[191] & b[56])^(a[190] & b[57])^(a[189] & b[58])^(a[188] & b[59])^(a[187] & b[60])^(a[186] & b[61])^(a[185] & b[62])^(a[184] & b[63])^(a[183] & b[64])^(a[182] & b[65])^(a[181] & b[66])^(a[180] & b[67])^(a[179] & b[68])^(a[178] & b[69])^(a[177] & b[70])^(a[176] & b[71])^(a[175] & b[72])^(a[174] & b[73])^(a[173] & b[74])^(a[172] & b[75])^(a[171] & b[76])^(a[170] & b[77])^(a[169] & b[78])^(a[168] & b[79])^(a[167] & b[80])^(a[166] & b[81])^(a[165] & b[82])^(a[164] & b[83])^(a[163] & b[84])^(a[162] & b[85])^(a[161] & b[86])^(a[160] & b[87])^(a[159] & b[88])^(a[158] & b[89])^(a[157] & b[90])^(a[156] & b[91])^(a[155] & b[92])^(a[154] & b[93])^(a[153] & b[94])^(a[152] & b[95])^(a[151] & b[96])^(a[150] & b[97])^(a[149] & b[98])^(a[148] & b[99])^(a[147] & b[100])^(a[146] & b[101])^(a[145] & b[102])^(a[144] & b[103])^(a[143] & b[104])^(a[142] & b[105])^(a[141] & b[106])^(a[140] & b[107])^(a[139] & b[108])^(a[138] & b[109])^(a[137] & b[110])^(a[136] & b[111])^(a[135] & b[112])^(a[134] & b[113])^(a[133] & b[114])^(a[132] & b[115])^(a[131] & b[116])^(a[130] & b[117])^(a[129] & b[118])^(a[128] & b[119])^(a[127] & b[120])^(a[126] & b[121])^(a[125] & b[122])^(a[124] & b[123])^(a[123] & b[124])^(a[122] & b[125])^(a[121] & b[126])^(a[120] & b[127])^(a[119] & b[128])^(a[118] & b[129])^(a[117] & b[130])^(a[116] & b[131])^(a[115] & b[132])^(a[114] & b[133])^(a[113] & b[134])^(a[112] & b[135])^(a[111] & b[136])^(a[110] & b[137])^(a[109] & b[138])^(a[108] & b[139])^(a[107] & b[140])^(a[106] & b[141])^(a[105] & b[142])^(a[104] & b[143])^(a[103] & b[144])^(a[102] & b[145])^(a[101] & b[146])^(a[100] & b[147])^(a[99] & b[148])^(a[98] & b[149])^(a[97] & b[150])^(a[96] & b[151])^(a[95] & b[152])^(a[94] & b[153])^(a[93] & b[154])^(a[92] & b[155])^(a[91] & b[156])^(a[90] & b[157])^(a[89] & b[158])^(a[88] & b[159])^(a[87] & b[160])^(a[86] & b[161])^(a[85] & b[162])^(a[84] & b[163])^(a[83] & b[164])^(a[82] & b[165])^(a[81] & b[166])^(a[80] & b[167])^(a[79] & b[168])^(a[78] & b[169])^(a[77] & b[170])^(a[76] & b[171])^(a[75] & b[172])^(a[74] & b[173])^(a[73] & b[174])^(a[72] & b[175])^(a[71] & b[176])^(a[70] & b[177])^(a[69] & b[178])^(a[68] & b[179])^(a[67] & b[180])^(a[66] & b[181])^(a[65] & b[182])^(a[64] & b[183])^(a[63] & b[184])^(a[62] & b[185])^(a[61] & b[186])^(a[60] & b[187])^(a[59] & b[188])^(a[58] & b[189])^(a[57] & b[190])^(a[56] & b[191])^(a[55] & b[192])^(a[54] & b[193])^(a[53] & b[194])^(a[52] & b[195])^(a[51] & b[196])^(a[50] & b[197])^(a[49] & b[198])^(a[48] & b[199])^(a[47] & b[200])^(a[46] & b[201])^(a[45] & b[202])^(a[44] & b[203])^(a[43] & b[204])^(a[42] & b[205])^(a[41] & b[206])^(a[40] & b[207])^(a[39] & b[208])^(a[38] & b[209])^(a[37] & b[210])^(a[36] & b[211])^(a[35] & b[212])^(a[34] & b[213])^(a[33] & b[214])^(a[32] & b[215])^(a[31] & b[216])^(a[30] & b[217])^(a[29] & b[218])^(a[28] & b[219])^(a[27] & b[220])^(a[26] & b[221])^(a[25] & b[222])^(a[24] & b[223])^(a[23] & b[224])^(a[22] & b[225])^(a[21] & b[226])^(a[20] & b[227])^(a[19] & b[228])^(a[18] & b[229])^(a[17] & b[230])^(a[16] & b[231])^(a[15] & b[232])^(a[14] & b[233])^(a[13] & b[234])^(a[12] & b[235])^(a[11] & b[236])^(a[10] & b[237])^(a[9] & b[238])^(a[8] & b[239])^(a[7] & b[240])^(a[6] & b[241])^(a[5] & b[242])^(a[4] & b[243])^(a[3] & b[244])^(a[2] & b[245])^(a[1] & b[246])^(a[0] & b[247]);
assign y[248] = (a[248] & b[0])^(a[247] & b[1])^(a[246] & b[2])^(a[245] & b[3])^(a[244] & b[4])^(a[243] & b[5])^(a[242] & b[6])^(a[241] & b[7])^(a[240] & b[8])^(a[239] & b[9])^(a[238] & b[10])^(a[237] & b[11])^(a[236] & b[12])^(a[235] & b[13])^(a[234] & b[14])^(a[233] & b[15])^(a[232] & b[16])^(a[231] & b[17])^(a[230] & b[18])^(a[229] & b[19])^(a[228] & b[20])^(a[227] & b[21])^(a[226] & b[22])^(a[225] & b[23])^(a[224] & b[24])^(a[223] & b[25])^(a[222] & b[26])^(a[221] & b[27])^(a[220] & b[28])^(a[219] & b[29])^(a[218] & b[30])^(a[217] & b[31])^(a[216] & b[32])^(a[215] & b[33])^(a[214] & b[34])^(a[213] & b[35])^(a[212] & b[36])^(a[211] & b[37])^(a[210] & b[38])^(a[209] & b[39])^(a[208] & b[40])^(a[207] & b[41])^(a[206] & b[42])^(a[205] & b[43])^(a[204] & b[44])^(a[203] & b[45])^(a[202] & b[46])^(a[201] & b[47])^(a[200] & b[48])^(a[199] & b[49])^(a[198] & b[50])^(a[197] & b[51])^(a[196] & b[52])^(a[195] & b[53])^(a[194] & b[54])^(a[193] & b[55])^(a[192] & b[56])^(a[191] & b[57])^(a[190] & b[58])^(a[189] & b[59])^(a[188] & b[60])^(a[187] & b[61])^(a[186] & b[62])^(a[185] & b[63])^(a[184] & b[64])^(a[183] & b[65])^(a[182] & b[66])^(a[181] & b[67])^(a[180] & b[68])^(a[179] & b[69])^(a[178] & b[70])^(a[177] & b[71])^(a[176] & b[72])^(a[175] & b[73])^(a[174] & b[74])^(a[173] & b[75])^(a[172] & b[76])^(a[171] & b[77])^(a[170] & b[78])^(a[169] & b[79])^(a[168] & b[80])^(a[167] & b[81])^(a[166] & b[82])^(a[165] & b[83])^(a[164] & b[84])^(a[163] & b[85])^(a[162] & b[86])^(a[161] & b[87])^(a[160] & b[88])^(a[159] & b[89])^(a[158] & b[90])^(a[157] & b[91])^(a[156] & b[92])^(a[155] & b[93])^(a[154] & b[94])^(a[153] & b[95])^(a[152] & b[96])^(a[151] & b[97])^(a[150] & b[98])^(a[149] & b[99])^(a[148] & b[100])^(a[147] & b[101])^(a[146] & b[102])^(a[145] & b[103])^(a[144] & b[104])^(a[143] & b[105])^(a[142] & b[106])^(a[141] & b[107])^(a[140] & b[108])^(a[139] & b[109])^(a[138] & b[110])^(a[137] & b[111])^(a[136] & b[112])^(a[135] & b[113])^(a[134] & b[114])^(a[133] & b[115])^(a[132] & b[116])^(a[131] & b[117])^(a[130] & b[118])^(a[129] & b[119])^(a[128] & b[120])^(a[127] & b[121])^(a[126] & b[122])^(a[125] & b[123])^(a[124] & b[124])^(a[123] & b[125])^(a[122] & b[126])^(a[121] & b[127])^(a[120] & b[128])^(a[119] & b[129])^(a[118] & b[130])^(a[117] & b[131])^(a[116] & b[132])^(a[115] & b[133])^(a[114] & b[134])^(a[113] & b[135])^(a[112] & b[136])^(a[111] & b[137])^(a[110] & b[138])^(a[109] & b[139])^(a[108] & b[140])^(a[107] & b[141])^(a[106] & b[142])^(a[105] & b[143])^(a[104] & b[144])^(a[103] & b[145])^(a[102] & b[146])^(a[101] & b[147])^(a[100] & b[148])^(a[99] & b[149])^(a[98] & b[150])^(a[97] & b[151])^(a[96] & b[152])^(a[95] & b[153])^(a[94] & b[154])^(a[93] & b[155])^(a[92] & b[156])^(a[91] & b[157])^(a[90] & b[158])^(a[89] & b[159])^(a[88] & b[160])^(a[87] & b[161])^(a[86] & b[162])^(a[85] & b[163])^(a[84] & b[164])^(a[83] & b[165])^(a[82] & b[166])^(a[81] & b[167])^(a[80] & b[168])^(a[79] & b[169])^(a[78] & b[170])^(a[77] & b[171])^(a[76] & b[172])^(a[75] & b[173])^(a[74] & b[174])^(a[73] & b[175])^(a[72] & b[176])^(a[71] & b[177])^(a[70] & b[178])^(a[69] & b[179])^(a[68] & b[180])^(a[67] & b[181])^(a[66] & b[182])^(a[65] & b[183])^(a[64] & b[184])^(a[63] & b[185])^(a[62] & b[186])^(a[61] & b[187])^(a[60] & b[188])^(a[59] & b[189])^(a[58] & b[190])^(a[57] & b[191])^(a[56] & b[192])^(a[55] & b[193])^(a[54] & b[194])^(a[53] & b[195])^(a[52] & b[196])^(a[51] & b[197])^(a[50] & b[198])^(a[49] & b[199])^(a[48] & b[200])^(a[47] & b[201])^(a[46] & b[202])^(a[45] & b[203])^(a[44] & b[204])^(a[43] & b[205])^(a[42] & b[206])^(a[41] & b[207])^(a[40] & b[208])^(a[39] & b[209])^(a[38] & b[210])^(a[37] & b[211])^(a[36] & b[212])^(a[35] & b[213])^(a[34] & b[214])^(a[33] & b[215])^(a[32] & b[216])^(a[31] & b[217])^(a[30] & b[218])^(a[29] & b[219])^(a[28] & b[220])^(a[27] & b[221])^(a[26] & b[222])^(a[25] & b[223])^(a[24] & b[224])^(a[23] & b[225])^(a[22] & b[226])^(a[21] & b[227])^(a[20] & b[228])^(a[19] & b[229])^(a[18] & b[230])^(a[17] & b[231])^(a[16] & b[232])^(a[15] & b[233])^(a[14] & b[234])^(a[13] & b[235])^(a[12] & b[236])^(a[11] & b[237])^(a[10] & b[238])^(a[9] & b[239])^(a[8] & b[240])^(a[7] & b[241])^(a[6] & b[242])^(a[5] & b[243])^(a[4] & b[244])^(a[3] & b[245])^(a[2] & b[246])^(a[1] & b[247])^(a[0] & b[248]);
assign y[249] = (a[249] & b[0])^(a[248] & b[1])^(a[247] & b[2])^(a[246] & b[3])^(a[245] & b[4])^(a[244] & b[5])^(a[243] & b[6])^(a[242] & b[7])^(a[241] & b[8])^(a[240] & b[9])^(a[239] & b[10])^(a[238] & b[11])^(a[237] & b[12])^(a[236] & b[13])^(a[235] & b[14])^(a[234] & b[15])^(a[233] & b[16])^(a[232] & b[17])^(a[231] & b[18])^(a[230] & b[19])^(a[229] & b[20])^(a[228] & b[21])^(a[227] & b[22])^(a[226] & b[23])^(a[225] & b[24])^(a[224] & b[25])^(a[223] & b[26])^(a[222] & b[27])^(a[221] & b[28])^(a[220] & b[29])^(a[219] & b[30])^(a[218] & b[31])^(a[217] & b[32])^(a[216] & b[33])^(a[215] & b[34])^(a[214] & b[35])^(a[213] & b[36])^(a[212] & b[37])^(a[211] & b[38])^(a[210] & b[39])^(a[209] & b[40])^(a[208] & b[41])^(a[207] & b[42])^(a[206] & b[43])^(a[205] & b[44])^(a[204] & b[45])^(a[203] & b[46])^(a[202] & b[47])^(a[201] & b[48])^(a[200] & b[49])^(a[199] & b[50])^(a[198] & b[51])^(a[197] & b[52])^(a[196] & b[53])^(a[195] & b[54])^(a[194] & b[55])^(a[193] & b[56])^(a[192] & b[57])^(a[191] & b[58])^(a[190] & b[59])^(a[189] & b[60])^(a[188] & b[61])^(a[187] & b[62])^(a[186] & b[63])^(a[185] & b[64])^(a[184] & b[65])^(a[183] & b[66])^(a[182] & b[67])^(a[181] & b[68])^(a[180] & b[69])^(a[179] & b[70])^(a[178] & b[71])^(a[177] & b[72])^(a[176] & b[73])^(a[175] & b[74])^(a[174] & b[75])^(a[173] & b[76])^(a[172] & b[77])^(a[171] & b[78])^(a[170] & b[79])^(a[169] & b[80])^(a[168] & b[81])^(a[167] & b[82])^(a[166] & b[83])^(a[165] & b[84])^(a[164] & b[85])^(a[163] & b[86])^(a[162] & b[87])^(a[161] & b[88])^(a[160] & b[89])^(a[159] & b[90])^(a[158] & b[91])^(a[157] & b[92])^(a[156] & b[93])^(a[155] & b[94])^(a[154] & b[95])^(a[153] & b[96])^(a[152] & b[97])^(a[151] & b[98])^(a[150] & b[99])^(a[149] & b[100])^(a[148] & b[101])^(a[147] & b[102])^(a[146] & b[103])^(a[145] & b[104])^(a[144] & b[105])^(a[143] & b[106])^(a[142] & b[107])^(a[141] & b[108])^(a[140] & b[109])^(a[139] & b[110])^(a[138] & b[111])^(a[137] & b[112])^(a[136] & b[113])^(a[135] & b[114])^(a[134] & b[115])^(a[133] & b[116])^(a[132] & b[117])^(a[131] & b[118])^(a[130] & b[119])^(a[129] & b[120])^(a[128] & b[121])^(a[127] & b[122])^(a[126] & b[123])^(a[125] & b[124])^(a[124] & b[125])^(a[123] & b[126])^(a[122] & b[127])^(a[121] & b[128])^(a[120] & b[129])^(a[119] & b[130])^(a[118] & b[131])^(a[117] & b[132])^(a[116] & b[133])^(a[115] & b[134])^(a[114] & b[135])^(a[113] & b[136])^(a[112] & b[137])^(a[111] & b[138])^(a[110] & b[139])^(a[109] & b[140])^(a[108] & b[141])^(a[107] & b[142])^(a[106] & b[143])^(a[105] & b[144])^(a[104] & b[145])^(a[103] & b[146])^(a[102] & b[147])^(a[101] & b[148])^(a[100] & b[149])^(a[99] & b[150])^(a[98] & b[151])^(a[97] & b[152])^(a[96] & b[153])^(a[95] & b[154])^(a[94] & b[155])^(a[93] & b[156])^(a[92] & b[157])^(a[91] & b[158])^(a[90] & b[159])^(a[89] & b[160])^(a[88] & b[161])^(a[87] & b[162])^(a[86] & b[163])^(a[85] & b[164])^(a[84] & b[165])^(a[83] & b[166])^(a[82] & b[167])^(a[81] & b[168])^(a[80] & b[169])^(a[79] & b[170])^(a[78] & b[171])^(a[77] & b[172])^(a[76] & b[173])^(a[75] & b[174])^(a[74] & b[175])^(a[73] & b[176])^(a[72] & b[177])^(a[71] & b[178])^(a[70] & b[179])^(a[69] & b[180])^(a[68] & b[181])^(a[67] & b[182])^(a[66] & b[183])^(a[65] & b[184])^(a[64] & b[185])^(a[63] & b[186])^(a[62] & b[187])^(a[61] & b[188])^(a[60] & b[189])^(a[59] & b[190])^(a[58] & b[191])^(a[57] & b[192])^(a[56] & b[193])^(a[55] & b[194])^(a[54] & b[195])^(a[53] & b[196])^(a[52] & b[197])^(a[51] & b[198])^(a[50] & b[199])^(a[49] & b[200])^(a[48] & b[201])^(a[47] & b[202])^(a[46] & b[203])^(a[45] & b[204])^(a[44] & b[205])^(a[43] & b[206])^(a[42] & b[207])^(a[41] & b[208])^(a[40] & b[209])^(a[39] & b[210])^(a[38] & b[211])^(a[37] & b[212])^(a[36] & b[213])^(a[35] & b[214])^(a[34] & b[215])^(a[33] & b[216])^(a[32] & b[217])^(a[31] & b[218])^(a[30] & b[219])^(a[29] & b[220])^(a[28] & b[221])^(a[27] & b[222])^(a[26] & b[223])^(a[25] & b[224])^(a[24] & b[225])^(a[23] & b[226])^(a[22] & b[227])^(a[21] & b[228])^(a[20] & b[229])^(a[19] & b[230])^(a[18] & b[231])^(a[17] & b[232])^(a[16] & b[233])^(a[15] & b[234])^(a[14] & b[235])^(a[13] & b[236])^(a[12] & b[237])^(a[11] & b[238])^(a[10] & b[239])^(a[9] & b[240])^(a[8] & b[241])^(a[7] & b[242])^(a[6] & b[243])^(a[5] & b[244])^(a[4] & b[245])^(a[3] & b[246])^(a[2] & b[247])^(a[1] & b[248])^(a[0] & b[249]);
assign y[250] = (a[250] & b[0])^(a[249] & b[1])^(a[248] & b[2])^(a[247] & b[3])^(a[246] & b[4])^(a[245] & b[5])^(a[244] & b[6])^(a[243] & b[7])^(a[242] & b[8])^(a[241] & b[9])^(a[240] & b[10])^(a[239] & b[11])^(a[238] & b[12])^(a[237] & b[13])^(a[236] & b[14])^(a[235] & b[15])^(a[234] & b[16])^(a[233] & b[17])^(a[232] & b[18])^(a[231] & b[19])^(a[230] & b[20])^(a[229] & b[21])^(a[228] & b[22])^(a[227] & b[23])^(a[226] & b[24])^(a[225] & b[25])^(a[224] & b[26])^(a[223] & b[27])^(a[222] & b[28])^(a[221] & b[29])^(a[220] & b[30])^(a[219] & b[31])^(a[218] & b[32])^(a[217] & b[33])^(a[216] & b[34])^(a[215] & b[35])^(a[214] & b[36])^(a[213] & b[37])^(a[212] & b[38])^(a[211] & b[39])^(a[210] & b[40])^(a[209] & b[41])^(a[208] & b[42])^(a[207] & b[43])^(a[206] & b[44])^(a[205] & b[45])^(a[204] & b[46])^(a[203] & b[47])^(a[202] & b[48])^(a[201] & b[49])^(a[200] & b[50])^(a[199] & b[51])^(a[198] & b[52])^(a[197] & b[53])^(a[196] & b[54])^(a[195] & b[55])^(a[194] & b[56])^(a[193] & b[57])^(a[192] & b[58])^(a[191] & b[59])^(a[190] & b[60])^(a[189] & b[61])^(a[188] & b[62])^(a[187] & b[63])^(a[186] & b[64])^(a[185] & b[65])^(a[184] & b[66])^(a[183] & b[67])^(a[182] & b[68])^(a[181] & b[69])^(a[180] & b[70])^(a[179] & b[71])^(a[178] & b[72])^(a[177] & b[73])^(a[176] & b[74])^(a[175] & b[75])^(a[174] & b[76])^(a[173] & b[77])^(a[172] & b[78])^(a[171] & b[79])^(a[170] & b[80])^(a[169] & b[81])^(a[168] & b[82])^(a[167] & b[83])^(a[166] & b[84])^(a[165] & b[85])^(a[164] & b[86])^(a[163] & b[87])^(a[162] & b[88])^(a[161] & b[89])^(a[160] & b[90])^(a[159] & b[91])^(a[158] & b[92])^(a[157] & b[93])^(a[156] & b[94])^(a[155] & b[95])^(a[154] & b[96])^(a[153] & b[97])^(a[152] & b[98])^(a[151] & b[99])^(a[150] & b[100])^(a[149] & b[101])^(a[148] & b[102])^(a[147] & b[103])^(a[146] & b[104])^(a[145] & b[105])^(a[144] & b[106])^(a[143] & b[107])^(a[142] & b[108])^(a[141] & b[109])^(a[140] & b[110])^(a[139] & b[111])^(a[138] & b[112])^(a[137] & b[113])^(a[136] & b[114])^(a[135] & b[115])^(a[134] & b[116])^(a[133] & b[117])^(a[132] & b[118])^(a[131] & b[119])^(a[130] & b[120])^(a[129] & b[121])^(a[128] & b[122])^(a[127] & b[123])^(a[126] & b[124])^(a[125] & b[125])^(a[124] & b[126])^(a[123] & b[127])^(a[122] & b[128])^(a[121] & b[129])^(a[120] & b[130])^(a[119] & b[131])^(a[118] & b[132])^(a[117] & b[133])^(a[116] & b[134])^(a[115] & b[135])^(a[114] & b[136])^(a[113] & b[137])^(a[112] & b[138])^(a[111] & b[139])^(a[110] & b[140])^(a[109] & b[141])^(a[108] & b[142])^(a[107] & b[143])^(a[106] & b[144])^(a[105] & b[145])^(a[104] & b[146])^(a[103] & b[147])^(a[102] & b[148])^(a[101] & b[149])^(a[100] & b[150])^(a[99] & b[151])^(a[98] & b[152])^(a[97] & b[153])^(a[96] & b[154])^(a[95] & b[155])^(a[94] & b[156])^(a[93] & b[157])^(a[92] & b[158])^(a[91] & b[159])^(a[90] & b[160])^(a[89] & b[161])^(a[88] & b[162])^(a[87] & b[163])^(a[86] & b[164])^(a[85] & b[165])^(a[84] & b[166])^(a[83] & b[167])^(a[82] & b[168])^(a[81] & b[169])^(a[80] & b[170])^(a[79] & b[171])^(a[78] & b[172])^(a[77] & b[173])^(a[76] & b[174])^(a[75] & b[175])^(a[74] & b[176])^(a[73] & b[177])^(a[72] & b[178])^(a[71] & b[179])^(a[70] & b[180])^(a[69] & b[181])^(a[68] & b[182])^(a[67] & b[183])^(a[66] & b[184])^(a[65] & b[185])^(a[64] & b[186])^(a[63] & b[187])^(a[62] & b[188])^(a[61] & b[189])^(a[60] & b[190])^(a[59] & b[191])^(a[58] & b[192])^(a[57] & b[193])^(a[56] & b[194])^(a[55] & b[195])^(a[54] & b[196])^(a[53] & b[197])^(a[52] & b[198])^(a[51] & b[199])^(a[50] & b[200])^(a[49] & b[201])^(a[48] & b[202])^(a[47] & b[203])^(a[46] & b[204])^(a[45] & b[205])^(a[44] & b[206])^(a[43] & b[207])^(a[42] & b[208])^(a[41] & b[209])^(a[40] & b[210])^(a[39] & b[211])^(a[38] & b[212])^(a[37] & b[213])^(a[36] & b[214])^(a[35] & b[215])^(a[34] & b[216])^(a[33] & b[217])^(a[32] & b[218])^(a[31] & b[219])^(a[30] & b[220])^(a[29] & b[221])^(a[28] & b[222])^(a[27] & b[223])^(a[26] & b[224])^(a[25] & b[225])^(a[24] & b[226])^(a[23] & b[227])^(a[22] & b[228])^(a[21] & b[229])^(a[20] & b[230])^(a[19] & b[231])^(a[18] & b[232])^(a[17] & b[233])^(a[16] & b[234])^(a[15] & b[235])^(a[14] & b[236])^(a[13] & b[237])^(a[12] & b[238])^(a[11] & b[239])^(a[10] & b[240])^(a[9] & b[241])^(a[8] & b[242])^(a[7] & b[243])^(a[6] & b[244])^(a[5] & b[245])^(a[4] & b[246])^(a[3] & b[247])^(a[2] & b[248])^(a[1] & b[249])^(a[0] & b[250]);
assign y[251] = (a[251] & b[0])^(a[250] & b[1])^(a[249] & b[2])^(a[248] & b[3])^(a[247] & b[4])^(a[246] & b[5])^(a[245] & b[6])^(a[244] & b[7])^(a[243] & b[8])^(a[242] & b[9])^(a[241] & b[10])^(a[240] & b[11])^(a[239] & b[12])^(a[238] & b[13])^(a[237] & b[14])^(a[236] & b[15])^(a[235] & b[16])^(a[234] & b[17])^(a[233] & b[18])^(a[232] & b[19])^(a[231] & b[20])^(a[230] & b[21])^(a[229] & b[22])^(a[228] & b[23])^(a[227] & b[24])^(a[226] & b[25])^(a[225] & b[26])^(a[224] & b[27])^(a[223] & b[28])^(a[222] & b[29])^(a[221] & b[30])^(a[220] & b[31])^(a[219] & b[32])^(a[218] & b[33])^(a[217] & b[34])^(a[216] & b[35])^(a[215] & b[36])^(a[214] & b[37])^(a[213] & b[38])^(a[212] & b[39])^(a[211] & b[40])^(a[210] & b[41])^(a[209] & b[42])^(a[208] & b[43])^(a[207] & b[44])^(a[206] & b[45])^(a[205] & b[46])^(a[204] & b[47])^(a[203] & b[48])^(a[202] & b[49])^(a[201] & b[50])^(a[200] & b[51])^(a[199] & b[52])^(a[198] & b[53])^(a[197] & b[54])^(a[196] & b[55])^(a[195] & b[56])^(a[194] & b[57])^(a[193] & b[58])^(a[192] & b[59])^(a[191] & b[60])^(a[190] & b[61])^(a[189] & b[62])^(a[188] & b[63])^(a[187] & b[64])^(a[186] & b[65])^(a[185] & b[66])^(a[184] & b[67])^(a[183] & b[68])^(a[182] & b[69])^(a[181] & b[70])^(a[180] & b[71])^(a[179] & b[72])^(a[178] & b[73])^(a[177] & b[74])^(a[176] & b[75])^(a[175] & b[76])^(a[174] & b[77])^(a[173] & b[78])^(a[172] & b[79])^(a[171] & b[80])^(a[170] & b[81])^(a[169] & b[82])^(a[168] & b[83])^(a[167] & b[84])^(a[166] & b[85])^(a[165] & b[86])^(a[164] & b[87])^(a[163] & b[88])^(a[162] & b[89])^(a[161] & b[90])^(a[160] & b[91])^(a[159] & b[92])^(a[158] & b[93])^(a[157] & b[94])^(a[156] & b[95])^(a[155] & b[96])^(a[154] & b[97])^(a[153] & b[98])^(a[152] & b[99])^(a[151] & b[100])^(a[150] & b[101])^(a[149] & b[102])^(a[148] & b[103])^(a[147] & b[104])^(a[146] & b[105])^(a[145] & b[106])^(a[144] & b[107])^(a[143] & b[108])^(a[142] & b[109])^(a[141] & b[110])^(a[140] & b[111])^(a[139] & b[112])^(a[138] & b[113])^(a[137] & b[114])^(a[136] & b[115])^(a[135] & b[116])^(a[134] & b[117])^(a[133] & b[118])^(a[132] & b[119])^(a[131] & b[120])^(a[130] & b[121])^(a[129] & b[122])^(a[128] & b[123])^(a[127] & b[124])^(a[126] & b[125])^(a[125] & b[126])^(a[124] & b[127])^(a[123] & b[128])^(a[122] & b[129])^(a[121] & b[130])^(a[120] & b[131])^(a[119] & b[132])^(a[118] & b[133])^(a[117] & b[134])^(a[116] & b[135])^(a[115] & b[136])^(a[114] & b[137])^(a[113] & b[138])^(a[112] & b[139])^(a[111] & b[140])^(a[110] & b[141])^(a[109] & b[142])^(a[108] & b[143])^(a[107] & b[144])^(a[106] & b[145])^(a[105] & b[146])^(a[104] & b[147])^(a[103] & b[148])^(a[102] & b[149])^(a[101] & b[150])^(a[100] & b[151])^(a[99] & b[152])^(a[98] & b[153])^(a[97] & b[154])^(a[96] & b[155])^(a[95] & b[156])^(a[94] & b[157])^(a[93] & b[158])^(a[92] & b[159])^(a[91] & b[160])^(a[90] & b[161])^(a[89] & b[162])^(a[88] & b[163])^(a[87] & b[164])^(a[86] & b[165])^(a[85] & b[166])^(a[84] & b[167])^(a[83] & b[168])^(a[82] & b[169])^(a[81] & b[170])^(a[80] & b[171])^(a[79] & b[172])^(a[78] & b[173])^(a[77] & b[174])^(a[76] & b[175])^(a[75] & b[176])^(a[74] & b[177])^(a[73] & b[178])^(a[72] & b[179])^(a[71] & b[180])^(a[70] & b[181])^(a[69] & b[182])^(a[68] & b[183])^(a[67] & b[184])^(a[66] & b[185])^(a[65] & b[186])^(a[64] & b[187])^(a[63] & b[188])^(a[62] & b[189])^(a[61] & b[190])^(a[60] & b[191])^(a[59] & b[192])^(a[58] & b[193])^(a[57] & b[194])^(a[56] & b[195])^(a[55] & b[196])^(a[54] & b[197])^(a[53] & b[198])^(a[52] & b[199])^(a[51] & b[200])^(a[50] & b[201])^(a[49] & b[202])^(a[48] & b[203])^(a[47] & b[204])^(a[46] & b[205])^(a[45] & b[206])^(a[44] & b[207])^(a[43] & b[208])^(a[42] & b[209])^(a[41] & b[210])^(a[40] & b[211])^(a[39] & b[212])^(a[38] & b[213])^(a[37] & b[214])^(a[36] & b[215])^(a[35] & b[216])^(a[34] & b[217])^(a[33] & b[218])^(a[32] & b[219])^(a[31] & b[220])^(a[30] & b[221])^(a[29] & b[222])^(a[28] & b[223])^(a[27] & b[224])^(a[26] & b[225])^(a[25] & b[226])^(a[24] & b[227])^(a[23] & b[228])^(a[22] & b[229])^(a[21] & b[230])^(a[20] & b[231])^(a[19] & b[232])^(a[18] & b[233])^(a[17] & b[234])^(a[16] & b[235])^(a[15] & b[236])^(a[14] & b[237])^(a[13] & b[238])^(a[12] & b[239])^(a[11] & b[240])^(a[10] & b[241])^(a[9] & b[242])^(a[8] & b[243])^(a[7] & b[244])^(a[6] & b[245])^(a[5] & b[246])^(a[4] & b[247])^(a[3] & b[248])^(a[2] & b[249])^(a[1] & b[250])^(a[0] & b[251]);
assign y[252] = (a[252] & b[0])^(a[251] & b[1])^(a[250] & b[2])^(a[249] & b[3])^(a[248] & b[4])^(a[247] & b[5])^(a[246] & b[6])^(a[245] & b[7])^(a[244] & b[8])^(a[243] & b[9])^(a[242] & b[10])^(a[241] & b[11])^(a[240] & b[12])^(a[239] & b[13])^(a[238] & b[14])^(a[237] & b[15])^(a[236] & b[16])^(a[235] & b[17])^(a[234] & b[18])^(a[233] & b[19])^(a[232] & b[20])^(a[231] & b[21])^(a[230] & b[22])^(a[229] & b[23])^(a[228] & b[24])^(a[227] & b[25])^(a[226] & b[26])^(a[225] & b[27])^(a[224] & b[28])^(a[223] & b[29])^(a[222] & b[30])^(a[221] & b[31])^(a[220] & b[32])^(a[219] & b[33])^(a[218] & b[34])^(a[217] & b[35])^(a[216] & b[36])^(a[215] & b[37])^(a[214] & b[38])^(a[213] & b[39])^(a[212] & b[40])^(a[211] & b[41])^(a[210] & b[42])^(a[209] & b[43])^(a[208] & b[44])^(a[207] & b[45])^(a[206] & b[46])^(a[205] & b[47])^(a[204] & b[48])^(a[203] & b[49])^(a[202] & b[50])^(a[201] & b[51])^(a[200] & b[52])^(a[199] & b[53])^(a[198] & b[54])^(a[197] & b[55])^(a[196] & b[56])^(a[195] & b[57])^(a[194] & b[58])^(a[193] & b[59])^(a[192] & b[60])^(a[191] & b[61])^(a[190] & b[62])^(a[189] & b[63])^(a[188] & b[64])^(a[187] & b[65])^(a[186] & b[66])^(a[185] & b[67])^(a[184] & b[68])^(a[183] & b[69])^(a[182] & b[70])^(a[181] & b[71])^(a[180] & b[72])^(a[179] & b[73])^(a[178] & b[74])^(a[177] & b[75])^(a[176] & b[76])^(a[175] & b[77])^(a[174] & b[78])^(a[173] & b[79])^(a[172] & b[80])^(a[171] & b[81])^(a[170] & b[82])^(a[169] & b[83])^(a[168] & b[84])^(a[167] & b[85])^(a[166] & b[86])^(a[165] & b[87])^(a[164] & b[88])^(a[163] & b[89])^(a[162] & b[90])^(a[161] & b[91])^(a[160] & b[92])^(a[159] & b[93])^(a[158] & b[94])^(a[157] & b[95])^(a[156] & b[96])^(a[155] & b[97])^(a[154] & b[98])^(a[153] & b[99])^(a[152] & b[100])^(a[151] & b[101])^(a[150] & b[102])^(a[149] & b[103])^(a[148] & b[104])^(a[147] & b[105])^(a[146] & b[106])^(a[145] & b[107])^(a[144] & b[108])^(a[143] & b[109])^(a[142] & b[110])^(a[141] & b[111])^(a[140] & b[112])^(a[139] & b[113])^(a[138] & b[114])^(a[137] & b[115])^(a[136] & b[116])^(a[135] & b[117])^(a[134] & b[118])^(a[133] & b[119])^(a[132] & b[120])^(a[131] & b[121])^(a[130] & b[122])^(a[129] & b[123])^(a[128] & b[124])^(a[127] & b[125])^(a[126] & b[126])^(a[125] & b[127])^(a[124] & b[128])^(a[123] & b[129])^(a[122] & b[130])^(a[121] & b[131])^(a[120] & b[132])^(a[119] & b[133])^(a[118] & b[134])^(a[117] & b[135])^(a[116] & b[136])^(a[115] & b[137])^(a[114] & b[138])^(a[113] & b[139])^(a[112] & b[140])^(a[111] & b[141])^(a[110] & b[142])^(a[109] & b[143])^(a[108] & b[144])^(a[107] & b[145])^(a[106] & b[146])^(a[105] & b[147])^(a[104] & b[148])^(a[103] & b[149])^(a[102] & b[150])^(a[101] & b[151])^(a[100] & b[152])^(a[99] & b[153])^(a[98] & b[154])^(a[97] & b[155])^(a[96] & b[156])^(a[95] & b[157])^(a[94] & b[158])^(a[93] & b[159])^(a[92] & b[160])^(a[91] & b[161])^(a[90] & b[162])^(a[89] & b[163])^(a[88] & b[164])^(a[87] & b[165])^(a[86] & b[166])^(a[85] & b[167])^(a[84] & b[168])^(a[83] & b[169])^(a[82] & b[170])^(a[81] & b[171])^(a[80] & b[172])^(a[79] & b[173])^(a[78] & b[174])^(a[77] & b[175])^(a[76] & b[176])^(a[75] & b[177])^(a[74] & b[178])^(a[73] & b[179])^(a[72] & b[180])^(a[71] & b[181])^(a[70] & b[182])^(a[69] & b[183])^(a[68] & b[184])^(a[67] & b[185])^(a[66] & b[186])^(a[65] & b[187])^(a[64] & b[188])^(a[63] & b[189])^(a[62] & b[190])^(a[61] & b[191])^(a[60] & b[192])^(a[59] & b[193])^(a[58] & b[194])^(a[57] & b[195])^(a[56] & b[196])^(a[55] & b[197])^(a[54] & b[198])^(a[53] & b[199])^(a[52] & b[200])^(a[51] & b[201])^(a[50] & b[202])^(a[49] & b[203])^(a[48] & b[204])^(a[47] & b[205])^(a[46] & b[206])^(a[45] & b[207])^(a[44] & b[208])^(a[43] & b[209])^(a[42] & b[210])^(a[41] & b[211])^(a[40] & b[212])^(a[39] & b[213])^(a[38] & b[214])^(a[37] & b[215])^(a[36] & b[216])^(a[35] & b[217])^(a[34] & b[218])^(a[33] & b[219])^(a[32] & b[220])^(a[31] & b[221])^(a[30] & b[222])^(a[29] & b[223])^(a[28] & b[224])^(a[27] & b[225])^(a[26] & b[226])^(a[25] & b[227])^(a[24] & b[228])^(a[23] & b[229])^(a[22] & b[230])^(a[21] & b[231])^(a[20] & b[232])^(a[19] & b[233])^(a[18] & b[234])^(a[17] & b[235])^(a[16] & b[236])^(a[15] & b[237])^(a[14] & b[238])^(a[13] & b[239])^(a[12] & b[240])^(a[11] & b[241])^(a[10] & b[242])^(a[9] & b[243])^(a[8] & b[244])^(a[7] & b[245])^(a[6] & b[246])^(a[5] & b[247])^(a[4] & b[248])^(a[3] & b[249])^(a[2] & b[250])^(a[1] & b[251])^(a[0] & b[252]);
assign y[253] = (a[253] & b[0])^(a[252] & b[1])^(a[251] & b[2])^(a[250] & b[3])^(a[249] & b[4])^(a[248] & b[5])^(a[247] & b[6])^(a[246] & b[7])^(a[245] & b[8])^(a[244] & b[9])^(a[243] & b[10])^(a[242] & b[11])^(a[241] & b[12])^(a[240] & b[13])^(a[239] & b[14])^(a[238] & b[15])^(a[237] & b[16])^(a[236] & b[17])^(a[235] & b[18])^(a[234] & b[19])^(a[233] & b[20])^(a[232] & b[21])^(a[231] & b[22])^(a[230] & b[23])^(a[229] & b[24])^(a[228] & b[25])^(a[227] & b[26])^(a[226] & b[27])^(a[225] & b[28])^(a[224] & b[29])^(a[223] & b[30])^(a[222] & b[31])^(a[221] & b[32])^(a[220] & b[33])^(a[219] & b[34])^(a[218] & b[35])^(a[217] & b[36])^(a[216] & b[37])^(a[215] & b[38])^(a[214] & b[39])^(a[213] & b[40])^(a[212] & b[41])^(a[211] & b[42])^(a[210] & b[43])^(a[209] & b[44])^(a[208] & b[45])^(a[207] & b[46])^(a[206] & b[47])^(a[205] & b[48])^(a[204] & b[49])^(a[203] & b[50])^(a[202] & b[51])^(a[201] & b[52])^(a[200] & b[53])^(a[199] & b[54])^(a[198] & b[55])^(a[197] & b[56])^(a[196] & b[57])^(a[195] & b[58])^(a[194] & b[59])^(a[193] & b[60])^(a[192] & b[61])^(a[191] & b[62])^(a[190] & b[63])^(a[189] & b[64])^(a[188] & b[65])^(a[187] & b[66])^(a[186] & b[67])^(a[185] & b[68])^(a[184] & b[69])^(a[183] & b[70])^(a[182] & b[71])^(a[181] & b[72])^(a[180] & b[73])^(a[179] & b[74])^(a[178] & b[75])^(a[177] & b[76])^(a[176] & b[77])^(a[175] & b[78])^(a[174] & b[79])^(a[173] & b[80])^(a[172] & b[81])^(a[171] & b[82])^(a[170] & b[83])^(a[169] & b[84])^(a[168] & b[85])^(a[167] & b[86])^(a[166] & b[87])^(a[165] & b[88])^(a[164] & b[89])^(a[163] & b[90])^(a[162] & b[91])^(a[161] & b[92])^(a[160] & b[93])^(a[159] & b[94])^(a[158] & b[95])^(a[157] & b[96])^(a[156] & b[97])^(a[155] & b[98])^(a[154] & b[99])^(a[153] & b[100])^(a[152] & b[101])^(a[151] & b[102])^(a[150] & b[103])^(a[149] & b[104])^(a[148] & b[105])^(a[147] & b[106])^(a[146] & b[107])^(a[145] & b[108])^(a[144] & b[109])^(a[143] & b[110])^(a[142] & b[111])^(a[141] & b[112])^(a[140] & b[113])^(a[139] & b[114])^(a[138] & b[115])^(a[137] & b[116])^(a[136] & b[117])^(a[135] & b[118])^(a[134] & b[119])^(a[133] & b[120])^(a[132] & b[121])^(a[131] & b[122])^(a[130] & b[123])^(a[129] & b[124])^(a[128] & b[125])^(a[127] & b[126])^(a[126] & b[127])^(a[125] & b[128])^(a[124] & b[129])^(a[123] & b[130])^(a[122] & b[131])^(a[121] & b[132])^(a[120] & b[133])^(a[119] & b[134])^(a[118] & b[135])^(a[117] & b[136])^(a[116] & b[137])^(a[115] & b[138])^(a[114] & b[139])^(a[113] & b[140])^(a[112] & b[141])^(a[111] & b[142])^(a[110] & b[143])^(a[109] & b[144])^(a[108] & b[145])^(a[107] & b[146])^(a[106] & b[147])^(a[105] & b[148])^(a[104] & b[149])^(a[103] & b[150])^(a[102] & b[151])^(a[101] & b[152])^(a[100] & b[153])^(a[99] & b[154])^(a[98] & b[155])^(a[97] & b[156])^(a[96] & b[157])^(a[95] & b[158])^(a[94] & b[159])^(a[93] & b[160])^(a[92] & b[161])^(a[91] & b[162])^(a[90] & b[163])^(a[89] & b[164])^(a[88] & b[165])^(a[87] & b[166])^(a[86] & b[167])^(a[85] & b[168])^(a[84] & b[169])^(a[83] & b[170])^(a[82] & b[171])^(a[81] & b[172])^(a[80] & b[173])^(a[79] & b[174])^(a[78] & b[175])^(a[77] & b[176])^(a[76] & b[177])^(a[75] & b[178])^(a[74] & b[179])^(a[73] & b[180])^(a[72] & b[181])^(a[71] & b[182])^(a[70] & b[183])^(a[69] & b[184])^(a[68] & b[185])^(a[67] & b[186])^(a[66] & b[187])^(a[65] & b[188])^(a[64] & b[189])^(a[63] & b[190])^(a[62] & b[191])^(a[61] & b[192])^(a[60] & b[193])^(a[59] & b[194])^(a[58] & b[195])^(a[57] & b[196])^(a[56] & b[197])^(a[55] & b[198])^(a[54] & b[199])^(a[53] & b[200])^(a[52] & b[201])^(a[51] & b[202])^(a[50] & b[203])^(a[49] & b[204])^(a[48] & b[205])^(a[47] & b[206])^(a[46] & b[207])^(a[45] & b[208])^(a[44] & b[209])^(a[43] & b[210])^(a[42] & b[211])^(a[41] & b[212])^(a[40] & b[213])^(a[39] & b[214])^(a[38] & b[215])^(a[37] & b[216])^(a[36] & b[217])^(a[35] & b[218])^(a[34] & b[219])^(a[33] & b[220])^(a[32] & b[221])^(a[31] & b[222])^(a[30] & b[223])^(a[29] & b[224])^(a[28] & b[225])^(a[27] & b[226])^(a[26] & b[227])^(a[25] & b[228])^(a[24] & b[229])^(a[23] & b[230])^(a[22] & b[231])^(a[21] & b[232])^(a[20] & b[233])^(a[19] & b[234])^(a[18] & b[235])^(a[17] & b[236])^(a[16] & b[237])^(a[15] & b[238])^(a[14] & b[239])^(a[13] & b[240])^(a[12] & b[241])^(a[11] & b[242])^(a[10] & b[243])^(a[9] & b[244])^(a[8] & b[245])^(a[7] & b[246])^(a[6] & b[247])^(a[5] & b[248])^(a[4] & b[249])^(a[3] & b[250])^(a[2] & b[251])^(a[1] & b[252])^(a[0] & b[253]);
assign y[254] = (a[254] & b[0])^(a[253] & b[1])^(a[252] & b[2])^(a[251] & b[3])^(a[250] & b[4])^(a[249] & b[5])^(a[248] & b[6])^(a[247] & b[7])^(a[246] & b[8])^(a[245] & b[9])^(a[244] & b[10])^(a[243] & b[11])^(a[242] & b[12])^(a[241] & b[13])^(a[240] & b[14])^(a[239] & b[15])^(a[238] & b[16])^(a[237] & b[17])^(a[236] & b[18])^(a[235] & b[19])^(a[234] & b[20])^(a[233] & b[21])^(a[232] & b[22])^(a[231] & b[23])^(a[230] & b[24])^(a[229] & b[25])^(a[228] & b[26])^(a[227] & b[27])^(a[226] & b[28])^(a[225] & b[29])^(a[224] & b[30])^(a[223] & b[31])^(a[222] & b[32])^(a[221] & b[33])^(a[220] & b[34])^(a[219] & b[35])^(a[218] & b[36])^(a[217] & b[37])^(a[216] & b[38])^(a[215] & b[39])^(a[214] & b[40])^(a[213] & b[41])^(a[212] & b[42])^(a[211] & b[43])^(a[210] & b[44])^(a[209] & b[45])^(a[208] & b[46])^(a[207] & b[47])^(a[206] & b[48])^(a[205] & b[49])^(a[204] & b[50])^(a[203] & b[51])^(a[202] & b[52])^(a[201] & b[53])^(a[200] & b[54])^(a[199] & b[55])^(a[198] & b[56])^(a[197] & b[57])^(a[196] & b[58])^(a[195] & b[59])^(a[194] & b[60])^(a[193] & b[61])^(a[192] & b[62])^(a[191] & b[63])^(a[190] & b[64])^(a[189] & b[65])^(a[188] & b[66])^(a[187] & b[67])^(a[186] & b[68])^(a[185] & b[69])^(a[184] & b[70])^(a[183] & b[71])^(a[182] & b[72])^(a[181] & b[73])^(a[180] & b[74])^(a[179] & b[75])^(a[178] & b[76])^(a[177] & b[77])^(a[176] & b[78])^(a[175] & b[79])^(a[174] & b[80])^(a[173] & b[81])^(a[172] & b[82])^(a[171] & b[83])^(a[170] & b[84])^(a[169] & b[85])^(a[168] & b[86])^(a[167] & b[87])^(a[166] & b[88])^(a[165] & b[89])^(a[164] & b[90])^(a[163] & b[91])^(a[162] & b[92])^(a[161] & b[93])^(a[160] & b[94])^(a[159] & b[95])^(a[158] & b[96])^(a[157] & b[97])^(a[156] & b[98])^(a[155] & b[99])^(a[154] & b[100])^(a[153] & b[101])^(a[152] & b[102])^(a[151] & b[103])^(a[150] & b[104])^(a[149] & b[105])^(a[148] & b[106])^(a[147] & b[107])^(a[146] & b[108])^(a[145] & b[109])^(a[144] & b[110])^(a[143] & b[111])^(a[142] & b[112])^(a[141] & b[113])^(a[140] & b[114])^(a[139] & b[115])^(a[138] & b[116])^(a[137] & b[117])^(a[136] & b[118])^(a[135] & b[119])^(a[134] & b[120])^(a[133] & b[121])^(a[132] & b[122])^(a[131] & b[123])^(a[130] & b[124])^(a[129] & b[125])^(a[128] & b[126])^(a[127] & b[127])^(a[126] & b[128])^(a[125] & b[129])^(a[124] & b[130])^(a[123] & b[131])^(a[122] & b[132])^(a[121] & b[133])^(a[120] & b[134])^(a[119] & b[135])^(a[118] & b[136])^(a[117] & b[137])^(a[116] & b[138])^(a[115] & b[139])^(a[114] & b[140])^(a[113] & b[141])^(a[112] & b[142])^(a[111] & b[143])^(a[110] & b[144])^(a[109] & b[145])^(a[108] & b[146])^(a[107] & b[147])^(a[106] & b[148])^(a[105] & b[149])^(a[104] & b[150])^(a[103] & b[151])^(a[102] & b[152])^(a[101] & b[153])^(a[100] & b[154])^(a[99] & b[155])^(a[98] & b[156])^(a[97] & b[157])^(a[96] & b[158])^(a[95] & b[159])^(a[94] & b[160])^(a[93] & b[161])^(a[92] & b[162])^(a[91] & b[163])^(a[90] & b[164])^(a[89] & b[165])^(a[88] & b[166])^(a[87] & b[167])^(a[86] & b[168])^(a[85] & b[169])^(a[84] & b[170])^(a[83] & b[171])^(a[82] & b[172])^(a[81] & b[173])^(a[80] & b[174])^(a[79] & b[175])^(a[78] & b[176])^(a[77] & b[177])^(a[76] & b[178])^(a[75] & b[179])^(a[74] & b[180])^(a[73] & b[181])^(a[72] & b[182])^(a[71] & b[183])^(a[70] & b[184])^(a[69] & b[185])^(a[68] & b[186])^(a[67] & b[187])^(a[66] & b[188])^(a[65] & b[189])^(a[64] & b[190])^(a[63] & b[191])^(a[62] & b[192])^(a[61] & b[193])^(a[60] & b[194])^(a[59] & b[195])^(a[58] & b[196])^(a[57] & b[197])^(a[56] & b[198])^(a[55] & b[199])^(a[54] & b[200])^(a[53] & b[201])^(a[52] & b[202])^(a[51] & b[203])^(a[50] & b[204])^(a[49] & b[205])^(a[48] & b[206])^(a[47] & b[207])^(a[46] & b[208])^(a[45] & b[209])^(a[44] & b[210])^(a[43] & b[211])^(a[42] & b[212])^(a[41] & b[213])^(a[40] & b[214])^(a[39] & b[215])^(a[38] & b[216])^(a[37] & b[217])^(a[36] & b[218])^(a[35] & b[219])^(a[34] & b[220])^(a[33] & b[221])^(a[32] & b[222])^(a[31] & b[223])^(a[30] & b[224])^(a[29] & b[225])^(a[28] & b[226])^(a[27] & b[227])^(a[26] & b[228])^(a[25] & b[229])^(a[24] & b[230])^(a[23] & b[231])^(a[22] & b[232])^(a[21] & b[233])^(a[20] & b[234])^(a[19] & b[235])^(a[18] & b[236])^(a[17] & b[237])^(a[16] & b[238])^(a[15] & b[239])^(a[14] & b[240])^(a[13] & b[241])^(a[12] & b[242])^(a[11] & b[243])^(a[10] & b[244])^(a[9] & b[245])^(a[8] & b[246])^(a[7] & b[247])^(a[6] & b[248])^(a[5] & b[249])^(a[4] & b[250])^(a[3] & b[251])^(a[2] & b[252])^(a[1] & b[253])^(a[0] & b[254]);
assign y[255] = (a[255] & b[0])^(a[254] & b[1])^(a[253] & b[2])^(a[252] & b[3])^(a[251] & b[4])^(a[250] & b[5])^(a[249] & b[6])^(a[248] & b[7])^(a[247] & b[8])^(a[246] & b[9])^(a[245] & b[10])^(a[244] & b[11])^(a[243] & b[12])^(a[242] & b[13])^(a[241] & b[14])^(a[240] & b[15])^(a[239] & b[16])^(a[238] & b[17])^(a[237] & b[18])^(a[236] & b[19])^(a[235] & b[20])^(a[234] & b[21])^(a[233] & b[22])^(a[232] & b[23])^(a[231] & b[24])^(a[230] & b[25])^(a[229] & b[26])^(a[228] & b[27])^(a[227] & b[28])^(a[226] & b[29])^(a[225] & b[30])^(a[224] & b[31])^(a[223] & b[32])^(a[222] & b[33])^(a[221] & b[34])^(a[220] & b[35])^(a[219] & b[36])^(a[218] & b[37])^(a[217] & b[38])^(a[216] & b[39])^(a[215] & b[40])^(a[214] & b[41])^(a[213] & b[42])^(a[212] & b[43])^(a[211] & b[44])^(a[210] & b[45])^(a[209] & b[46])^(a[208] & b[47])^(a[207] & b[48])^(a[206] & b[49])^(a[205] & b[50])^(a[204] & b[51])^(a[203] & b[52])^(a[202] & b[53])^(a[201] & b[54])^(a[200] & b[55])^(a[199] & b[56])^(a[198] & b[57])^(a[197] & b[58])^(a[196] & b[59])^(a[195] & b[60])^(a[194] & b[61])^(a[193] & b[62])^(a[192] & b[63])^(a[191] & b[64])^(a[190] & b[65])^(a[189] & b[66])^(a[188] & b[67])^(a[187] & b[68])^(a[186] & b[69])^(a[185] & b[70])^(a[184] & b[71])^(a[183] & b[72])^(a[182] & b[73])^(a[181] & b[74])^(a[180] & b[75])^(a[179] & b[76])^(a[178] & b[77])^(a[177] & b[78])^(a[176] & b[79])^(a[175] & b[80])^(a[174] & b[81])^(a[173] & b[82])^(a[172] & b[83])^(a[171] & b[84])^(a[170] & b[85])^(a[169] & b[86])^(a[168] & b[87])^(a[167] & b[88])^(a[166] & b[89])^(a[165] & b[90])^(a[164] & b[91])^(a[163] & b[92])^(a[162] & b[93])^(a[161] & b[94])^(a[160] & b[95])^(a[159] & b[96])^(a[158] & b[97])^(a[157] & b[98])^(a[156] & b[99])^(a[155] & b[100])^(a[154] & b[101])^(a[153] & b[102])^(a[152] & b[103])^(a[151] & b[104])^(a[150] & b[105])^(a[149] & b[106])^(a[148] & b[107])^(a[147] & b[108])^(a[146] & b[109])^(a[145] & b[110])^(a[144] & b[111])^(a[143] & b[112])^(a[142] & b[113])^(a[141] & b[114])^(a[140] & b[115])^(a[139] & b[116])^(a[138] & b[117])^(a[137] & b[118])^(a[136] & b[119])^(a[135] & b[120])^(a[134] & b[121])^(a[133] & b[122])^(a[132] & b[123])^(a[131] & b[124])^(a[130] & b[125])^(a[129] & b[126])^(a[128] & b[127])^(a[127] & b[128])^(a[126] & b[129])^(a[125] & b[130])^(a[124] & b[131])^(a[123] & b[132])^(a[122] & b[133])^(a[121] & b[134])^(a[120] & b[135])^(a[119] & b[136])^(a[118] & b[137])^(a[117] & b[138])^(a[116] & b[139])^(a[115] & b[140])^(a[114] & b[141])^(a[113] & b[142])^(a[112] & b[143])^(a[111] & b[144])^(a[110] & b[145])^(a[109] & b[146])^(a[108] & b[147])^(a[107] & b[148])^(a[106] & b[149])^(a[105] & b[150])^(a[104] & b[151])^(a[103] & b[152])^(a[102] & b[153])^(a[101] & b[154])^(a[100] & b[155])^(a[99] & b[156])^(a[98] & b[157])^(a[97] & b[158])^(a[96] & b[159])^(a[95] & b[160])^(a[94] & b[161])^(a[93] & b[162])^(a[92] & b[163])^(a[91] & b[164])^(a[90] & b[165])^(a[89] & b[166])^(a[88] & b[167])^(a[87] & b[168])^(a[86] & b[169])^(a[85] & b[170])^(a[84] & b[171])^(a[83] & b[172])^(a[82] & b[173])^(a[81] & b[174])^(a[80] & b[175])^(a[79] & b[176])^(a[78] & b[177])^(a[77] & b[178])^(a[76] & b[179])^(a[75] & b[180])^(a[74] & b[181])^(a[73] & b[182])^(a[72] & b[183])^(a[71] & b[184])^(a[70] & b[185])^(a[69] & b[186])^(a[68] & b[187])^(a[67] & b[188])^(a[66] & b[189])^(a[65] & b[190])^(a[64] & b[191])^(a[63] & b[192])^(a[62] & b[193])^(a[61] & b[194])^(a[60] & b[195])^(a[59] & b[196])^(a[58] & b[197])^(a[57] & b[198])^(a[56] & b[199])^(a[55] & b[200])^(a[54] & b[201])^(a[53] & b[202])^(a[52] & b[203])^(a[51] & b[204])^(a[50] & b[205])^(a[49] & b[206])^(a[48] & b[207])^(a[47] & b[208])^(a[46] & b[209])^(a[45] & b[210])^(a[44] & b[211])^(a[43] & b[212])^(a[42] & b[213])^(a[41] & b[214])^(a[40] & b[215])^(a[39] & b[216])^(a[38] & b[217])^(a[37] & b[218])^(a[36] & b[219])^(a[35] & b[220])^(a[34] & b[221])^(a[33] & b[222])^(a[32] & b[223])^(a[31] & b[224])^(a[30] & b[225])^(a[29] & b[226])^(a[28] & b[227])^(a[27] & b[228])^(a[26] & b[229])^(a[25] & b[230])^(a[24] & b[231])^(a[23] & b[232])^(a[22] & b[233])^(a[21] & b[234])^(a[20] & b[235])^(a[19] & b[236])^(a[18] & b[237])^(a[17] & b[238])^(a[16] & b[239])^(a[15] & b[240])^(a[14] & b[241])^(a[13] & b[242])^(a[12] & b[243])^(a[11] & b[244])^(a[10] & b[245])^(a[9] & b[246])^(a[8] & b[247])^(a[7] & b[248])^(a[6] & b[249])^(a[5] & b[250])^(a[4] & b[251])^(a[3] & b[252])^(a[2] & b[253])^(a[1] & b[254])^(a[0] & b[255]);
assign y[256] = (a[256] & b[0])^(a[255] & b[1])^(a[254] & b[2])^(a[253] & b[3])^(a[252] & b[4])^(a[251] & b[5])^(a[250] & b[6])^(a[249] & b[7])^(a[248] & b[8])^(a[247] & b[9])^(a[246] & b[10])^(a[245] & b[11])^(a[244] & b[12])^(a[243] & b[13])^(a[242] & b[14])^(a[241] & b[15])^(a[240] & b[16])^(a[239] & b[17])^(a[238] & b[18])^(a[237] & b[19])^(a[236] & b[20])^(a[235] & b[21])^(a[234] & b[22])^(a[233] & b[23])^(a[232] & b[24])^(a[231] & b[25])^(a[230] & b[26])^(a[229] & b[27])^(a[228] & b[28])^(a[227] & b[29])^(a[226] & b[30])^(a[225] & b[31])^(a[224] & b[32])^(a[223] & b[33])^(a[222] & b[34])^(a[221] & b[35])^(a[220] & b[36])^(a[219] & b[37])^(a[218] & b[38])^(a[217] & b[39])^(a[216] & b[40])^(a[215] & b[41])^(a[214] & b[42])^(a[213] & b[43])^(a[212] & b[44])^(a[211] & b[45])^(a[210] & b[46])^(a[209] & b[47])^(a[208] & b[48])^(a[207] & b[49])^(a[206] & b[50])^(a[205] & b[51])^(a[204] & b[52])^(a[203] & b[53])^(a[202] & b[54])^(a[201] & b[55])^(a[200] & b[56])^(a[199] & b[57])^(a[198] & b[58])^(a[197] & b[59])^(a[196] & b[60])^(a[195] & b[61])^(a[194] & b[62])^(a[193] & b[63])^(a[192] & b[64])^(a[191] & b[65])^(a[190] & b[66])^(a[189] & b[67])^(a[188] & b[68])^(a[187] & b[69])^(a[186] & b[70])^(a[185] & b[71])^(a[184] & b[72])^(a[183] & b[73])^(a[182] & b[74])^(a[181] & b[75])^(a[180] & b[76])^(a[179] & b[77])^(a[178] & b[78])^(a[177] & b[79])^(a[176] & b[80])^(a[175] & b[81])^(a[174] & b[82])^(a[173] & b[83])^(a[172] & b[84])^(a[171] & b[85])^(a[170] & b[86])^(a[169] & b[87])^(a[168] & b[88])^(a[167] & b[89])^(a[166] & b[90])^(a[165] & b[91])^(a[164] & b[92])^(a[163] & b[93])^(a[162] & b[94])^(a[161] & b[95])^(a[160] & b[96])^(a[159] & b[97])^(a[158] & b[98])^(a[157] & b[99])^(a[156] & b[100])^(a[155] & b[101])^(a[154] & b[102])^(a[153] & b[103])^(a[152] & b[104])^(a[151] & b[105])^(a[150] & b[106])^(a[149] & b[107])^(a[148] & b[108])^(a[147] & b[109])^(a[146] & b[110])^(a[145] & b[111])^(a[144] & b[112])^(a[143] & b[113])^(a[142] & b[114])^(a[141] & b[115])^(a[140] & b[116])^(a[139] & b[117])^(a[138] & b[118])^(a[137] & b[119])^(a[136] & b[120])^(a[135] & b[121])^(a[134] & b[122])^(a[133] & b[123])^(a[132] & b[124])^(a[131] & b[125])^(a[130] & b[126])^(a[129] & b[127])^(a[128] & b[128])^(a[127] & b[129])^(a[126] & b[130])^(a[125] & b[131])^(a[124] & b[132])^(a[123] & b[133])^(a[122] & b[134])^(a[121] & b[135])^(a[120] & b[136])^(a[119] & b[137])^(a[118] & b[138])^(a[117] & b[139])^(a[116] & b[140])^(a[115] & b[141])^(a[114] & b[142])^(a[113] & b[143])^(a[112] & b[144])^(a[111] & b[145])^(a[110] & b[146])^(a[109] & b[147])^(a[108] & b[148])^(a[107] & b[149])^(a[106] & b[150])^(a[105] & b[151])^(a[104] & b[152])^(a[103] & b[153])^(a[102] & b[154])^(a[101] & b[155])^(a[100] & b[156])^(a[99] & b[157])^(a[98] & b[158])^(a[97] & b[159])^(a[96] & b[160])^(a[95] & b[161])^(a[94] & b[162])^(a[93] & b[163])^(a[92] & b[164])^(a[91] & b[165])^(a[90] & b[166])^(a[89] & b[167])^(a[88] & b[168])^(a[87] & b[169])^(a[86] & b[170])^(a[85] & b[171])^(a[84] & b[172])^(a[83] & b[173])^(a[82] & b[174])^(a[81] & b[175])^(a[80] & b[176])^(a[79] & b[177])^(a[78] & b[178])^(a[77] & b[179])^(a[76] & b[180])^(a[75] & b[181])^(a[74] & b[182])^(a[73] & b[183])^(a[72] & b[184])^(a[71] & b[185])^(a[70] & b[186])^(a[69] & b[187])^(a[68] & b[188])^(a[67] & b[189])^(a[66] & b[190])^(a[65] & b[191])^(a[64] & b[192])^(a[63] & b[193])^(a[62] & b[194])^(a[61] & b[195])^(a[60] & b[196])^(a[59] & b[197])^(a[58] & b[198])^(a[57] & b[199])^(a[56] & b[200])^(a[55] & b[201])^(a[54] & b[202])^(a[53] & b[203])^(a[52] & b[204])^(a[51] & b[205])^(a[50] & b[206])^(a[49] & b[207])^(a[48] & b[208])^(a[47] & b[209])^(a[46] & b[210])^(a[45] & b[211])^(a[44] & b[212])^(a[43] & b[213])^(a[42] & b[214])^(a[41] & b[215])^(a[40] & b[216])^(a[39] & b[217])^(a[38] & b[218])^(a[37] & b[219])^(a[36] & b[220])^(a[35] & b[221])^(a[34] & b[222])^(a[33] & b[223])^(a[32] & b[224])^(a[31] & b[225])^(a[30] & b[226])^(a[29] & b[227])^(a[28] & b[228])^(a[27] & b[229])^(a[26] & b[230])^(a[25] & b[231])^(a[24] & b[232])^(a[23] & b[233])^(a[22] & b[234])^(a[21] & b[235])^(a[20] & b[236])^(a[19] & b[237])^(a[18] & b[238])^(a[17] & b[239])^(a[16] & b[240])^(a[15] & b[241])^(a[14] & b[242])^(a[13] & b[243])^(a[12] & b[244])^(a[11] & b[245])^(a[10] & b[246])^(a[9] & b[247])^(a[8] & b[248])^(a[7] & b[249])^(a[6] & b[250])^(a[5] & b[251])^(a[4] & b[252])^(a[3] & b[253])^(a[2] & b[254])^(a[1] & b[255])^(a[0] & b[256]);
assign y[257] = (a[257] & b[0])^(a[256] & b[1])^(a[255] & b[2])^(a[254] & b[3])^(a[253] & b[4])^(a[252] & b[5])^(a[251] & b[6])^(a[250] & b[7])^(a[249] & b[8])^(a[248] & b[9])^(a[247] & b[10])^(a[246] & b[11])^(a[245] & b[12])^(a[244] & b[13])^(a[243] & b[14])^(a[242] & b[15])^(a[241] & b[16])^(a[240] & b[17])^(a[239] & b[18])^(a[238] & b[19])^(a[237] & b[20])^(a[236] & b[21])^(a[235] & b[22])^(a[234] & b[23])^(a[233] & b[24])^(a[232] & b[25])^(a[231] & b[26])^(a[230] & b[27])^(a[229] & b[28])^(a[228] & b[29])^(a[227] & b[30])^(a[226] & b[31])^(a[225] & b[32])^(a[224] & b[33])^(a[223] & b[34])^(a[222] & b[35])^(a[221] & b[36])^(a[220] & b[37])^(a[219] & b[38])^(a[218] & b[39])^(a[217] & b[40])^(a[216] & b[41])^(a[215] & b[42])^(a[214] & b[43])^(a[213] & b[44])^(a[212] & b[45])^(a[211] & b[46])^(a[210] & b[47])^(a[209] & b[48])^(a[208] & b[49])^(a[207] & b[50])^(a[206] & b[51])^(a[205] & b[52])^(a[204] & b[53])^(a[203] & b[54])^(a[202] & b[55])^(a[201] & b[56])^(a[200] & b[57])^(a[199] & b[58])^(a[198] & b[59])^(a[197] & b[60])^(a[196] & b[61])^(a[195] & b[62])^(a[194] & b[63])^(a[193] & b[64])^(a[192] & b[65])^(a[191] & b[66])^(a[190] & b[67])^(a[189] & b[68])^(a[188] & b[69])^(a[187] & b[70])^(a[186] & b[71])^(a[185] & b[72])^(a[184] & b[73])^(a[183] & b[74])^(a[182] & b[75])^(a[181] & b[76])^(a[180] & b[77])^(a[179] & b[78])^(a[178] & b[79])^(a[177] & b[80])^(a[176] & b[81])^(a[175] & b[82])^(a[174] & b[83])^(a[173] & b[84])^(a[172] & b[85])^(a[171] & b[86])^(a[170] & b[87])^(a[169] & b[88])^(a[168] & b[89])^(a[167] & b[90])^(a[166] & b[91])^(a[165] & b[92])^(a[164] & b[93])^(a[163] & b[94])^(a[162] & b[95])^(a[161] & b[96])^(a[160] & b[97])^(a[159] & b[98])^(a[158] & b[99])^(a[157] & b[100])^(a[156] & b[101])^(a[155] & b[102])^(a[154] & b[103])^(a[153] & b[104])^(a[152] & b[105])^(a[151] & b[106])^(a[150] & b[107])^(a[149] & b[108])^(a[148] & b[109])^(a[147] & b[110])^(a[146] & b[111])^(a[145] & b[112])^(a[144] & b[113])^(a[143] & b[114])^(a[142] & b[115])^(a[141] & b[116])^(a[140] & b[117])^(a[139] & b[118])^(a[138] & b[119])^(a[137] & b[120])^(a[136] & b[121])^(a[135] & b[122])^(a[134] & b[123])^(a[133] & b[124])^(a[132] & b[125])^(a[131] & b[126])^(a[130] & b[127])^(a[129] & b[128])^(a[128] & b[129])^(a[127] & b[130])^(a[126] & b[131])^(a[125] & b[132])^(a[124] & b[133])^(a[123] & b[134])^(a[122] & b[135])^(a[121] & b[136])^(a[120] & b[137])^(a[119] & b[138])^(a[118] & b[139])^(a[117] & b[140])^(a[116] & b[141])^(a[115] & b[142])^(a[114] & b[143])^(a[113] & b[144])^(a[112] & b[145])^(a[111] & b[146])^(a[110] & b[147])^(a[109] & b[148])^(a[108] & b[149])^(a[107] & b[150])^(a[106] & b[151])^(a[105] & b[152])^(a[104] & b[153])^(a[103] & b[154])^(a[102] & b[155])^(a[101] & b[156])^(a[100] & b[157])^(a[99] & b[158])^(a[98] & b[159])^(a[97] & b[160])^(a[96] & b[161])^(a[95] & b[162])^(a[94] & b[163])^(a[93] & b[164])^(a[92] & b[165])^(a[91] & b[166])^(a[90] & b[167])^(a[89] & b[168])^(a[88] & b[169])^(a[87] & b[170])^(a[86] & b[171])^(a[85] & b[172])^(a[84] & b[173])^(a[83] & b[174])^(a[82] & b[175])^(a[81] & b[176])^(a[80] & b[177])^(a[79] & b[178])^(a[78] & b[179])^(a[77] & b[180])^(a[76] & b[181])^(a[75] & b[182])^(a[74] & b[183])^(a[73] & b[184])^(a[72] & b[185])^(a[71] & b[186])^(a[70] & b[187])^(a[69] & b[188])^(a[68] & b[189])^(a[67] & b[190])^(a[66] & b[191])^(a[65] & b[192])^(a[64] & b[193])^(a[63] & b[194])^(a[62] & b[195])^(a[61] & b[196])^(a[60] & b[197])^(a[59] & b[198])^(a[58] & b[199])^(a[57] & b[200])^(a[56] & b[201])^(a[55] & b[202])^(a[54] & b[203])^(a[53] & b[204])^(a[52] & b[205])^(a[51] & b[206])^(a[50] & b[207])^(a[49] & b[208])^(a[48] & b[209])^(a[47] & b[210])^(a[46] & b[211])^(a[45] & b[212])^(a[44] & b[213])^(a[43] & b[214])^(a[42] & b[215])^(a[41] & b[216])^(a[40] & b[217])^(a[39] & b[218])^(a[38] & b[219])^(a[37] & b[220])^(a[36] & b[221])^(a[35] & b[222])^(a[34] & b[223])^(a[33] & b[224])^(a[32] & b[225])^(a[31] & b[226])^(a[30] & b[227])^(a[29] & b[228])^(a[28] & b[229])^(a[27] & b[230])^(a[26] & b[231])^(a[25] & b[232])^(a[24] & b[233])^(a[23] & b[234])^(a[22] & b[235])^(a[21] & b[236])^(a[20] & b[237])^(a[19] & b[238])^(a[18] & b[239])^(a[17] & b[240])^(a[16] & b[241])^(a[15] & b[242])^(a[14] & b[243])^(a[13] & b[244])^(a[12] & b[245])^(a[11] & b[246])^(a[10] & b[247])^(a[9] & b[248])^(a[8] & b[249])^(a[7] & b[250])^(a[6] & b[251])^(a[5] & b[252])^(a[4] & b[253])^(a[3] & b[254])^(a[2] & b[255])^(a[1] & b[256])^(a[0] & b[257]);
assign y[258] = (a[258] & b[0])^(a[257] & b[1])^(a[256] & b[2])^(a[255] & b[3])^(a[254] & b[4])^(a[253] & b[5])^(a[252] & b[6])^(a[251] & b[7])^(a[250] & b[8])^(a[249] & b[9])^(a[248] & b[10])^(a[247] & b[11])^(a[246] & b[12])^(a[245] & b[13])^(a[244] & b[14])^(a[243] & b[15])^(a[242] & b[16])^(a[241] & b[17])^(a[240] & b[18])^(a[239] & b[19])^(a[238] & b[20])^(a[237] & b[21])^(a[236] & b[22])^(a[235] & b[23])^(a[234] & b[24])^(a[233] & b[25])^(a[232] & b[26])^(a[231] & b[27])^(a[230] & b[28])^(a[229] & b[29])^(a[228] & b[30])^(a[227] & b[31])^(a[226] & b[32])^(a[225] & b[33])^(a[224] & b[34])^(a[223] & b[35])^(a[222] & b[36])^(a[221] & b[37])^(a[220] & b[38])^(a[219] & b[39])^(a[218] & b[40])^(a[217] & b[41])^(a[216] & b[42])^(a[215] & b[43])^(a[214] & b[44])^(a[213] & b[45])^(a[212] & b[46])^(a[211] & b[47])^(a[210] & b[48])^(a[209] & b[49])^(a[208] & b[50])^(a[207] & b[51])^(a[206] & b[52])^(a[205] & b[53])^(a[204] & b[54])^(a[203] & b[55])^(a[202] & b[56])^(a[201] & b[57])^(a[200] & b[58])^(a[199] & b[59])^(a[198] & b[60])^(a[197] & b[61])^(a[196] & b[62])^(a[195] & b[63])^(a[194] & b[64])^(a[193] & b[65])^(a[192] & b[66])^(a[191] & b[67])^(a[190] & b[68])^(a[189] & b[69])^(a[188] & b[70])^(a[187] & b[71])^(a[186] & b[72])^(a[185] & b[73])^(a[184] & b[74])^(a[183] & b[75])^(a[182] & b[76])^(a[181] & b[77])^(a[180] & b[78])^(a[179] & b[79])^(a[178] & b[80])^(a[177] & b[81])^(a[176] & b[82])^(a[175] & b[83])^(a[174] & b[84])^(a[173] & b[85])^(a[172] & b[86])^(a[171] & b[87])^(a[170] & b[88])^(a[169] & b[89])^(a[168] & b[90])^(a[167] & b[91])^(a[166] & b[92])^(a[165] & b[93])^(a[164] & b[94])^(a[163] & b[95])^(a[162] & b[96])^(a[161] & b[97])^(a[160] & b[98])^(a[159] & b[99])^(a[158] & b[100])^(a[157] & b[101])^(a[156] & b[102])^(a[155] & b[103])^(a[154] & b[104])^(a[153] & b[105])^(a[152] & b[106])^(a[151] & b[107])^(a[150] & b[108])^(a[149] & b[109])^(a[148] & b[110])^(a[147] & b[111])^(a[146] & b[112])^(a[145] & b[113])^(a[144] & b[114])^(a[143] & b[115])^(a[142] & b[116])^(a[141] & b[117])^(a[140] & b[118])^(a[139] & b[119])^(a[138] & b[120])^(a[137] & b[121])^(a[136] & b[122])^(a[135] & b[123])^(a[134] & b[124])^(a[133] & b[125])^(a[132] & b[126])^(a[131] & b[127])^(a[130] & b[128])^(a[129] & b[129])^(a[128] & b[130])^(a[127] & b[131])^(a[126] & b[132])^(a[125] & b[133])^(a[124] & b[134])^(a[123] & b[135])^(a[122] & b[136])^(a[121] & b[137])^(a[120] & b[138])^(a[119] & b[139])^(a[118] & b[140])^(a[117] & b[141])^(a[116] & b[142])^(a[115] & b[143])^(a[114] & b[144])^(a[113] & b[145])^(a[112] & b[146])^(a[111] & b[147])^(a[110] & b[148])^(a[109] & b[149])^(a[108] & b[150])^(a[107] & b[151])^(a[106] & b[152])^(a[105] & b[153])^(a[104] & b[154])^(a[103] & b[155])^(a[102] & b[156])^(a[101] & b[157])^(a[100] & b[158])^(a[99] & b[159])^(a[98] & b[160])^(a[97] & b[161])^(a[96] & b[162])^(a[95] & b[163])^(a[94] & b[164])^(a[93] & b[165])^(a[92] & b[166])^(a[91] & b[167])^(a[90] & b[168])^(a[89] & b[169])^(a[88] & b[170])^(a[87] & b[171])^(a[86] & b[172])^(a[85] & b[173])^(a[84] & b[174])^(a[83] & b[175])^(a[82] & b[176])^(a[81] & b[177])^(a[80] & b[178])^(a[79] & b[179])^(a[78] & b[180])^(a[77] & b[181])^(a[76] & b[182])^(a[75] & b[183])^(a[74] & b[184])^(a[73] & b[185])^(a[72] & b[186])^(a[71] & b[187])^(a[70] & b[188])^(a[69] & b[189])^(a[68] & b[190])^(a[67] & b[191])^(a[66] & b[192])^(a[65] & b[193])^(a[64] & b[194])^(a[63] & b[195])^(a[62] & b[196])^(a[61] & b[197])^(a[60] & b[198])^(a[59] & b[199])^(a[58] & b[200])^(a[57] & b[201])^(a[56] & b[202])^(a[55] & b[203])^(a[54] & b[204])^(a[53] & b[205])^(a[52] & b[206])^(a[51] & b[207])^(a[50] & b[208])^(a[49] & b[209])^(a[48] & b[210])^(a[47] & b[211])^(a[46] & b[212])^(a[45] & b[213])^(a[44] & b[214])^(a[43] & b[215])^(a[42] & b[216])^(a[41] & b[217])^(a[40] & b[218])^(a[39] & b[219])^(a[38] & b[220])^(a[37] & b[221])^(a[36] & b[222])^(a[35] & b[223])^(a[34] & b[224])^(a[33] & b[225])^(a[32] & b[226])^(a[31] & b[227])^(a[30] & b[228])^(a[29] & b[229])^(a[28] & b[230])^(a[27] & b[231])^(a[26] & b[232])^(a[25] & b[233])^(a[24] & b[234])^(a[23] & b[235])^(a[22] & b[236])^(a[21] & b[237])^(a[20] & b[238])^(a[19] & b[239])^(a[18] & b[240])^(a[17] & b[241])^(a[16] & b[242])^(a[15] & b[243])^(a[14] & b[244])^(a[13] & b[245])^(a[12] & b[246])^(a[11] & b[247])^(a[10] & b[248])^(a[9] & b[249])^(a[8] & b[250])^(a[7] & b[251])^(a[6] & b[252])^(a[5] & b[253])^(a[4] & b[254])^(a[3] & b[255])^(a[2] & b[256])^(a[1] & b[257])^(a[0] & b[258]);
assign y[259] = (a[259] & b[0])^(a[258] & b[1])^(a[257] & b[2])^(a[256] & b[3])^(a[255] & b[4])^(a[254] & b[5])^(a[253] & b[6])^(a[252] & b[7])^(a[251] & b[8])^(a[250] & b[9])^(a[249] & b[10])^(a[248] & b[11])^(a[247] & b[12])^(a[246] & b[13])^(a[245] & b[14])^(a[244] & b[15])^(a[243] & b[16])^(a[242] & b[17])^(a[241] & b[18])^(a[240] & b[19])^(a[239] & b[20])^(a[238] & b[21])^(a[237] & b[22])^(a[236] & b[23])^(a[235] & b[24])^(a[234] & b[25])^(a[233] & b[26])^(a[232] & b[27])^(a[231] & b[28])^(a[230] & b[29])^(a[229] & b[30])^(a[228] & b[31])^(a[227] & b[32])^(a[226] & b[33])^(a[225] & b[34])^(a[224] & b[35])^(a[223] & b[36])^(a[222] & b[37])^(a[221] & b[38])^(a[220] & b[39])^(a[219] & b[40])^(a[218] & b[41])^(a[217] & b[42])^(a[216] & b[43])^(a[215] & b[44])^(a[214] & b[45])^(a[213] & b[46])^(a[212] & b[47])^(a[211] & b[48])^(a[210] & b[49])^(a[209] & b[50])^(a[208] & b[51])^(a[207] & b[52])^(a[206] & b[53])^(a[205] & b[54])^(a[204] & b[55])^(a[203] & b[56])^(a[202] & b[57])^(a[201] & b[58])^(a[200] & b[59])^(a[199] & b[60])^(a[198] & b[61])^(a[197] & b[62])^(a[196] & b[63])^(a[195] & b[64])^(a[194] & b[65])^(a[193] & b[66])^(a[192] & b[67])^(a[191] & b[68])^(a[190] & b[69])^(a[189] & b[70])^(a[188] & b[71])^(a[187] & b[72])^(a[186] & b[73])^(a[185] & b[74])^(a[184] & b[75])^(a[183] & b[76])^(a[182] & b[77])^(a[181] & b[78])^(a[180] & b[79])^(a[179] & b[80])^(a[178] & b[81])^(a[177] & b[82])^(a[176] & b[83])^(a[175] & b[84])^(a[174] & b[85])^(a[173] & b[86])^(a[172] & b[87])^(a[171] & b[88])^(a[170] & b[89])^(a[169] & b[90])^(a[168] & b[91])^(a[167] & b[92])^(a[166] & b[93])^(a[165] & b[94])^(a[164] & b[95])^(a[163] & b[96])^(a[162] & b[97])^(a[161] & b[98])^(a[160] & b[99])^(a[159] & b[100])^(a[158] & b[101])^(a[157] & b[102])^(a[156] & b[103])^(a[155] & b[104])^(a[154] & b[105])^(a[153] & b[106])^(a[152] & b[107])^(a[151] & b[108])^(a[150] & b[109])^(a[149] & b[110])^(a[148] & b[111])^(a[147] & b[112])^(a[146] & b[113])^(a[145] & b[114])^(a[144] & b[115])^(a[143] & b[116])^(a[142] & b[117])^(a[141] & b[118])^(a[140] & b[119])^(a[139] & b[120])^(a[138] & b[121])^(a[137] & b[122])^(a[136] & b[123])^(a[135] & b[124])^(a[134] & b[125])^(a[133] & b[126])^(a[132] & b[127])^(a[131] & b[128])^(a[130] & b[129])^(a[129] & b[130])^(a[128] & b[131])^(a[127] & b[132])^(a[126] & b[133])^(a[125] & b[134])^(a[124] & b[135])^(a[123] & b[136])^(a[122] & b[137])^(a[121] & b[138])^(a[120] & b[139])^(a[119] & b[140])^(a[118] & b[141])^(a[117] & b[142])^(a[116] & b[143])^(a[115] & b[144])^(a[114] & b[145])^(a[113] & b[146])^(a[112] & b[147])^(a[111] & b[148])^(a[110] & b[149])^(a[109] & b[150])^(a[108] & b[151])^(a[107] & b[152])^(a[106] & b[153])^(a[105] & b[154])^(a[104] & b[155])^(a[103] & b[156])^(a[102] & b[157])^(a[101] & b[158])^(a[100] & b[159])^(a[99] & b[160])^(a[98] & b[161])^(a[97] & b[162])^(a[96] & b[163])^(a[95] & b[164])^(a[94] & b[165])^(a[93] & b[166])^(a[92] & b[167])^(a[91] & b[168])^(a[90] & b[169])^(a[89] & b[170])^(a[88] & b[171])^(a[87] & b[172])^(a[86] & b[173])^(a[85] & b[174])^(a[84] & b[175])^(a[83] & b[176])^(a[82] & b[177])^(a[81] & b[178])^(a[80] & b[179])^(a[79] & b[180])^(a[78] & b[181])^(a[77] & b[182])^(a[76] & b[183])^(a[75] & b[184])^(a[74] & b[185])^(a[73] & b[186])^(a[72] & b[187])^(a[71] & b[188])^(a[70] & b[189])^(a[69] & b[190])^(a[68] & b[191])^(a[67] & b[192])^(a[66] & b[193])^(a[65] & b[194])^(a[64] & b[195])^(a[63] & b[196])^(a[62] & b[197])^(a[61] & b[198])^(a[60] & b[199])^(a[59] & b[200])^(a[58] & b[201])^(a[57] & b[202])^(a[56] & b[203])^(a[55] & b[204])^(a[54] & b[205])^(a[53] & b[206])^(a[52] & b[207])^(a[51] & b[208])^(a[50] & b[209])^(a[49] & b[210])^(a[48] & b[211])^(a[47] & b[212])^(a[46] & b[213])^(a[45] & b[214])^(a[44] & b[215])^(a[43] & b[216])^(a[42] & b[217])^(a[41] & b[218])^(a[40] & b[219])^(a[39] & b[220])^(a[38] & b[221])^(a[37] & b[222])^(a[36] & b[223])^(a[35] & b[224])^(a[34] & b[225])^(a[33] & b[226])^(a[32] & b[227])^(a[31] & b[228])^(a[30] & b[229])^(a[29] & b[230])^(a[28] & b[231])^(a[27] & b[232])^(a[26] & b[233])^(a[25] & b[234])^(a[24] & b[235])^(a[23] & b[236])^(a[22] & b[237])^(a[21] & b[238])^(a[20] & b[239])^(a[19] & b[240])^(a[18] & b[241])^(a[17] & b[242])^(a[16] & b[243])^(a[15] & b[244])^(a[14] & b[245])^(a[13] & b[246])^(a[12] & b[247])^(a[11] & b[248])^(a[10] & b[249])^(a[9] & b[250])^(a[8] & b[251])^(a[7] & b[252])^(a[6] & b[253])^(a[5] & b[254])^(a[4] & b[255])^(a[3] & b[256])^(a[2] & b[257])^(a[1] & b[258])^(a[0] & b[259]);
assign y[260] = (a[260] & b[0])^(a[259] & b[1])^(a[258] & b[2])^(a[257] & b[3])^(a[256] & b[4])^(a[255] & b[5])^(a[254] & b[6])^(a[253] & b[7])^(a[252] & b[8])^(a[251] & b[9])^(a[250] & b[10])^(a[249] & b[11])^(a[248] & b[12])^(a[247] & b[13])^(a[246] & b[14])^(a[245] & b[15])^(a[244] & b[16])^(a[243] & b[17])^(a[242] & b[18])^(a[241] & b[19])^(a[240] & b[20])^(a[239] & b[21])^(a[238] & b[22])^(a[237] & b[23])^(a[236] & b[24])^(a[235] & b[25])^(a[234] & b[26])^(a[233] & b[27])^(a[232] & b[28])^(a[231] & b[29])^(a[230] & b[30])^(a[229] & b[31])^(a[228] & b[32])^(a[227] & b[33])^(a[226] & b[34])^(a[225] & b[35])^(a[224] & b[36])^(a[223] & b[37])^(a[222] & b[38])^(a[221] & b[39])^(a[220] & b[40])^(a[219] & b[41])^(a[218] & b[42])^(a[217] & b[43])^(a[216] & b[44])^(a[215] & b[45])^(a[214] & b[46])^(a[213] & b[47])^(a[212] & b[48])^(a[211] & b[49])^(a[210] & b[50])^(a[209] & b[51])^(a[208] & b[52])^(a[207] & b[53])^(a[206] & b[54])^(a[205] & b[55])^(a[204] & b[56])^(a[203] & b[57])^(a[202] & b[58])^(a[201] & b[59])^(a[200] & b[60])^(a[199] & b[61])^(a[198] & b[62])^(a[197] & b[63])^(a[196] & b[64])^(a[195] & b[65])^(a[194] & b[66])^(a[193] & b[67])^(a[192] & b[68])^(a[191] & b[69])^(a[190] & b[70])^(a[189] & b[71])^(a[188] & b[72])^(a[187] & b[73])^(a[186] & b[74])^(a[185] & b[75])^(a[184] & b[76])^(a[183] & b[77])^(a[182] & b[78])^(a[181] & b[79])^(a[180] & b[80])^(a[179] & b[81])^(a[178] & b[82])^(a[177] & b[83])^(a[176] & b[84])^(a[175] & b[85])^(a[174] & b[86])^(a[173] & b[87])^(a[172] & b[88])^(a[171] & b[89])^(a[170] & b[90])^(a[169] & b[91])^(a[168] & b[92])^(a[167] & b[93])^(a[166] & b[94])^(a[165] & b[95])^(a[164] & b[96])^(a[163] & b[97])^(a[162] & b[98])^(a[161] & b[99])^(a[160] & b[100])^(a[159] & b[101])^(a[158] & b[102])^(a[157] & b[103])^(a[156] & b[104])^(a[155] & b[105])^(a[154] & b[106])^(a[153] & b[107])^(a[152] & b[108])^(a[151] & b[109])^(a[150] & b[110])^(a[149] & b[111])^(a[148] & b[112])^(a[147] & b[113])^(a[146] & b[114])^(a[145] & b[115])^(a[144] & b[116])^(a[143] & b[117])^(a[142] & b[118])^(a[141] & b[119])^(a[140] & b[120])^(a[139] & b[121])^(a[138] & b[122])^(a[137] & b[123])^(a[136] & b[124])^(a[135] & b[125])^(a[134] & b[126])^(a[133] & b[127])^(a[132] & b[128])^(a[131] & b[129])^(a[130] & b[130])^(a[129] & b[131])^(a[128] & b[132])^(a[127] & b[133])^(a[126] & b[134])^(a[125] & b[135])^(a[124] & b[136])^(a[123] & b[137])^(a[122] & b[138])^(a[121] & b[139])^(a[120] & b[140])^(a[119] & b[141])^(a[118] & b[142])^(a[117] & b[143])^(a[116] & b[144])^(a[115] & b[145])^(a[114] & b[146])^(a[113] & b[147])^(a[112] & b[148])^(a[111] & b[149])^(a[110] & b[150])^(a[109] & b[151])^(a[108] & b[152])^(a[107] & b[153])^(a[106] & b[154])^(a[105] & b[155])^(a[104] & b[156])^(a[103] & b[157])^(a[102] & b[158])^(a[101] & b[159])^(a[100] & b[160])^(a[99] & b[161])^(a[98] & b[162])^(a[97] & b[163])^(a[96] & b[164])^(a[95] & b[165])^(a[94] & b[166])^(a[93] & b[167])^(a[92] & b[168])^(a[91] & b[169])^(a[90] & b[170])^(a[89] & b[171])^(a[88] & b[172])^(a[87] & b[173])^(a[86] & b[174])^(a[85] & b[175])^(a[84] & b[176])^(a[83] & b[177])^(a[82] & b[178])^(a[81] & b[179])^(a[80] & b[180])^(a[79] & b[181])^(a[78] & b[182])^(a[77] & b[183])^(a[76] & b[184])^(a[75] & b[185])^(a[74] & b[186])^(a[73] & b[187])^(a[72] & b[188])^(a[71] & b[189])^(a[70] & b[190])^(a[69] & b[191])^(a[68] & b[192])^(a[67] & b[193])^(a[66] & b[194])^(a[65] & b[195])^(a[64] & b[196])^(a[63] & b[197])^(a[62] & b[198])^(a[61] & b[199])^(a[60] & b[200])^(a[59] & b[201])^(a[58] & b[202])^(a[57] & b[203])^(a[56] & b[204])^(a[55] & b[205])^(a[54] & b[206])^(a[53] & b[207])^(a[52] & b[208])^(a[51] & b[209])^(a[50] & b[210])^(a[49] & b[211])^(a[48] & b[212])^(a[47] & b[213])^(a[46] & b[214])^(a[45] & b[215])^(a[44] & b[216])^(a[43] & b[217])^(a[42] & b[218])^(a[41] & b[219])^(a[40] & b[220])^(a[39] & b[221])^(a[38] & b[222])^(a[37] & b[223])^(a[36] & b[224])^(a[35] & b[225])^(a[34] & b[226])^(a[33] & b[227])^(a[32] & b[228])^(a[31] & b[229])^(a[30] & b[230])^(a[29] & b[231])^(a[28] & b[232])^(a[27] & b[233])^(a[26] & b[234])^(a[25] & b[235])^(a[24] & b[236])^(a[23] & b[237])^(a[22] & b[238])^(a[21] & b[239])^(a[20] & b[240])^(a[19] & b[241])^(a[18] & b[242])^(a[17] & b[243])^(a[16] & b[244])^(a[15] & b[245])^(a[14] & b[246])^(a[13] & b[247])^(a[12] & b[248])^(a[11] & b[249])^(a[10] & b[250])^(a[9] & b[251])^(a[8] & b[252])^(a[7] & b[253])^(a[6] & b[254])^(a[5] & b[255])^(a[4] & b[256])^(a[3] & b[257])^(a[2] & b[258])^(a[1] & b[259])^(a[0] & b[260]);
assign y[261] = (a[261] & b[0])^(a[260] & b[1])^(a[259] & b[2])^(a[258] & b[3])^(a[257] & b[4])^(a[256] & b[5])^(a[255] & b[6])^(a[254] & b[7])^(a[253] & b[8])^(a[252] & b[9])^(a[251] & b[10])^(a[250] & b[11])^(a[249] & b[12])^(a[248] & b[13])^(a[247] & b[14])^(a[246] & b[15])^(a[245] & b[16])^(a[244] & b[17])^(a[243] & b[18])^(a[242] & b[19])^(a[241] & b[20])^(a[240] & b[21])^(a[239] & b[22])^(a[238] & b[23])^(a[237] & b[24])^(a[236] & b[25])^(a[235] & b[26])^(a[234] & b[27])^(a[233] & b[28])^(a[232] & b[29])^(a[231] & b[30])^(a[230] & b[31])^(a[229] & b[32])^(a[228] & b[33])^(a[227] & b[34])^(a[226] & b[35])^(a[225] & b[36])^(a[224] & b[37])^(a[223] & b[38])^(a[222] & b[39])^(a[221] & b[40])^(a[220] & b[41])^(a[219] & b[42])^(a[218] & b[43])^(a[217] & b[44])^(a[216] & b[45])^(a[215] & b[46])^(a[214] & b[47])^(a[213] & b[48])^(a[212] & b[49])^(a[211] & b[50])^(a[210] & b[51])^(a[209] & b[52])^(a[208] & b[53])^(a[207] & b[54])^(a[206] & b[55])^(a[205] & b[56])^(a[204] & b[57])^(a[203] & b[58])^(a[202] & b[59])^(a[201] & b[60])^(a[200] & b[61])^(a[199] & b[62])^(a[198] & b[63])^(a[197] & b[64])^(a[196] & b[65])^(a[195] & b[66])^(a[194] & b[67])^(a[193] & b[68])^(a[192] & b[69])^(a[191] & b[70])^(a[190] & b[71])^(a[189] & b[72])^(a[188] & b[73])^(a[187] & b[74])^(a[186] & b[75])^(a[185] & b[76])^(a[184] & b[77])^(a[183] & b[78])^(a[182] & b[79])^(a[181] & b[80])^(a[180] & b[81])^(a[179] & b[82])^(a[178] & b[83])^(a[177] & b[84])^(a[176] & b[85])^(a[175] & b[86])^(a[174] & b[87])^(a[173] & b[88])^(a[172] & b[89])^(a[171] & b[90])^(a[170] & b[91])^(a[169] & b[92])^(a[168] & b[93])^(a[167] & b[94])^(a[166] & b[95])^(a[165] & b[96])^(a[164] & b[97])^(a[163] & b[98])^(a[162] & b[99])^(a[161] & b[100])^(a[160] & b[101])^(a[159] & b[102])^(a[158] & b[103])^(a[157] & b[104])^(a[156] & b[105])^(a[155] & b[106])^(a[154] & b[107])^(a[153] & b[108])^(a[152] & b[109])^(a[151] & b[110])^(a[150] & b[111])^(a[149] & b[112])^(a[148] & b[113])^(a[147] & b[114])^(a[146] & b[115])^(a[145] & b[116])^(a[144] & b[117])^(a[143] & b[118])^(a[142] & b[119])^(a[141] & b[120])^(a[140] & b[121])^(a[139] & b[122])^(a[138] & b[123])^(a[137] & b[124])^(a[136] & b[125])^(a[135] & b[126])^(a[134] & b[127])^(a[133] & b[128])^(a[132] & b[129])^(a[131] & b[130])^(a[130] & b[131])^(a[129] & b[132])^(a[128] & b[133])^(a[127] & b[134])^(a[126] & b[135])^(a[125] & b[136])^(a[124] & b[137])^(a[123] & b[138])^(a[122] & b[139])^(a[121] & b[140])^(a[120] & b[141])^(a[119] & b[142])^(a[118] & b[143])^(a[117] & b[144])^(a[116] & b[145])^(a[115] & b[146])^(a[114] & b[147])^(a[113] & b[148])^(a[112] & b[149])^(a[111] & b[150])^(a[110] & b[151])^(a[109] & b[152])^(a[108] & b[153])^(a[107] & b[154])^(a[106] & b[155])^(a[105] & b[156])^(a[104] & b[157])^(a[103] & b[158])^(a[102] & b[159])^(a[101] & b[160])^(a[100] & b[161])^(a[99] & b[162])^(a[98] & b[163])^(a[97] & b[164])^(a[96] & b[165])^(a[95] & b[166])^(a[94] & b[167])^(a[93] & b[168])^(a[92] & b[169])^(a[91] & b[170])^(a[90] & b[171])^(a[89] & b[172])^(a[88] & b[173])^(a[87] & b[174])^(a[86] & b[175])^(a[85] & b[176])^(a[84] & b[177])^(a[83] & b[178])^(a[82] & b[179])^(a[81] & b[180])^(a[80] & b[181])^(a[79] & b[182])^(a[78] & b[183])^(a[77] & b[184])^(a[76] & b[185])^(a[75] & b[186])^(a[74] & b[187])^(a[73] & b[188])^(a[72] & b[189])^(a[71] & b[190])^(a[70] & b[191])^(a[69] & b[192])^(a[68] & b[193])^(a[67] & b[194])^(a[66] & b[195])^(a[65] & b[196])^(a[64] & b[197])^(a[63] & b[198])^(a[62] & b[199])^(a[61] & b[200])^(a[60] & b[201])^(a[59] & b[202])^(a[58] & b[203])^(a[57] & b[204])^(a[56] & b[205])^(a[55] & b[206])^(a[54] & b[207])^(a[53] & b[208])^(a[52] & b[209])^(a[51] & b[210])^(a[50] & b[211])^(a[49] & b[212])^(a[48] & b[213])^(a[47] & b[214])^(a[46] & b[215])^(a[45] & b[216])^(a[44] & b[217])^(a[43] & b[218])^(a[42] & b[219])^(a[41] & b[220])^(a[40] & b[221])^(a[39] & b[222])^(a[38] & b[223])^(a[37] & b[224])^(a[36] & b[225])^(a[35] & b[226])^(a[34] & b[227])^(a[33] & b[228])^(a[32] & b[229])^(a[31] & b[230])^(a[30] & b[231])^(a[29] & b[232])^(a[28] & b[233])^(a[27] & b[234])^(a[26] & b[235])^(a[25] & b[236])^(a[24] & b[237])^(a[23] & b[238])^(a[22] & b[239])^(a[21] & b[240])^(a[20] & b[241])^(a[19] & b[242])^(a[18] & b[243])^(a[17] & b[244])^(a[16] & b[245])^(a[15] & b[246])^(a[14] & b[247])^(a[13] & b[248])^(a[12] & b[249])^(a[11] & b[250])^(a[10] & b[251])^(a[9] & b[252])^(a[8] & b[253])^(a[7] & b[254])^(a[6] & b[255])^(a[5] & b[256])^(a[4] & b[257])^(a[3] & b[258])^(a[2] & b[259])^(a[1] & b[260])^(a[0] & b[261]);
assign y[262] = (a[262] & b[0])^(a[261] & b[1])^(a[260] & b[2])^(a[259] & b[3])^(a[258] & b[4])^(a[257] & b[5])^(a[256] & b[6])^(a[255] & b[7])^(a[254] & b[8])^(a[253] & b[9])^(a[252] & b[10])^(a[251] & b[11])^(a[250] & b[12])^(a[249] & b[13])^(a[248] & b[14])^(a[247] & b[15])^(a[246] & b[16])^(a[245] & b[17])^(a[244] & b[18])^(a[243] & b[19])^(a[242] & b[20])^(a[241] & b[21])^(a[240] & b[22])^(a[239] & b[23])^(a[238] & b[24])^(a[237] & b[25])^(a[236] & b[26])^(a[235] & b[27])^(a[234] & b[28])^(a[233] & b[29])^(a[232] & b[30])^(a[231] & b[31])^(a[230] & b[32])^(a[229] & b[33])^(a[228] & b[34])^(a[227] & b[35])^(a[226] & b[36])^(a[225] & b[37])^(a[224] & b[38])^(a[223] & b[39])^(a[222] & b[40])^(a[221] & b[41])^(a[220] & b[42])^(a[219] & b[43])^(a[218] & b[44])^(a[217] & b[45])^(a[216] & b[46])^(a[215] & b[47])^(a[214] & b[48])^(a[213] & b[49])^(a[212] & b[50])^(a[211] & b[51])^(a[210] & b[52])^(a[209] & b[53])^(a[208] & b[54])^(a[207] & b[55])^(a[206] & b[56])^(a[205] & b[57])^(a[204] & b[58])^(a[203] & b[59])^(a[202] & b[60])^(a[201] & b[61])^(a[200] & b[62])^(a[199] & b[63])^(a[198] & b[64])^(a[197] & b[65])^(a[196] & b[66])^(a[195] & b[67])^(a[194] & b[68])^(a[193] & b[69])^(a[192] & b[70])^(a[191] & b[71])^(a[190] & b[72])^(a[189] & b[73])^(a[188] & b[74])^(a[187] & b[75])^(a[186] & b[76])^(a[185] & b[77])^(a[184] & b[78])^(a[183] & b[79])^(a[182] & b[80])^(a[181] & b[81])^(a[180] & b[82])^(a[179] & b[83])^(a[178] & b[84])^(a[177] & b[85])^(a[176] & b[86])^(a[175] & b[87])^(a[174] & b[88])^(a[173] & b[89])^(a[172] & b[90])^(a[171] & b[91])^(a[170] & b[92])^(a[169] & b[93])^(a[168] & b[94])^(a[167] & b[95])^(a[166] & b[96])^(a[165] & b[97])^(a[164] & b[98])^(a[163] & b[99])^(a[162] & b[100])^(a[161] & b[101])^(a[160] & b[102])^(a[159] & b[103])^(a[158] & b[104])^(a[157] & b[105])^(a[156] & b[106])^(a[155] & b[107])^(a[154] & b[108])^(a[153] & b[109])^(a[152] & b[110])^(a[151] & b[111])^(a[150] & b[112])^(a[149] & b[113])^(a[148] & b[114])^(a[147] & b[115])^(a[146] & b[116])^(a[145] & b[117])^(a[144] & b[118])^(a[143] & b[119])^(a[142] & b[120])^(a[141] & b[121])^(a[140] & b[122])^(a[139] & b[123])^(a[138] & b[124])^(a[137] & b[125])^(a[136] & b[126])^(a[135] & b[127])^(a[134] & b[128])^(a[133] & b[129])^(a[132] & b[130])^(a[131] & b[131])^(a[130] & b[132])^(a[129] & b[133])^(a[128] & b[134])^(a[127] & b[135])^(a[126] & b[136])^(a[125] & b[137])^(a[124] & b[138])^(a[123] & b[139])^(a[122] & b[140])^(a[121] & b[141])^(a[120] & b[142])^(a[119] & b[143])^(a[118] & b[144])^(a[117] & b[145])^(a[116] & b[146])^(a[115] & b[147])^(a[114] & b[148])^(a[113] & b[149])^(a[112] & b[150])^(a[111] & b[151])^(a[110] & b[152])^(a[109] & b[153])^(a[108] & b[154])^(a[107] & b[155])^(a[106] & b[156])^(a[105] & b[157])^(a[104] & b[158])^(a[103] & b[159])^(a[102] & b[160])^(a[101] & b[161])^(a[100] & b[162])^(a[99] & b[163])^(a[98] & b[164])^(a[97] & b[165])^(a[96] & b[166])^(a[95] & b[167])^(a[94] & b[168])^(a[93] & b[169])^(a[92] & b[170])^(a[91] & b[171])^(a[90] & b[172])^(a[89] & b[173])^(a[88] & b[174])^(a[87] & b[175])^(a[86] & b[176])^(a[85] & b[177])^(a[84] & b[178])^(a[83] & b[179])^(a[82] & b[180])^(a[81] & b[181])^(a[80] & b[182])^(a[79] & b[183])^(a[78] & b[184])^(a[77] & b[185])^(a[76] & b[186])^(a[75] & b[187])^(a[74] & b[188])^(a[73] & b[189])^(a[72] & b[190])^(a[71] & b[191])^(a[70] & b[192])^(a[69] & b[193])^(a[68] & b[194])^(a[67] & b[195])^(a[66] & b[196])^(a[65] & b[197])^(a[64] & b[198])^(a[63] & b[199])^(a[62] & b[200])^(a[61] & b[201])^(a[60] & b[202])^(a[59] & b[203])^(a[58] & b[204])^(a[57] & b[205])^(a[56] & b[206])^(a[55] & b[207])^(a[54] & b[208])^(a[53] & b[209])^(a[52] & b[210])^(a[51] & b[211])^(a[50] & b[212])^(a[49] & b[213])^(a[48] & b[214])^(a[47] & b[215])^(a[46] & b[216])^(a[45] & b[217])^(a[44] & b[218])^(a[43] & b[219])^(a[42] & b[220])^(a[41] & b[221])^(a[40] & b[222])^(a[39] & b[223])^(a[38] & b[224])^(a[37] & b[225])^(a[36] & b[226])^(a[35] & b[227])^(a[34] & b[228])^(a[33] & b[229])^(a[32] & b[230])^(a[31] & b[231])^(a[30] & b[232])^(a[29] & b[233])^(a[28] & b[234])^(a[27] & b[235])^(a[26] & b[236])^(a[25] & b[237])^(a[24] & b[238])^(a[23] & b[239])^(a[22] & b[240])^(a[21] & b[241])^(a[20] & b[242])^(a[19] & b[243])^(a[18] & b[244])^(a[17] & b[245])^(a[16] & b[246])^(a[15] & b[247])^(a[14] & b[248])^(a[13] & b[249])^(a[12] & b[250])^(a[11] & b[251])^(a[10] & b[252])^(a[9] & b[253])^(a[8] & b[254])^(a[7] & b[255])^(a[6] & b[256])^(a[5] & b[257])^(a[4] & b[258])^(a[3] & b[259])^(a[2] & b[260])^(a[1] & b[261])^(a[0] & b[262]);
assign y[263] = (a[263] & b[0])^(a[262] & b[1])^(a[261] & b[2])^(a[260] & b[3])^(a[259] & b[4])^(a[258] & b[5])^(a[257] & b[6])^(a[256] & b[7])^(a[255] & b[8])^(a[254] & b[9])^(a[253] & b[10])^(a[252] & b[11])^(a[251] & b[12])^(a[250] & b[13])^(a[249] & b[14])^(a[248] & b[15])^(a[247] & b[16])^(a[246] & b[17])^(a[245] & b[18])^(a[244] & b[19])^(a[243] & b[20])^(a[242] & b[21])^(a[241] & b[22])^(a[240] & b[23])^(a[239] & b[24])^(a[238] & b[25])^(a[237] & b[26])^(a[236] & b[27])^(a[235] & b[28])^(a[234] & b[29])^(a[233] & b[30])^(a[232] & b[31])^(a[231] & b[32])^(a[230] & b[33])^(a[229] & b[34])^(a[228] & b[35])^(a[227] & b[36])^(a[226] & b[37])^(a[225] & b[38])^(a[224] & b[39])^(a[223] & b[40])^(a[222] & b[41])^(a[221] & b[42])^(a[220] & b[43])^(a[219] & b[44])^(a[218] & b[45])^(a[217] & b[46])^(a[216] & b[47])^(a[215] & b[48])^(a[214] & b[49])^(a[213] & b[50])^(a[212] & b[51])^(a[211] & b[52])^(a[210] & b[53])^(a[209] & b[54])^(a[208] & b[55])^(a[207] & b[56])^(a[206] & b[57])^(a[205] & b[58])^(a[204] & b[59])^(a[203] & b[60])^(a[202] & b[61])^(a[201] & b[62])^(a[200] & b[63])^(a[199] & b[64])^(a[198] & b[65])^(a[197] & b[66])^(a[196] & b[67])^(a[195] & b[68])^(a[194] & b[69])^(a[193] & b[70])^(a[192] & b[71])^(a[191] & b[72])^(a[190] & b[73])^(a[189] & b[74])^(a[188] & b[75])^(a[187] & b[76])^(a[186] & b[77])^(a[185] & b[78])^(a[184] & b[79])^(a[183] & b[80])^(a[182] & b[81])^(a[181] & b[82])^(a[180] & b[83])^(a[179] & b[84])^(a[178] & b[85])^(a[177] & b[86])^(a[176] & b[87])^(a[175] & b[88])^(a[174] & b[89])^(a[173] & b[90])^(a[172] & b[91])^(a[171] & b[92])^(a[170] & b[93])^(a[169] & b[94])^(a[168] & b[95])^(a[167] & b[96])^(a[166] & b[97])^(a[165] & b[98])^(a[164] & b[99])^(a[163] & b[100])^(a[162] & b[101])^(a[161] & b[102])^(a[160] & b[103])^(a[159] & b[104])^(a[158] & b[105])^(a[157] & b[106])^(a[156] & b[107])^(a[155] & b[108])^(a[154] & b[109])^(a[153] & b[110])^(a[152] & b[111])^(a[151] & b[112])^(a[150] & b[113])^(a[149] & b[114])^(a[148] & b[115])^(a[147] & b[116])^(a[146] & b[117])^(a[145] & b[118])^(a[144] & b[119])^(a[143] & b[120])^(a[142] & b[121])^(a[141] & b[122])^(a[140] & b[123])^(a[139] & b[124])^(a[138] & b[125])^(a[137] & b[126])^(a[136] & b[127])^(a[135] & b[128])^(a[134] & b[129])^(a[133] & b[130])^(a[132] & b[131])^(a[131] & b[132])^(a[130] & b[133])^(a[129] & b[134])^(a[128] & b[135])^(a[127] & b[136])^(a[126] & b[137])^(a[125] & b[138])^(a[124] & b[139])^(a[123] & b[140])^(a[122] & b[141])^(a[121] & b[142])^(a[120] & b[143])^(a[119] & b[144])^(a[118] & b[145])^(a[117] & b[146])^(a[116] & b[147])^(a[115] & b[148])^(a[114] & b[149])^(a[113] & b[150])^(a[112] & b[151])^(a[111] & b[152])^(a[110] & b[153])^(a[109] & b[154])^(a[108] & b[155])^(a[107] & b[156])^(a[106] & b[157])^(a[105] & b[158])^(a[104] & b[159])^(a[103] & b[160])^(a[102] & b[161])^(a[101] & b[162])^(a[100] & b[163])^(a[99] & b[164])^(a[98] & b[165])^(a[97] & b[166])^(a[96] & b[167])^(a[95] & b[168])^(a[94] & b[169])^(a[93] & b[170])^(a[92] & b[171])^(a[91] & b[172])^(a[90] & b[173])^(a[89] & b[174])^(a[88] & b[175])^(a[87] & b[176])^(a[86] & b[177])^(a[85] & b[178])^(a[84] & b[179])^(a[83] & b[180])^(a[82] & b[181])^(a[81] & b[182])^(a[80] & b[183])^(a[79] & b[184])^(a[78] & b[185])^(a[77] & b[186])^(a[76] & b[187])^(a[75] & b[188])^(a[74] & b[189])^(a[73] & b[190])^(a[72] & b[191])^(a[71] & b[192])^(a[70] & b[193])^(a[69] & b[194])^(a[68] & b[195])^(a[67] & b[196])^(a[66] & b[197])^(a[65] & b[198])^(a[64] & b[199])^(a[63] & b[200])^(a[62] & b[201])^(a[61] & b[202])^(a[60] & b[203])^(a[59] & b[204])^(a[58] & b[205])^(a[57] & b[206])^(a[56] & b[207])^(a[55] & b[208])^(a[54] & b[209])^(a[53] & b[210])^(a[52] & b[211])^(a[51] & b[212])^(a[50] & b[213])^(a[49] & b[214])^(a[48] & b[215])^(a[47] & b[216])^(a[46] & b[217])^(a[45] & b[218])^(a[44] & b[219])^(a[43] & b[220])^(a[42] & b[221])^(a[41] & b[222])^(a[40] & b[223])^(a[39] & b[224])^(a[38] & b[225])^(a[37] & b[226])^(a[36] & b[227])^(a[35] & b[228])^(a[34] & b[229])^(a[33] & b[230])^(a[32] & b[231])^(a[31] & b[232])^(a[30] & b[233])^(a[29] & b[234])^(a[28] & b[235])^(a[27] & b[236])^(a[26] & b[237])^(a[25] & b[238])^(a[24] & b[239])^(a[23] & b[240])^(a[22] & b[241])^(a[21] & b[242])^(a[20] & b[243])^(a[19] & b[244])^(a[18] & b[245])^(a[17] & b[246])^(a[16] & b[247])^(a[15] & b[248])^(a[14] & b[249])^(a[13] & b[250])^(a[12] & b[251])^(a[11] & b[252])^(a[10] & b[253])^(a[9] & b[254])^(a[8] & b[255])^(a[7] & b[256])^(a[6] & b[257])^(a[5] & b[258])^(a[4] & b[259])^(a[3] & b[260])^(a[2] & b[261])^(a[1] & b[262])^(a[0] & b[263]);
assign y[264] = (a[264] & b[0])^(a[263] & b[1])^(a[262] & b[2])^(a[261] & b[3])^(a[260] & b[4])^(a[259] & b[5])^(a[258] & b[6])^(a[257] & b[7])^(a[256] & b[8])^(a[255] & b[9])^(a[254] & b[10])^(a[253] & b[11])^(a[252] & b[12])^(a[251] & b[13])^(a[250] & b[14])^(a[249] & b[15])^(a[248] & b[16])^(a[247] & b[17])^(a[246] & b[18])^(a[245] & b[19])^(a[244] & b[20])^(a[243] & b[21])^(a[242] & b[22])^(a[241] & b[23])^(a[240] & b[24])^(a[239] & b[25])^(a[238] & b[26])^(a[237] & b[27])^(a[236] & b[28])^(a[235] & b[29])^(a[234] & b[30])^(a[233] & b[31])^(a[232] & b[32])^(a[231] & b[33])^(a[230] & b[34])^(a[229] & b[35])^(a[228] & b[36])^(a[227] & b[37])^(a[226] & b[38])^(a[225] & b[39])^(a[224] & b[40])^(a[223] & b[41])^(a[222] & b[42])^(a[221] & b[43])^(a[220] & b[44])^(a[219] & b[45])^(a[218] & b[46])^(a[217] & b[47])^(a[216] & b[48])^(a[215] & b[49])^(a[214] & b[50])^(a[213] & b[51])^(a[212] & b[52])^(a[211] & b[53])^(a[210] & b[54])^(a[209] & b[55])^(a[208] & b[56])^(a[207] & b[57])^(a[206] & b[58])^(a[205] & b[59])^(a[204] & b[60])^(a[203] & b[61])^(a[202] & b[62])^(a[201] & b[63])^(a[200] & b[64])^(a[199] & b[65])^(a[198] & b[66])^(a[197] & b[67])^(a[196] & b[68])^(a[195] & b[69])^(a[194] & b[70])^(a[193] & b[71])^(a[192] & b[72])^(a[191] & b[73])^(a[190] & b[74])^(a[189] & b[75])^(a[188] & b[76])^(a[187] & b[77])^(a[186] & b[78])^(a[185] & b[79])^(a[184] & b[80])^(a[183] & b[81])^(a[182] & b[82])^(a[181] & b[83])^(a[180] & b[84])^(a[179] & b[85])^(a[178] & b[86])^(a[177] & b[87])^(a[176] & b[88])^(a[175] & b[89])^(a[174] & b[90])^(a[173] & b[91])^(a[172] & b[92])^(a[171] & b[93])^(a[170] & b[94])^(a[169] & b[95])^(a[168] & b[96])^(a[167] & b[97])^(a[166] & b[98])^(a[165] & b[99])^(a[164] & b[100])^(a[163] & b[101])^(a[162] & b[102])^(a[161] & b[103])^(a[160] & b[104])^(a[159] & b[105])^(a[158] & b[106])^(a[157] & b[107])^(a[156] & b[108])^(a[155] & b[109])^(a[154] & b[110])^(a[153] & b[111])^(a[152] & b[112])^(a[151] & b[113])^(a[150] & b[114])^(a[149] & b[115])^(a[148] & b[116])^(a[147] & b[117])^(a[146] & b[118])^(a[145] & b[119])^(a[144] & b[120])^(a[143] & b[121])^(a[142] & b[122])^(a[141] & b[123])^(a[140] & b[124])^(a[139] & b[125])^(a[138] & b[126])^(a[137] & b[127])^(a[136] & b[128])^(a[135] & b[129])^(a[134] & b[130])^(a[133] & b[131])^(a[132] & b[132])^(a[131] & b[133])^(a[130] & b[134])^(a[129] & b[135])^(a[128] & b[136])^(a[127] & b[137])^(a[126] & b[138])^(a[125] & b[139])^(a[124] & b[140])^(a[123] & b[141])^(a[122] & b[142])^(a[121] & b[143])^(a[120] & b[144])^(a[119] & b[145])^(a[118] & b[146])^(a[117] & b[147])^(a[116] & b[148])^(a[115] & b[149])^(a[114] & b[150])^(a[113] & b[151])^(a[112] & b[152])^(a[111] & b[153])^(a[110] & b[154])^(a[109] & b[155])^(a[108] & b[156])^(a[107] & b[157])^(a[106] & b[158])^(a[105] & b[159])^(a[104] & b[160])^(a[103] & b[161])^(a[102] & b[162])^(a[101] & b[163])^(a[100] & b[164])^(a[99] & b[165])^(a[98] & b[166])^(a[97] & b[167])^(a[96] & b[168])^(a[95] & b[169])^(a[94] & b[170])^(a[93] & b[171])^(a[92] & b[172])^(a[91] & b[173])^(a[90] & b[174])^(a[89] & b[175])^(a[88] & b[176])^(a[87] & b[177])^(a[86] & b[178])^(a[85] & b[179])^(a[84] & b[180])^(a[83] & b[181])^(a[82] & b[182])^(a[81] & b[183])^(a[80] & b[184])^(a[79] & b[185])^(a[78] & b[186])^(a[77] & b[187])^(a[76] & b[188])^(a[75] & b[189])^(a[74] & b[190])^(a[73] & b[191])^(a[72] & b[192])^(a[71] & b[193])^(a[70] & b[194])^(a[69] & b[195])^(a[68] & b[196])^(a[67] & b[197])^(a[66] & b[198])^(a[65] & b[199])^(a[64] & b[200])^(a[63] & b[201])^(a[62] & b[202])^(a[61] & b[203])^(a[60] & b[204])^(a[59] & b[205])^(a[58] & b[206])^(a[57] & b[207])^(a[56] & b[208])^(a[55] & b[209])^(a[54] & b[210])^(a[53] & b[211])^(a[52] & b[212])^(a[51] & b[213])^(a[50] & b[214])^(a[49] & b[215])^(a[48] & b[216])^(a[47] & b[217])^(a[46] & b[218])^(a[45] & b[219])^(a[44] & b[220])^(a[43] & b[221])^(a[42] & b[222])^(a[41] & b[223])^(a[40] & b[224])^(a[39] & b[225])^(a[38] & b[226])^(a[37] & b[227])^(a[36] & b[228])^(a[35] & b[229])^(a[34] & b[230])^(a[33] & b[231])^(a[32] & b[232])^(a[31] & b[233])^(a[30] & b[234])^(a[29] & b[235])^(a[28] & b[236])^(a[27] & b[237])^(a[26] & b[238])^(a[25] & b[239])^(a[24] & b[240])^(a[23] & b[241])^(a[22] & b[242])^(a[21] & b[243])^(a[20] & b[244])^(a[19] & b[245])^(a[18] & b[246])^(a[17] & b[247])^(a[16] & b[248])^(a[15] & b[249])^(a[14] & b[250])^(a[13] & b[251])^(a[12] & b[252])^(a[11] & b[253])^(a[10] & b[254])^(a[9] & b[255])^(a[8] & b[256])^(a[7] & b[257])^(a[6] & b[258])^(a[5] & b[259])^(a[4] & b[260])^(a[3] & b[261])^(a[2] & b[262])^(a[1] & b[263])^(a[0] & b[264]);
assign y[265] = (a[265] & b[0])^(a[264] & b[1])^(a[263] & b[2])^(a[262] & b[3])^(a[261] & b[4])^(a[260] & b[5])^(a[259] & b[6])^(a[258] & b[7])^(a[257] & b[8])^(a[256] & b[9])^(a[255] & b[10])^(a[254] & b[11])^(a[253] & b[12])^(a[252] & b[13])^(a[251] & b[14])^(a[250] & b[15])^(a[249] & b[16])^(a[248] & b[17])^(a[247] & b[18])^(a[246] & b[19])^(a[245] & b[20])^(a[244] & b[21])^(a[243] & b[22])^(a[242] & b[23])^(a[241] & b[24])^(a[240] & b[25])^(a[239] & b[26])^(a[238] & b[27])^(a[237] & b[28])^(a[236] & b[29])^(a[235] & b[30])^(a[234] & b[31])^(a[233] & b[32])^(a[232] & b[33])^(a[231] & b[34])^(a[230] & b[35])^(a[229] & b[36])^(a[228] & b[37])^(a[227] & b[38])^(a[226] & b[39])^(a[225] & b[40])^(a[224] & b[41])^(a[223] & b[42])^(a[222] & b[43])^(a[221] & b[44])^(a[220] & b[45])^(a[219] & b[46])^(a[218] & b[47])^(a[217] & b[48])^(a[216] & b[49])^(a[215] & b[50])^(a[214] & b[51])^(a[213] & b[52])^(a[212] & b[53])^(a[211] & b[54])^(a[210] & b[55])^(a[209] & b[56])^(a[208] & b[57])^(a[207] & b[58])^(a[206] & b[59])^(a[205] & b[60])^(a[204] & b[61])^(a[203] & b[62])^(a[202] & b[63])^(a[201] & b[64])^(a[200] & b[65])^(a[199] & b[66])^(a[198] & b[67])^(a[197] & b[68])^(a[196] & b[69])^(a[195] & b[70])^(a[194] & b[71])^(a[193] & b[72])^(a[192] & b[73])^(a[191] & b[74])^(a[190] & b[75])^(a[189] & b[76])^(a[188] & b[77])^(a[187] & b[78])^(a[186] & b[79])^(a[185] & b[80])^(a[184] & b[81])^(a[183] & b[82])^(a[182] & b[83])^(a[181] & b[84])^(a[180] & b[85])^(a[179] & b[86])^(a[178] & b[87])^(a[177] & b[88])^(a[176] & b[89])^(a[175] & b[90])^(a[174] & b[91])^(a[173] & b[92])^(a[172] & b[93])^(a[171] & b[94])^(a[170] & b[95])^(a[169] & b[96])^(a[168] & b[97])^(a[167] & b[98])^(a[166] & b[99])^(a[165] & b[100])^(a[164] & b[101])^(a[163] & b[102])^(a[162] & b[103])^(a[161] & b[104])^(a[160] & b[105])^(a[159] & b[106])^(a[158] & b[107])^(a[157] & b[108])^(a[156] & b[109])^(a[155] & b[110])^(a[154] & b[111])^(a[153] & b[112])^(a[152] & b[113])^(a[151] & b[114])^(a[150] & b[115])^(a[149] & b[116])^(a[148] & b[117])^(a[147] & b[118])^(a[146] & b[119])^(a[145] & b[120])^(a[144] & b[121])^(a[143] & b[122])^(a[142] & b[123])^(a[141] & b[124])^(a[140] & b[125])^(a[139] & b[126])^(a[138] & b[127])^(a[137] & b[128])^(a[136] & b[129])^(a[135] & b[130])^(a[134] & b[131])^(a[133] & b[132])^(a[132] & b[133])^(a[131] & b[134])^(a[130] & b[135])^(a[129] & b[136])^(a[128] & b[137])^(a[127] & b[138])^(a[126] & b[139])^(a[125] & b[140])^(a[124] & b[141])^(a[123] & b[142])^(a[122] & b[143])^(a[121] & b[144])^(a[120] & b[145])^(a[119] & b[146])^(a[118] & b[147])^(a[117] & b[148])^(a[116] & b[149])^(a[115] & b[150])^(a[114] & b[151])^(a[113] & b[152])^(a[112] & b[153])^(a[111] & b[154])^(a[110] & b[155])^(a[109] & b[156])^(a[108] & b[157])^(a[107] & b[158])^(a[106] & b[159])^(a[105] & b[160])^(a[104] & b[161])^(a[103] & b[162])^(a[102] & b[163])^(a[101] & b[164])^(a[100] & b[165])^(a[99] & b[166])^(a[98] & b[167])^(a[97] & b[168])^(a[96] & b[169])^(a[95] & b[170])^(a[94] & b[171])^(a[93] & b[172])^(a[92] & b[173])^(a[91] & b[174])^(a[90] & b[175])^(a[89] & b[176])^(a[88] & b[177])^(a[87] & b[178])^(a[86] & b[179])^(a[85] & b[180])^(a[84] & b[181])^(a[83] & b[182])^(a[82] & b[183])^(a[81] & b[184])^(a[80] & b[185])^(a[79] & b[186])^(a[78] & b[187])^(a[77] & b[188])^(a[76] & b[189])^(a[75] & b[190])^(a[74] & b[191])^(a[73] & b[192])^(a[72] & b[193])^(a[71] & b[194])^(a[70] & b[195])^(a[69] & b[196])^(a[68] & b[197])^(a[67] & b[198])^(a[66] & b[199])^(a[65] & b[200])^(a[64] & b[201])^(a[63] & b[202])^(a[62] & b[203])^(a[61] & b[204])^(a[60] & b[205])^(a[59] & b[206])^(a[58] & b[207])^(a[57] & b[208])^(a[56] & b[209])^(a[55] & b[210])^(a[54] & b[211])^(a[53] & b[212])^(a[52] & b[213])^(a[51] & b[214])^(a[50] & b[215])^(a[49] & b[216])^(a[48] & b[217])^(a[47] & b[218])^(a[46] & b[219])^(a[45] & b[220])^(a[44] & b[221])^(a[43] & b[222])^(a[42] & b[223])^(a[41] & b[224])^(a[40] & b[225])^(a[39] & b[226])^(a[38] & b[227])^(a[37] & b[228])^(a[36] & b[229])^(a[35] & b[230])^(a[34] & b[231])^(a[33] & b[232])^(a[32] & b[233])^(a[31] & b[234])^(a[30] & b[235])^(a[29] & b[236])^(a[28] & b[237])^(a[27] & b[238])^(a[26] & b[239])^(a[25] & b[240])^(a[24] & b[241])^(a[23] & b[242])^(a[22] & b[243])^(a[21] & b[244])^(a[20] & b[245])^(a[19] & b[246])^(a[18] & b[247])^(a[17] & b[248])^(a[16] & b[249])^(a[15] & b[250])^(a[14] & b[251])^(a[13] & b[252])^(a[12] & b[253])^(a[11] & b[254])^(a[10] & b[255])^(a[9] & b[256])^(a[8] & b[257])^(a[7] & b[258])^(a[6] & b[259])^(a[5] & b[260])^(a[4] & b[261])^(a[3] & b[262])^(a[2] & b[263])^(a[1] & b[264])^(a[0] & b[265]);
assign y[266] = (a[266] & b[0])^(a[265] & b[1])^(a[264] & b[2])^(a[263] & b[3])^(a[262] & b[4])^(a[261] & b[5])^(a[260] & b[6])^(a[259] & b[7])^(a[258] & b[8])^(a[257] & b[9])^(a[256] & b[10])^(a[255] & b[11])^(a[254] & b[12])^(a[253] & b[13])^(a[252] & b[14])^(a[251] & b[15])^(a[250] & b[16])^(a[249] & b[17])^(a[248] & b[18])^(a[247] & b[19])^(a[246] & b[20])^(a[245] & b[21])^(a[244] & b[22])^(a[243] & b[23])^(a[242] & b[24])^(a[241] & b[25])^(a[240] & b[26])^(a[239] & b[27])^(a[238] & b[28])^(a[237] & b[29])^(a[236] & b[30])^(a[235] & b[31])^(a[234] & b[32])^(a[233] & b[33])^(a[232] & b[34])^(a[231] & b[35])^(a[230] & b[36])^(a[229] & b[37])^(a[228] & b[38])^(a[227] & b[39])^(a[226] & b[40])^(a[225] & b[41])^(a[224] & b[42])^(a[223] & b[43])^(a[222] & b[44])^(a[221] & b[45])^(a[220] & b[46])^(a[219] & b[47])^(a[218] & b[48])^(a[217] & b[49])^(a[216] & b[50])^(a[215] & b[51])^(a[214] & b[52])^(a[213] & b[53])^(a[212] & b[54])^(a[211] & b[55])^(a[210] & b[56])^(a[209] & b[57])^(a[208] & b[58])^(a[207] & b[59])^(a[206] & b[60])^(a[205] & b[61])^(a[204] & b[62])^(a[203] & b[63])^(a[202] & b[64])^(a[201] & b[65])^(a[200] & b[66])^(a[199] & b[67])^(a[198] & b[68])^(a[197] & b[69])^(a[196] & b[70])^(a[195] & b[71])^(a[194] & b[72])^(a[193] & b[73])^(a[192] & b[74])^(a[191] & b[75])^(a[190] & b[76])^(a[189] & b[77])^(a[188] & b[78])^(a[187] & b[79])^(a[186] & b[80])^(a[185] & b[81])^(a[184] & b[82])^(a[183] & b[83])^(a[182] & b[84])^(a[181] & b[85])^(a[180] & b[86])^(a[179] & b[87])^(a[178] & b[88])^(a[177] & b[89])^(a[176] & b[90])^(a[175] & b[91])^(a[174] & b[92])^(a[173] & b[93])^(a[172] & b[94])^(a[171] & b[95])^(a[170] & b[96])^(a[169] & b[97])^(a[168] & b[98])^(a[167] & b[99])^(a[166] & b[100])^(a[165] & b[101])^(a[164] & b[102])^(a[163] & b[103])^(a[162] & b[104])^(a[161] & b[105])^(a[160] & b[106])^(a[159] & b[107])^(a[158] & b[108])^(a[157] & b[109])^(a[156] & b[110])^(a[155] & b[111])^(a[154] & b[112])^(a[153] & b[113])^(a[152] & b[114])^(a[151] & b[115])^(a[150] & b[116])^(a[149] & b[117])^(a[148] & b[118])^(a[147] & b[119])^(a[146] & b[120])^(a[145] & b[121])^(a[144] & b[122])^(a[143] & b[123])^(a[142] & b[124])^(a[141] & b[125])^(a[140] & b[126])^(a[139] & b[127])^(a[138] & b[128])^(a[137] & b[129])^(a[136] & b[130])^(a[135] & b[131])^(a[134] & b[132])^(a[133] & b[133])^(a[132] & b[134])^(a[131] & b[135])^(a[130] & b[136])^(a[129] & b[137])^(a[128] & b[138])^(a[127] & b[139])^(a[126] & b[140])^(a[125] & b[141])^(a[124] & b[142])^(a[123] & b[143])^(a[122] & b[144])^(a[121] & b[145])^(a[120] & b[146])^(a[119] & b[147])^(a[118] & b[148])^(a[117] & b[149])^(a[116] & b[150])^(a[115] & b[151])^(a[114] & b[152])^(a[113] & b[153])^(a[112] & b[154])^(a[111] & b[155])^(a[110] & b[156])^(a[109] & b[157])^(a[108] & b[158])^(a[107] & b[159])^(a[106] & b[160])^(a[105] & b[161])^(a[104] & b[162])^(a[103] & b[163])^(a[102] & b[164])^(a[101] & b[165])^(a[100] & b[166])^(a[99] & b[167])^(a[98] & b[168])^(a[97] & b[169])^(a[96] & b[170])^(a[95] & b[171])^(a[94] & b[172])^(a[93] & b[173])^(a[92] & b[174])^(a[91] & b[175])^(a[90] & b[176])^(a[89] & b[177])^(a[88] & b[178])^(a[87] & b[179])^(a[86] & b[180])^(a[85] & b[181])^(a[84] & b[182])^(a[83] & b[183])^(a[82] & b[184])^(a[81] & b[185])^(a[80] & b[186])^(a[79] & b[187])^(a[78] & b[188])^(a[77] & b[189])^(a[76] & b[190])^(a[75] & b[191])^(a[74] & b[192])^(a[73] & b[193])^(a[72] & b[194])^(a[71] & b[195])^(a[70] & b[196])^(a[69] & b[197])^(a[68] & b[198])^(a[67] & b[199])^(a[66] & b[200])^(a[65] & b[201])^(a[64] & b[202])^(a[63] & b[203])^(a[62] & b[204])^(a[61] & b[205])^(a[60] & b[206])^(a[59] & b[207])^(a[58] & b[208])^(a[57] & b[209])^(a[56] & b[210])^(a[55] & b[211])^(a[54] & b[212])^(a[53] & b[213])^(a[52] & b[214])^(a[51] & b[215])^(a[50] & b[216])^(a[49] & b[217])^(a[48] & b[218])^(a[47] & b[219])^(a[46] & b[220])^(a[45] & b[221])^(a[44] & b[222])^(a[43] & b[223])^(a[42] & b[224])^(a[41] & b[225])^(a[40] & b[226])^(a[39] & b[227])^(a[38] & b[228])^(a[37] & b[229])^(a[36] & b[230])^(a[35] & b[231])^(a[34] & b[232])^(a[33] & b[233])^(a[32] & b[234])^(a[31] & b[235])^(a[30] & b[236])^(a[29] & b[237])^(a[28] & b[238])^(a[27] & b[239])^(a[26] & b[240])^(a[25] & b[241])^(a[24] & b[242])^(a[23] & b[243])^(a[22] & b[244])^(a[21] & b[245])^(a[20] & b[246])^(a[19] & b[247])^(a[18] & b[248])^(a[17] & b[249])^(a[16] & b[250])^(a[15] & b[251])^(a[14] & b[252])^(a[13] & b[253])^(a[12] & b[254])^(a[11] & b[255])^(a[10] & b[256])^(a[9] & b[257])^(a[8] & b[258])^(a[7] & b[259])^(a[6] & b[260])^(a[5] & b[261])^(a[4] & b[262])^(a[3] & b[263])^(a[2] & b[264])^(a[1] & b[265])^(a[0] & b[266]);
assign y[267] = (a[267] & b[0])^(a[266] & b[1])^(a[265] & b[2])^(a[264] & b[3])^(a[263] & b[4])^(a[262] & b[5])^(a[261] & b[6])^(a[260] & b[7])^(a[259] & b[8])^(a[258] & b[9])^(a[257] & b[10])^(a[256] & b[11])^(a[255] & b[12])^(a[254] & b[13])^(a[253] & b[14])^(a[252] & b[15])^(a[251] & b[16])^(a[250] & b[17])^(a[249] & b[18])^(a[248] & b[19])^(a[247] & b[20])^(a[246] & b[21])^(a[245] & b[22])^(a[244] & b[23])^(a[243] & b[24])^(a[242] & b[25])^(a[241] & b[26])^(a[240] & b[27])^(a[239] & b[28])^(a[238] & b[29])^(a[237] & b[30])^(a[236] & b[31])^(a[235] & b[32])^(a[234] & b[33])^(a[233] & b[34])^(a[232] & b[35])^(a[231] & b[36])^(a[230] & b[37])^(a[229] & b[38])^(a[228] & b[39])^(a[227] & b[40])^(a[226] & b[41])^(a[225] & b[42])^(a[224] & b[43])^(a[223] & b[44])^(a[222] & b[45])^(a[221] & b[46])^(a[220] & b[47])^(a[219] & b[48])^(a[218] & b[49])^(a[217] & b[50])^(a[216] & b[51])^(a[215] & b[52])^(a[214] & b[53])^(a[213] & b[54])^(a[212] & b[55])^(a[211] & b[56])^(a[210] & b[57])^(a[209] & b[58])^(a[208] & b[59])^(a[207] & b[60])^(a[206] & b[61])^(a[205] & b[62])^(a[204] & b[63])^(a[203] & b[64])^(a[202] & b[65])^(a[201] & b[66])^(a[200] & b[67])^(a[199] & b[68])^(a[198] & b[69])^(a[197] & b[70])^(a[196] & b[71])^(a[195] & b[72])^(a[194] & b[73])^(a[193] & b[74])^(a[192] & b[75])^(a[191] & b[76])^(a[190] & b[77])^(a[189] & b[78])^(a[188] & b[79])^(a[187] & b[80])^(a[186] & b[81])^(a[185] & b[82])^(a[184] & b[83])^(a[183] & b[84])^(a[182] & b[85])^(a[181] & b[86])^(a[180] & b[87])^(a[179] & b[88])^(a[178] & b[89])^(a[177] & b[90])^(a[176] & b[91])^(a[175] & b[92])^(a[174] & b[93])^(a[173] & b[94])^(a[172] & b[95])^(a[171] & b[96])^(a[170] & b[97])^(a[169] & b[98])^(a[168] & b[99])^(a[167] & b[100])^(a[166] & b[101])^(a[165] & b[102])^(a[164] & b[103])^(a[163] & b[104])^(a[162] & b[105])^(a[161] & b[106])^(a[160] & b[107])^(a[159] & b[108])^(a[158] & b[109])^(a[157] & b[110])^(a[156] & b[111])^(a[155] & b[112])^(a[154] & b[113])^(a[153] & b[114])^(a[152] & b[115])^(a[151] & b[116])^(a[150] & b[117])^(a[149] & b[118])^(a[148] & b[119])^(a[147] & b[120])^(a[146] & b[121])^(a[145] & b[122])^(a[144] & b[123])^(a[143] & b[124])^(a[142] & b[125])^(a[141] & b[126])^(a[140] & b[127])^(a[139] & b[128])^(a[138] & b[129])^(a[137] & b[130])^(a[136] & b[131])^(a[135] & b[132])^(a[134] & b[133])^(a[133] & b[134])^(a[132] & b[135])^(a[131] & b[136])^(a[130] & b[137])^(a[129] & b[138])^(a[128] & b[139])^(a[127] & b[140])^(a[126] & b[141])^(a[125] & b[142])^(a[124] & b[143])^(a[123] & b[144])^(a[122] & b[145])^(a[121] & b[146])^(a[120] & b[147])^(a[119] & b[148])^(a[118] & b[149])^(a[117] & b[150])^(a[116] & b[151])^(a[115] & b[152])^(a[114] & b[153])^(a[113] & b[154])^(a[112] & b[155])^(a[111] & b[156])^(a[110] & b[157])^(a[109] & b[158])^(a[108] & b[159])^(a[107] & b[160])^(a[106] & b[161])^(a[105] & b[162])^(a[104] & b[163])^(a[103] & b[164])^(a[102] & b[165])^(a[101] & b[166])^(a[100] & b[167])^(a[99] & b[168])^(a[98] & b[169])^(a[97] & b[170])^(a[96] & b[171])^(a[95] & b[172])^(a[94] & b[173])^(a[93] & b[174])^(a[92] & b[175])^(a[91] & b[176])^(a[90] & b[177])^(a[89] & b[178])^(a[88] & b[179])^(a[87] & b[180])^(a[86] & b[181])^(a[85] & b[182])^(a[84] & b[183])^(a[83] & b[184])^(a[82] & b[185])^(a[81] & b[186])^(a[80] & b[187])^(a[79] & b[188])^(a[78] & b[189])^(a[77] & b[190])^(a[76] & b[191])^(a[75] & b[192])^(a[74] & b[193])^(a[73] & b[194])^(a[72] & b[195])^(a[71] & b[196])^(a[70] & b[197])^(a[69] & b[198])^(a[68] & b[199])^(a[67] & b[200])^(a[66] & b[201])^(a[65] & b[202])^(a[64] & b[203])^(a[63] & b[204])^(a[62] & b[205])^(a[61] & b[206])^(a[60] & b[207])^(a[59] & b[208])^(a[58] & b[209])^(a[57] & b[210])^(a[56] & b[211])^(a[55] & b[212])^(a[54] & b[213])^(a[53] & b[214])^(a[52] & b[215])^(a[51] & b[216])^(a[50] & b[217])^(a[49] & b[218])^(a[48] & b[219])^(a[47] & b[220])^(a[46] & b[221])^(a[45] & b[222])^(a[44] & b[223])^(a[43] & b[224])^(a[42] & b[225])^(a[41] & b[226])^(a[40] & b[227])^(a[39] & b[228])^(a[38] & b[229])^(a[37] & b[230])^(a[36] & b[231])^(a[35] & b[232])^(a[34] & b[233])^(a[33] & b[234])^(a[32] & b[235])^(a[31] & b[236])^(a[30] & b[237])^(a[29] & b[238])^(a[28] & b[239])^(a[27] & b[240])^(a[26] & b[241])^(a[25] & b[242])^(a[24] & b[243])^(a[23] & b[244])^(a[22] & b[245])^(a[21] & b[246])^(a[20] & b[247])^(a[19] & b[248])^(a[18] & b[249])^(a[17] & b[250])^(a[16] & b[251])^(a[15] & b[252])^(a[14] & b[253])^(a[13] & b[254])^(a[12] & b[255])^(a[11] & b[256])^(a[10] & b[257])^(a[9] & b[258])^(a[8] & b[259])^(a[7] & b[260])^(a[6] & b[261])^(a[5] & b[262])^(a[4] & b[263])^(a[3] & b[264])^(a[2] & b[265])^(a[1] & b[266])^(a[0] & b[267]);
assign y[268] = (a[268] & b[0])^(a[267] & b[1])^(a[266] & b[2])^(a[265] & b[3])^(a[264] & b[4])^(a[263] & b[5])^(a[262] & b[6])^(a[261] & b[7])^(a[260] & b[8])^(a[259] & b[9])^(a[258] & b[10])^(a[257] & b[11])^(a[256] & b[12])^(a[255] & b[13])^(a[254] & b[14])^(a[253] & b[15])^(a[252] & b[16])^(a[251] & b[17])^(a[250] & b[18])^(a[249] & b[19])^(a[248] & b[20])^(a[247] & b[21])^(a[246] & b[22])^(a[245] & b[23])^(a[244] & b[24])^(a[243] & b[25])^(a[242] & b[26])^(a[241] & b[27])^(a[240] & b[28])^(a[239] & b[29])^(a[238] & b[30])^(a[237] & b[31])^(a[236] & b[32])^(a[235] & b[33])^(a[234] & b[34])^(a[233] & b[35])^(a[232] & b[36])^(a[231] & b[37])^(a[230] & b[38])^(a[229] & b[39])^(a[228] & b[40])^(a[227] & b[41])^(a[226] & b[42])^(a[225] & b[43])^(a[224] & b[44])^(a[223] & b[45])^(a[222] & b[46])^(a[221] & b[47])^(a[220] & b[48])^(a[219] & b[49])^(a[218] & b[50])^(a[217] & b[51])^(a[216] & b[52])^(a[215] & b[53])^(a[214] & b[54])^(a[213] & b[55])^(a[212] & b[56])^(a[211] & b[57])^(a[210] & b[58])^(a[209] & b[59])^(a[208] & b[60])^(a[207] & b[61])^(a[206] & b[62])^(a[205] & b[63])^(a[204] & b[64])^(a[203] & b[65])^(a[202] & b[66])^(a[201] & b[67])^(a[200] & b[68])^(a[199] & b[69])^(a[198] & b[70])^(a[197] & b[71])^(a[196] & b[72])^(a[195] & b[73])^(a[194] & b[74])^(a[193] & b[75])^(a[192] & b[76])^(a[191] & b[77])^(a[190] & b[78])^(a[189] & b[79])^(a[188] & b[80])^(a[187] & b[81])^(a[186] & b[82])^(a[185] & b[83])^(a[184] & b[84])^(a[183] & b[85])^(a[182] & b[86])^(a[181] & b[87])^(a[180] & b[88])^(a[179] & b[89])^(a[178] & b[90])^(a[177] & b[91])^(a[176] & b[92])^(a[175] & b[93])^(a[174] & b[94])^(a[173] & b[95])^(a[172] & b[96])^(a[171] & b[97])^(a[170] & b[98])^(a[169] & b[99])^(a[168] & b[100])^(a[167] & b[101])^(a[166] & b[102])^(a[165] & b[103])^(a[164] & b[104])^(a[163] & b[105])^(a[162] & b[106])^(a[161] & b[107])^(a[160] & b[108])^(a[159] & b[109])^(a[158] & b[110])^(a[157] & b[111])^(a[156] & b[112])^(a[155] & b[113])^(a[154] & b[114])^(a[153] & b[115])^(a[152] & b[116])^(a[151] & b[117])^(a[150] & b[118])^(a[149] & b[119])^(a[148] & b[120])^(a[147] & b[121])^(a[146] & b[122])^(a[145] & b[123])^(a[144] & b[124])^(a[143] & b[125])^(a[142] & b[126])^(a[141] & b[127])^(a[140] & b[128])^(a[139] & b[129])^(a[138] & b[130])^(a[137] & b[131])^(a[136] & b[132])^(a[135] & b[133])^(a[134] & b[134])^(a[133] & b[135])^(a[132] & b[136])^(a[131] & b[137])^(a[130] & b[138])^(a[129] & b[139])^(a[128] & b[140])^(a[127] & b[141])^(a[126] & b[142])^(a[125] & b[143])^(a[124] & b[144])^(a[123] & b[145])^(a[122] & b[146])^(a[121] & b[147])^(a[120] & b[148])^(a[119] & b[149])^(a[118] & b[150])^(a[117] & b[151])^(a[116] & b[152])^(a[115] & b[153])^(a[114] & b[154])^(a[113] & b[155])^(a[112] & b[156])^(a[111] & b[157])^(a[110] & b[158])^(a[109] & b[159])^(a[108] & b[160])^(a[107] & b[161])^(a[106] & b[162])^(a[105] & b[163])^(a[104] & b[164])^(a[103] & b[165])^(a[102] & b[166])^(a[101] & b[167])^(a[100] & b[168])^(a[99] & b[169])^(a[98] & b[170])^(a[97] & b[171])^(a[96] & b[172])^(a[95] & b[173])^(a[94] & b[174])^(a[93] & b[175])^(a[92] & b[176])^(a[91] & b[177])^(a[90] & b[178])^(a[89] & b[179])^(a[88] & b[180])^(a[87] & b[181])^(a[86] & b[182])^(a[85] & b[183])^(a[84] & b[184])^(a[83] & b[185])^(a[82] & b[186])^(a[81] & b[187])^(a[80] & b[188])^(a[79] & b[189])^(a[78] & b[190])^(a[77] & b[191])^(a[76] & b[192])^(a[75] & b[193])^(a[74] & b[194])^(a[73] & b[195])^(a[72] & b[196])^(a[71] & b[197])^(a[70] & b[198])^(a[69] & b[199])^(a[68] & b[200])^(a[67] & b[201])^(a[66] & b[202])^(a[65] & b[203])^(a[64] & b[204])^(a[63] & b[205])^(a[62] & b[206])^(a[61] & b[207])^(a[60] & b[208])^(a[59] & b[209])^(a[58] & b[210])^(a[57] & b[211])^(a[56] & b[212])^(a[55] & b[213])^(a[54] & b[214])^(a[53] & b[215])^(a[52] & b[216])^(a[51] & b[217])^(a[50] & b[218])^(a[49] & b[219])^(a[48] & b[220])^(a[47] & b[221])^(a[46] & b[222])^(a[45] & b[223])^(a[44] & b[224])^(a[43] & b[225])^(a[42] & b[226])^(a[41] & b[227])^(a[40] & b[228])^(a[39] & b[229])^(a[38] & b[230])^(a[37] & b[231])^(a[36] & b[232])^(a[35] & b[233])^(a[34] & b[234])^(a[33] & b[235])^(a[32] & b[236])^(a[31] & b[237])^(a[30] & b[238])^(a[29] & b[239])^(a[28] & b[240])^(a[27] & b[241])^(a[26] & b[242])^(a[25] & b[243])^(a[24] & b[244])^(a[23] & b[245])^(a[22] & b[246])^(a[21] & b[247])^(a[20] & b[248])^(a[19] & b[249])^(a[18] & b[250])^(a[17] & b[251])^(a[16] & b[252])^(a[15] & b[253])^(a[14] & b[254])^(a[13] & b[255])^(a[12] & b[256])^(a[11] & b[257])^(a[10] & b[258])^(a[9] & b[259])^(a[8] & b[260])^(a[7] & b[261])^(a[6] & b[262])^(a[5] & b[263])^(a[4] & b[264])^(a[3] & b[265])^(a[2] & b[266])^(a[1] & b[267])^(a[0] & b[268]);
assign y[269] = (a[269] & b[0])^(a[268] & b[1])^(a[267] & b[2])^(a[266] & b[3])^(a[265] & b[4])^(a[264] & b[5])^(a[263] & b[6])^(a[262] & b[7])^(a[261] & b[8])^(a[260] & b[9])^(a[259] & b[10])^(a[258] & b[11])^(a[257] & b[12])^(a[256] & b[13])^(a[255] & b[14])^(a[254] & b[15])^(a[253] & b[16])^(a[252] & b[17])^(a[251] & b[18])^(a[250] & b[19])^(a[249] & b[20])^(a[248] & b[21])^(a[247] & b[22])^(a[246] & b[23])^(a[245] & b[24])^(a[244] & b[25])^(a[243] & b[26])^(a[242] & b[27])^(a[241] & b[28])^(a[240] & b[29])^(a[239] & b[30])^(a[238] & b[31])^(a[237] & b[32])^(a[236] & b[33])^(a[235] & b[34])^(a[234] & b[35])^(a[233] & b[36])^(a[232] & b[37])^(a[231] & b[38])^(a[230] & b[39])^(a[229] & b[40])^(a[228] & b[41])^(a[227] & b[42])^(a[226] & b[43])^(a[225] & b[44])^(a[224] & b[45])^(a[223] & b[46])^(a[222] & b[47])^(a[221] & b[48])^(a[220] & b[49])^(a[219] & b[50])^(a[218] & b[51])^(a[217] & b[52])^(a[216] & b[53])^(a[215] & b[54])^(a[214] & b[55])^(a[213] & b[56])^(a[212] & b[57])^(a[211] & b[58])^(a[210] & b[59])^(a[209] & b[60])^(a[208] & b[61])^(a[207] & b[62])^(a[206] & b[63])^(a[205] & b[64])^(a[204] & b[65])^(a[203] & b[66])^(a[202] & b[67])^(a[201] & b[68])^(a[200] & b[69])^(a[199] & b[70])^(a[198] & b[71])^(a[197] & b[72])^(a[196] & b[73])^(a[195] & b[74])^(a[194] & b[75])^(a[193] & b[76])^(a[192] & b[77])^(a[191] & b[78])^(a[190] & b[79])^(a[189] & b[80])^(a[188] & b[81])^(a[187] & b[82])^(a[186] & b[83])^(a[185] & b[84])^(a[184] & b[85])^(a[183] & b[86])^(a[182] & b[87])^(a[181] & b[88])^(a[180] & b[89])^(a[179] & b[90])^(a[178] & b[91])^(a[177] & b[92])^(a[176] & b[93])^(a[175] & b[94])^(a[174] & b[95])^(a[173] & b[96])^(a[172] & b[97])^(a[171] & b[98])^(a[170] & b[99])^(a[169] & b[100])^(a[168] & b[101])^(a[167] & b[102])^(a[166] & b[103])^(a[165] & b[104])^(a[164] & b[105])^(a[163] & b[106])^(a[162] & b[107])^(a[161] & b[108])^(a[160] & b[109])^(a[159] & b[110])^(a[158] & b[111])^(a[157] & b[112])^(a[156] & b[113])^(a[155] & b[114])^(a[154] & b[115])^(a[153] & b[116])^(a[152] & b[117])^(a[151] & b[118])^(a[150] & b[119])^(a[149] & b[120])^(a[148] & b[121])^(a[147] & b[122])^(a[146] & b[123])^(a[145] & b[124])^(a[144] & b[125])^(a[143] & b[126])^(a[142] & b[127])^(a[141] & b[128])^(a[140] & b[129])^(a[139] & b[130])^(a[138] & b[131])^(a[137] & b[132])^(a[136] & b[133])^(a[135] & b[134])^(a[134] & b[135])^(a[133] & b[136])^(a[132] & b[137])^(a[131] & b[138])^(a[130] & b[139])^(a[129] & b[140])^(a[128] & b[141])^(a[127] & b[142])^(a[126] & b[143])^(a[125] & b[144])^(a[124] & b[145])^(a[123] & b[146])^(a[122] & b[147])^(a[121] & b[148])^(a[120] & b[149])^(a[119] & b[150])^(a[118] & b[151])^(a[117] & b[152])^(a[116] & b[153])^(a[115] & b[154])^(a[114] & b[155])^(a[113] & b[156])^(a[112] & b[157])^(a[111] & b[158])^(a[110] & b[159])^(a[109] & b[160])^(a[108] & b[161])^(a[107] & b[162])^(a[106] & b[163])^(a[105] & b[164])^(a[104] & b[165])^(a[103] & b[166])^(a[102] & b[167])^(a[101] & b[168])^(a[100] & b[169])^(a[99] & b[170])^(a[98] & b[171])^(a[97] & b[172])^(a[96] & b[173])^(a[95] & b[174])^(a[94] & b[175])^(a[93] & b[176])^(a[92] & b[177])^(a[91] & b[178])^(a[90] & b[179])^(a[89] & b[180])^(a[88] & b[181])^(a[87] & b[182])^(a[86] & b[183])^(a[85] & b[184])^(a[84] & b[185])^(a[83] & b[186])^(a[82] & b[187])^(a[81] & b[188])^(a[80] & b[189])^(a[79] & b[190])^(a[78] & b[191])^(a[77] & b[192])^(a[76] & b[193])^(a[75] & b[194])^(a[74] & b[195])^(a[73] & b[196])^(a[72] & b[197])^(a[71] & b[198])^(a[70] & b[199])^(a[69] & b[200])^(a[68] & b[201])^(a[67] & b[202])^(a[66] & b[203])^(a[65] & b[204])^(a[64] & b[205])^(a[63] & b[206])^(a[62] & b[207])^(a[61] & b[208])^(a[60] & b[209])^(a[59] & b[210])^(a[58] & b[211])^(a[57] & b[212])^(a[56] & b[213])^(a[55] & b[214])^(a[54] & b[215])^(a[53] & b[216])^(a[52] & b[217])^(a[51] & b[218])^(a[50] & b[219])^(a[49] & b[220])^(a[48] & b[221])^(a[47] & b[222])^(a[46] & b[223])^(a[45] & b[224])^(a[44] & b[225])^(a[43] & b[226])^(a[42] & b[227])^(a[41] & b[228])^(a[40] & b[229])^(a[39] & b[230])^(a[38] & b[231])^(a[37] & b[232])^(a[36] & b[233])^(a[35] & b[234])^(a[34] & b[235])^(a[33] & b[236])^(a[32] & b[237])^(a[31] & b[238])^(a[30] & b[239])^(a[29] & b[240])^(a[28] & b[241])^(a[27] & b[242])^(a[26] & b[243])^(a[25] & b[244])^(a[24] & b[245])^(a[23] & b[246])^(a[22] & b[247])^(a[21] & b[248])^(a[20] & b[249])^(a[19] & b[250])^(a[18] & b[251])^(a[17] & b[252])^(a[16] & b[253])^(a[15] & b[254])^(a[14] & b[255])^(a[13] & b[256])^(a[12] & b[257])^(a[11] & b[258])^(a[10] & b[259])^(a[9] & b[260])^(a[8] & b[261])^(a[7] & b[262])^(a[6] & b[263])^(a[5] & b[264])^(a[4] & b[265])^(a[3] & b[266])^(a[2] & b[267])^(a[1] & b[268])^(a[0] & b[269]);
assign y[270] = (a[270] & b[0])^(a[269] & b[1])^(a[268] & b[2])^(a[267] & b[3])^(a[266] & b[4])^(a[265] & b[5])^(a[264] & b[6])^(a[263] & b[7])^(a[262] & b[8])^(a[261] & b[9])^(a[260] & b[10])^(a[259] & b[11])^(a[258] & b[12])^(a[257] & b[13])^(a[256] & b[14])^(a[255] & b[15])^(a[254] & b[16])^(a[253] & b[17])^(a[252] & b[18])^(a[251] & b[19])^(a[250] & b[20])^(a[249] & b[21])^(a[248] & b[22])^(a[247] & b[23])^(a[246] & b[24])^(a[245] & b[25])^(a[244] & b[26])^(a[243] & b[27])^(a[242] & b[28])^(a[241] & b[29])^(a[240] & b[30])^(a[239] & b[31])^(a[238] & b[32])^(a[237] & b[33])^(a[236] & b[34])^(a[235] & b[35])^(a[234] & b[36])^(a[233] & b[37])^(a[232] & b[38])^(a[231] & b[39])^(a[230] & b[40])^(a[229] & b[41])^(a[228] & b[42])^(a[227] & b[43])^(a[226] & b[44])^(a[225] & b[45])^(a[224] & b[46])^(a[223] & b[47])^(a[222] & b[48])^(a[221] & b[49])^(a[220] & b[50])^(a[219] & b[51])^(a[218] & b[52])^(a[217] & b[53])^(a[216] & b[54])^(a[215] & b[55])^(a[214] & b[56])^(a[213] & b[57])^(a[212] & b[58])^(a[211] & b[59])^(a[210] & b[60])^(a[209] & b[61])^(a[208] & b[62])^(a[207] & b[63])^(a[206] & b[64])^(a[205] & b[65])^(a[204] & b[66])^(a[203] & b[67])^(a[202] & b[68])^(a[201] & b[69])^(a[200] & b[70])^(a[199] & b[71])^(a[198] & b[72])^(a[197] & b[73])^(a[196] & b[74])^(a[195] & b[75])^(a[194] & b[76])^(a[193] & b[77])^(a[192] & b[78])^(a[191] & b[79])^(a[190] & b[80])^(a[189] & b[81])^(a[188] & b[82])^(a[187] & b[83])^(a[186] & b[84])^(a[185] & b[85])^(a[184] & b[86])^(a[183] & b[87])^(a[182] & b[88])^(a[181] & b[89])^(a[180] & b[90])^(a[179] & b[91])^(a[178] & b[92])^(a[177] & b[93])^(a[176] & b[94])^(a[175] & b[95])^(a[174] & b[96])^(a[173] & b[97])^(a[172] & b[98])^(a[171] & b[99])^(a[170] & b[100])^(a[169] & b[101])^(a[168] & b[102])^(a[167] & b[103])^(a[166] & b[104])^(a[165] & b[105])^(a[164] & b[106])^(a[163] & b[107])^(a[162] & b[108])^(a[161] & b[109])^(a[160] & b[110])^(a[159] & b[111])^(a[158] & b[112])^(a[157] & b[113])^(a[156] & b[114])^(a[155] & b[115])^(a[154] & b[116])^(a[153] & b[117])^(a[152] & b[118])^(a[151] & b[119])^(a[150] & b[120])^(a[149] & b[121])^(a[148] & b[122])^(a[147] & b[123])^(a[146] & b[124])^(a[145] & b[125])^(a[144] & b[126])^(a[143] & b[127])^(a[142] & b[128])^(a[141] & b[129])^(a[140] & b[130])^(a[139] & b[131])^(a[138] & b[132])^(a[137] & b[133])^(a[136] & b[134])^(a[135] & b[135])^(a[134] & b[136])^(a[133] & b[137])^(a[132] & b[138])^(a[131] & b[139])^(a[130] & b[140])^(a[129] & b[141])^(a[128] & b[142])^(a[127] & b[143])^(a[126] & b[144])^(a[125] & b[145])^(a[124] & b[146])^(a[123] & b[147])^(a[122] & b[148])^(a[121] & b[149])^(a[120] & b[150])^(a[119] & b[151])^(a[118] & b[152])^(a[117] & b[153])^(a[116] & b[154])^(a[115] & b[155])^(a[114] & b[156])^(a[113] & b[157])^(a[112] & b[158])^(a[111] & b[159])^(a[110] & b[160])^(a[109] & b[161])^(a[108] & b[162])^(a[107] & b[163])^(a[106] & b[164])^(a[105] & b[165])^(a[104] & b[166])^(a[103] & b[167])^(a[102] & b[168])^(a[101] & b[169])^(a[100] & b[170])^(a[99] & b[171])^(a[98] & b[172])^(a[97] & b[173])^(a[96] & b[174])^(a[95] & b[175])^(a[94] & b[176])^(a[93] & b[177])^(a[92] & b[178])^(a[91] & b[179])^(a[90] & b[180])^(a[89] & b[181])^(a[88] & b[182])^(a[87] & b[183])^(a[86] & b[184])^(a[85] & b[185])^(a[84] & b[186])^(a[83] & b[187])^(a[82] & b[188])^(a[81] & b[189])^(a[80] & b[190])^(a[79] & b[191])^(a[78] & b[192])^(a[77] & b[193])^(a[76] & b[194])^(a[75] & b[195])^(a[74] & b[196])^(a[73] & b[197])^(a[72] & b[198])^(a[71] & b[199])^(a[70] & b[200])^(a[69] & b[201])^(a[68] & b[202])^(a[67] & b[203])^(a[66] & b[204])^(a[65] & b[205])^(a[64] & b[206])^(a[63] & b[207])^(a[62] & b[208])^(a[61] & b[209])^(a[60] & b[210])^(a[59] & b[211])^(a[58] & b[212])^(a[57] & b[213])^(a[56] & b[214])^(a[55] & b[215])^(a[54] & b[216])^(a[53] & b[217])^(a[52] & b[218])^(a[51] & b[219])^(a[50] & b[220])^(a[49] & b[221])^(a[48] & b[222])^(a[47] & b[223])^(a[46] & b[224])^(a[45] & b[225])^(a[44] & b[226])^(a[43] & b[227])^(a[42] & b[228])^(a[41] & b[229])^(a[40] & b[230])^(a[39] & b[231])^(a[38] & b[232])^(a[37] & b[233])^(a[36] & b[234])^(a[35] & b[235])^(a[34] & b[236])^(a[33] & b[237])^(a[32] & b[238])^(a[31] & b[239])^(a[30] & b[240])^(a[29] & b[241])^(a[28] & b[242])^(a[27] & b[243])^(a[26] & b[244])^(a[25] & b[245])^(a[24] & b[246])^(a[23] & b[247])^(a[22] & b[248])^(a[21] & b[249])^(a[20] & b[250])^(a[19] & b[251])^(a[18] & b[252])^(a[17] & b[253])^(a[16] & b[254])^(a[15] & b[255])^(a[14] & b[256])^(a[13] & b[257])^(a[12] & b[258])^(a[11] & b[259])^(a[10] & b[260])^(a[9] & b[261])^(a[8] & b[262])^(a[7] & b[263])^(a[6] & b[264])^(a[5] & b[265])^(a[4] & b[266])^(a[3] & b[267])^(a[2] & b[268])^(a[1] & b[269])^(a[0] & b[270]);
assign y[271] = (a[271] & b[0])^(a[270] & b[1])^(a[269] & b[2])^(a[268] & b[3])^(a[267] & b[4])^(a[266] & b[5])^(a[265] & b[6])^(a[264] & b[7])^(a[263] & b[8])^(a[262] & b[9])^(a[261] & b[10])^(a[260] & b[11])^(a[259] & b[12])^(a[258] & b[13])^(a[257] & b[14])^(a[256] & b[15])^(a[255] & b[16])^(a[254] & b[17])^(a[253] & b[18])^(a[252] & b[19])^(a[251] & b[20])^(a[250] & b[21])^(a[249] & b[22])^(a[248] & b[23])^(a[247] & b[24])^(a[246] & b[25])^(a[245] & b[26])^(a[244] & b[27])^(a[243] & b[28])^(a[242] & b[29])^(a[241] & b[30])^(a[240] & b[31])^(a[239] & b[32])^(a[238] & b[33])^(a[237] & b[34])^(a[236] & b[35])^(a[235] & b[36])^(a[234] & b[37])^(a[233] & b[38])^(a[232] & b[39])^(a[231] & b[40])^(a[230] & b[41])^(a[229] & b[42])^(a[228] & b[43])^(a[227] & b[44])^(a[226] & b[45])^(a[225] & b[46])^(a[224] & b[47])^(a[223] & b[48])^(a[222] & b[49])^(a[221] & b[50])^(a[220] & b[51])^(a[219] & b[52])^(a[218] & b[53])^(a[217] & b[54])^(a[216] & b[55])^(a[215] & b[56])^(a[214] & b[57])^(a[213] & b[58])^(a[212] & b[59])^(a[211] & b[60])^(a[210] & b[61])^(a[209] & b[62])^(a[208] & b[63])^(a[207] & b[64])^(a[206] & b[65])^(a[205] & b[66])^(a[204] & b[67])^(a[203] & b[68])^(a[202] & b[69])^(a[201] & b[70])^(a[200] & b[71])^(a[199] & b[72])^(a[198] & b[73])^(a[197] & b[74])^(a[196] & b[75])^(a[195] & b[76])^(a[194] & b[77])^(a[193] & b[78])^(a[192] & b[79])^(a[191] & b[80])^(a[190] & b[81])^(a[189] & b[82])^(a[188] & b[83])^(a[187] & b[84])^(a[186] & b[85])^(a[185] & b[86])^(a[184] & b[87])^(a[183] & b[88])^(a[182] & b[89])^(a[181] & b[90])^(a[180] & b[91])^(a[179] & b[92])^(a[178] & b[93])^(a[177] & b[94])^(a[176] & b[95])^(a[175] & b[96])^(a[174] & b[97])^(a[173] & b[98])^(a[172] & b[99])^(a[171] & b[100])^(a[170] & b[101])^(a[169] & b[102])^(a[168] & b[103])^(a[167] & b[104])^(a[166] & b[105])^(a[165] & b[106])^(a[164] & b[107])^(a[163] & b[108])^(a[162] & b[109])^(a[161] & b[110])^(a[160] & b[111])^(a[159] & b[112])^(a[158] & b[113])^(a[157] & b[114])^(a[156] & b[115])^(a[155] & b[116])^(a[154] & b[117])^(a[153] & b[118])^(a[152] & b[119])^(a[151] & b[120])^(a[150] & b[121])^(a[149] & b[122])^(a[148] & b[123])^(a[147] & b[124])^(a[146] & b[125])^(a[145] & b[126])^(a[144] & b[127])^(a[143] & b[128])^(a[142] & b[129])^(a[141] & b[130])^(a[140] & b[131])^(a[139] & b[132])^(a[138] & b[133])^(a[137] & b[134])^(a[136] & b[135])^(a[135] & b[136])^(a[134] & b[137])^(a[133] & b[138])^(a[132] & b[139])^(a[131] & b[140])^(a[130] & b[141])^(a[129] & b[142])^(a[128] & b[143])^(a[127] & b[144])^(a[126] & b[145])^(a[125] & b[146])^(a[124] & b[147])^(a[123] & b[148])^(a[122] & b[149])^(a[121] & b[150])^(a[120] & b[151])^(a[119] & b[152])^(a[118] & b[153])^(a[117] & b[154])^(a[116] & b[155])^(a[115] & b[156])^(a[114] & b[157])^(a[113] & b[158])^(a[112] & b[159])^(a[111] & b[160])^(a[110] & b[161])^(a[109] & b[162])^(a[108] & b[163])^(a[107] & b[164])^(a[106] & b[165])^(a[105] & b[166])^(a[104] & b[167])^(a[103] & b[168])^(a[102] & b[169])^(a[101] & b[170])^(a[100] & b[171])^(a[99] & b[172])^(a[98] & b[173])^(a[97] & b[174])^(a[96] & b[175])^(a[95] & b[176])^(a[94] & b[177])^(a[93] & b[178])^(a[92] & b[179])^(a[91] & b[180])^(a[90] & b[181])^(a[89] & b[182])^(a[88] & b[183])^(a[87] & b[184])^(a[86] & b[185])^(a[85] & b[186])^(a[84] & b[187])^(a[83] & b[188])^(a[82] & b[189])^(a[81] & b[190])^(a[80] & b[191])^(a[79] & b[192])^(a[78] & b[193])^(a[77] & b[194])^(a[76] & b[195])^(a[75] & b[196])^(a[74] & b[197])^(a[73] & b[198])^(a[72] & b[199])^(a[71] & b[200])^(a[70] & b[201])^(a[69] & b[202])^(a[68] & b[203])^(a[67] & b[204])^(a[66] & b[205])^(a[65] & b[206])^(a[64] & b[207])^(a[63] & b[208])^(a[62] & b[209])^(a[61] & b[210])^(a[60] & b[211])^(a[59] & b[212])^(a[58] & b[213])^(a[57] & b[214])^(a[56] & b[215])^(a[55] & b[216])^(a[54] & b[217])^(a[53] & b[218])^(a[52] & b[219])^(a[51] & b[220])^(a[50] & b[221])^(a[49] & b[222])^(a[48] & b[223])^(a[47] & b[224])^(a[46] & b[225])^(a[45] & b[226])^(a[44] & b[227])^(a[43] & b[228])^(a[42] & b[229])^(a[41] & b[230])^(a[40] & b[231])^(a[39] & b[232])^(a[38] & b[233])^(a[37] & b[234])^(a[36] & b[235])^(a[35] & b[236])^(a[34] & b[237])^(a[33] & b[238])^(a[32] & b[239])^(a[31] & b[240])^(a[30] & b[241])^(a[29] & b[242])^(a[28] & b[243])^(a[27] & b[244])^(a[26] & b[245])^(a[25] & b[246])^(a[24] & b[247])^(a[23] & b[248])^(a[22] & b[249])^(a[21] & b[250])^(a[20] & b[251])^(a[19] & b[252])^(a[18] & b[253])^(a[17] & b[254])^(a[16] & b[255])^(a[15] & b[256])^(a[14] & b[257])^(a[13] & b[258])^(a[12] & b[259])^(a[11] & b[260])^(a[10] & b[261])^(a[9] & b[262])^(a[8] & b[263])^(a[7] & b[264])^(a[6] & b[265])^(a[5] & b[266])^(a[4] & b[267])^(a[3] & b[268])^(a[2] & b[269])^(a[1] & b[270])^(a[0] & b[271]);
assign y[272] = (a[272] & b[0])^(a[271] & b[1])^(a[270] & b[2])^(a[269] & b[3])^(a[268] & b[4])^(a[267] & b[5])^(a[266] & b[6])^(a[265] & b[7])^(a[264] & b[8])^(a[263] & b[9])^(a[262] & b[10])^(a[261] & b[11])^(a[260] & b[12])^(a[259] & b[13])^(a[258] & b[14])^(a[257] & b[15])^(a[256] & b[16])^(a[255] & b[17])^(a[254] & b[18])^(a[253] & b[19])^(a[252] & b[20])^(a[251] & b[21])^(a[250] & b[22])^(a[249] & b[23])^(a[248] & b[24])^(a[247] & b[25])^(a[246] & b[26])^(a[245] & b[27])^(a[244] & b[28])^(a[243] & b[29])^(a[242] & b[30])^(a[241] & b[31])^(a[240] & b[32])^(a[239] & b[33])^(a[238] & b[34])^(a[237] & b[35])^(a[236] & b[36])^(a[235] & b[37])^(a[234] & b[38])^(a[233] & b[39])^(a[232] & b[40])^(a[231] & b[41])^(a[230] & b[42])^(a[229] & b[43])^(a[228] & b[44])^(a[227] & b[45])^(a[226] & b[46])^(a[225] & b[47])^(a[224] & b[48])^(a[223] & b[49])^(a[222] & b[50])^(a[221] & b[51])^(a[220] & b[52])^(a[219] & b[53])^(a[218] & b[54])^(a[217] & b[55])^(a[216] & b[56])^(a[215] & b[57])^(a[214] & b[58])^(a[213] & b[59])^(a[212] & b[60])^(a[211] & b[61])^(a[210] & b[62])^(a[209] & b[63])^(a[208] & b[64])^(a[207] & b[65])^(a[206] & b[66])^(a[205] & b[67])^(a[204] & b[68])^(a[203] & b[69])^(a[202] & b[70])^(a[201] & b[71])^(a[200] & b[72])^(a[199] & b[73])^(a[198] & b[74])^(a[197] & b[75])^(a[196] & b[76])^(a[195] & b[77])^(a[194] & b[78])^(a[193] & b[79])^(a[192] & b[80])^(a[191] & b[81])^(a[190] & b[82])^(a[189] & b[83])^(a[188] & b[84])^(a[187] & b[85])^(a[186] & b[86])^(a[185] & b[87])^(a[184] & b[88])^(a[183] & b[89])^(a[182] & b[90])^(a[181] & b[91])^(a[180] & b[92])^(a[179] & b[93])^(a[178] & b[94])^(a[177] & b[95])^(a[176] & b[96])^(a[175] & b[97])^(a[174] & b[98])^(a[173] & b[99])^(a[172] & b[100])^(a[171] & b[101])^(a[170] & b[102])^(a[169] & b[103])^(a[168] & b[104])^(a[167] & b[105])^(a[166] & b[106])^(a[165] & b[107])^(a[164] & b[108])^(a[163] & b[109])^(a[162] & b[110])^(a[161] & b[111])^(a[160] & b[112])^(a[159] & b[113])^(a[158] & b[114])^(a[157] & b[115])^(a[156] & b[116])^(a[155] & b[117])^(a[154] & b[118])^(a[153] & b[119])^(a[152] & b[120])^(a[151] & b[121])^(a[150] & b[122])^(a[149] & b[123])^(a[148] & b[124])^(a[147] & b[125])^(a[146] & b[126])^(a[145] & b[127])^(a[144] & b[128])^(a[143] & b[129])^(a[142] & b[130])^(a[141] & b[131])^(a[140] & b[132])^(a[139] & b[133])^(a[138] & b[134])^(a[137] & b[135])^(a[136] & b[136])^(a[135] & b[137])^(a[134] & b[138])^(a[133] & b[139])^(a[132] & b[140])^(a[131] & b[141])^(a[130] & b[142])^(a[129] & b[143])^(a[128] & b[144])^(a[127] & b[145])^(a[126] & b[146])^(a[125] & b[147])^(a[124] & b[148])^(a[123] & b[149])^(a[122] & b[150])^(a[121] & b[151])^(a[120] & b[152])^(a[119] & b[153])^(a[118] & b[154])^(a[117] & b[155])^(a[116] & b[156])^(a[115] & b[157])^(a[114] & b[158])^(a[113] & b[159])^(a[112] & b[160])^(a[111] & b[161])^(a[110] & b[162])^(a[109] & b[163])^(a[108] & b[164])^(a[107] & b[165])^(a[106] & b[166])^(a[105] & b[167])^(a[104] & b[168])^(a[103] & b[169])^(a[102] & b[170])^(a[101] & b[171])^(a[100] & b[172])^(a[99] & b[173])^(a[98] & b[174])^(a[97] & b[175])^(a[96] & b[176])^(a[95] & b[177])^(a[94] & b[178])^(a[93] & b[179])^(a[92] & b[180])^(a[91] & b[181])^(a[90] & b[182])^(a[89] & b[183])^(a[88] & b[184])^(a[87] & b[185])^(a[86] & b[186])^(a[85] & b[187])^(a[84] & b[188])^(a[83] & b[189])^(a[82] & b[190])^(a[81] & b[191])^(a[80] & b[192])^(a[79] & b[193])^(a[78] & b[194])^(a[77] & b[195])^(a[76] & b[196])^(a[75] & b[197])^(a[74] & b[198])^(a[73] & b[199])^(a[72] & b[200])^(a[71] & b[201])^(a[70] & b[202])^(a[69] & b[203])^(a[68] & b[204])^(a[67] & b[205])^(a[66] & b[206])^(a[65] & b[207])^(a[64] & b[208])^(a[63] & b[209])^(a[62] & b[210])^(a[61] & b[211])^(a[60] & b[212])^(a[59] & b[213])^(a[58] & b[214])^(a[57] & b[215])^(a[56] & b[216])^(a[55] & b[217])^(a[54] & b[218])^(a[53] & b[219])^(a[52] & b[220])^(a[51] & b[221])^(a[50] & b[222])^(a[49] & b[223])^(a[48] & b[224])^(a[47] & b[225])^(a[46] & b[226])^(a[45] & b[227])^(a[44] & b[228])^(a[43] & b[229])^(a[42] & b[230])^(a[41] & b[231])^(a[40] & b[232])^(a[39] & b[233])^(a[38] & b[234])^(a[37] & b[235])^(a[36] & b[236])^(a[35] & b[237])^(a[34] & b[238])^(a[33] & b[239])^(a[32] & b[240])^(a[31] & b[241])^(a[30] & b[242])^(a[29] & b[243])^(a[28] & b[244])^(a[27] & b[245])^(a[26] & b[246])^(a[25] & b[247])^(a[24] & b[248])^(a[23] & b[249])^(a[22] & b[250])^(a[21] & b[251])^(a[20] & b[252])^(a[19] & b[253])^(a[18] & b[254])^(a[17] & b[255])^(a[16] & b[256])^(a[15] & b[257])^(a[14] & b[258])^(a[13] & b[259])^(a[12] & b[260])^(a[11] & b[261])^(a[10] & b[262])^(a[9] & b[263])^(a[8] & b[264])^(a[7] & b[265])^(a[6] & b[266])^(a[5] & b[267])^(a[4] & b[268])^(a[3] & b[269])^(a[2] & b[270])^(a[1] & b[271])^(a[0] & b[272]);
assign y[273] = (a[273] & b[0])^(a[272] & b[1])^(a[271] & b[2])^(a[270] & b[3])^(a[269] & b[4])^(a[268] & b[5])^(a[267] & b[6])^(a[266] & b[7])^(a[265] & b[8])^(a[264] & b[9])^(a[263] & b[10])^(a[262] & b[11])^(a[261] & b[12])^(a[260] & b[13])^(a[259] & b[14])^(a[258] & b[15])^(a[257] & b[16])^(a[256] & b[17])^(a[255] & b[18])^(a[254] & b[19])^(a[253] & b[20])^(a[252] & b[21])^(a[251] & b[22])^(a[250] & b[23])^(a[249] & b[24])^(a[248] & b[25])^(a[247] & b[26])^(a[246] & b[27])^(a[245] & b[28])^(a[244] & b[29])^(a[243] & b[30])^(a[242] & b[31])^(a[241] & b[32])^(a[240] & b[33])^(a[239] & b[34])^(a[238] & b[35])^(a[237] & b[36])^(a[236] & b[37])^(a[235] & b[38])^(a[234] & b[39])^(a[233] & b[40])^(a[232] & b[41])^(a[231] & b[42])^(a[230] & b[43])^(a[229] & b[44])^(a[228] & b[45])^(a[227] & b[46])^(a[226] & b[47])^(a[225] & b[48])^(a[224] & b[49])^(a[223] & b[50])^(a[222] & b[51])^(a[221] & b[52])^(a[220] & b[53])^(a[219] & b[54])^(a[218] & b[55])^(a[217] & b[56])^(a[216] & b[57])^(a[215] & b[58])^(a[214] & b[59])^(a[213] & b[60])^(a[212] & b[61])^(a[211] & b[62])^(a[210] & b[63])^(a[209] & b[64])^(a[208] & b[65])^(a[207] & b[66])^(a[206] & b[67])^(a[205] & b[68])^(a[204] & b[69])^(a[203] & b[70])^(a[202] & b[71])^(a[201] & b[72])^(a[200] & b[73])^(a[199] & b[74])^(a[198] & b[75])^(a[197] & b[76])^(a[196] & b[77])^(a[195] & b[78])^(a[194] & b[79])^(a[193] & b[80])^(a[192] & b[81])^(a[191] & b[82])^(a[190] & b[83])^(a[189] & b[84])^(a[188] & b[85])^(a[187] & b[86])^(a[186] & b[87])^(a[185] & b[88])^(a[184] & b[89])^(a[183] & b[90])^(a[182] & b[91])^(a[181] & b[92])^(a[180] & b[93])^(a[179] & b[94])^(a[178] & b[95])^(a[177] & b[96])^(a[176] & b[97])^(a[175] & b[98])^(a[174] & b[99])^(a[173] & b[100])^(a[172] & b[101])^(a[171] & b[102])^(a[170] & b[103])^(a[169] & b[104])^(a[168] & b[105])^(a[167] & b[106])^(a[166] & b[107])^(a[165] & b[108])^(a[164] & b[109])^(a[163] & b[110])^(a[162] & b[111])^(a[161] & b[112])^(a[160] & b[113])^(a[159] & b[114])^(a[158] & b[115])^(a[157] & b[116])^(a[156] & b[117])^(a[155] & b[118])^(a[154] & b[119])^(a[153] & b[120])^(a[152] & b[121])^(a[151] & b[122])^(a[150] & b[123])^(a[149] & b[124])^(a[148] & b[125])^(a[147] & b[126])^(a[146] & b[127])^(a[145] & b[128])^(a[144] & b[129])^(a[143] & b[130])^(a[142] & b[131])^(a[141] & b[132])^(a[140] & b[133])^(a[139] & b[134])^(a[138] & b[135])^(a[137] & b[136])^(a[136] & b[137])^(a[135] & b[138])^(a[134] & b[139])^(a[133] & b[140])^(a[132] & b[141])^(a[131] & b[142])^(a[130] & b[143])^(a[129] & b[144])^(a[128] & b[145])^(a[127] & b[146])^(a[126] & b[147])^(a[125] & b[148])^(a[124] & b[149])^(a[123] & b[150])^(a[122] & b[151])^(a[121] & b[152])^(a[120] & b[153])^(a[119] & b[154])^(a[118] & b[155])^(a[117] & b[156])^(a[116] & b[157])^(a[115] & b[158])^(a[114] & b[159])^(a[113] & b[160])^(a[112] & b[161])^(a[111] & b[162])^(a[110] & b[163])^(a[109] & b[164])^(a[108] & b[165])^(a[107] & b[166])^(a[106] & b[167])^(a[105] & b[168])^(a[104] & b[169])^(a[103] & b[170])^(a[102] & b[171])^(a[101] & b[172])^(a[100] & b[173])^(a[99] & b[174])^(a[98] & b[175])^(a[97] & b[176])^(a[96] & b[177])^(a[95] & b[178])^(a[94] & b[179])^(a[93] & b[180])^(a[92] & b[181])^(a[91] & b[182])^(a[90] & b[183])^(a[89] & b[184])^(a[88] & b[185])^(a[87] & b[186])^(a[86] & b[187])^(a[85] & b[188])^(a[84] & b[189])^(a[83] & b[190])^(a[82] & b[191])^(a[81] & b[192])^(a[80] & b[193])^(a[79] & b[194])^(a[78] & b[195])^(a[77] & b[196])^(a[76] & b[197])^(a[75] & b[198])^(a[74] & b[199])^(a[73] & b[200])^(a[72] & b[201])^(a[71] & b[202])^(a[70] & b[203])^(a[69] & b[204])^(a[68] & b[205])^(a[67] & b[206])^(a[66] & b[207])^(a[65] & b[208])^(a[64] & b[209])^(a[63] & b[210])^(a[62] & b[211])^(a[61] & b[212])^(a[60] & b[213])^(a[59] & b[214])^(a[58] & b[215])^(a[57] & b[216])^(a[56] & b[217])^(a[55] & b[218])^(a[54] & b[219])^(a[53] & b[220])^(a[52] & b[221])^(a[51] & b[222])^(a[50] & b[223])^(a[49] & b[224])^(a[48] & b[225])^(a[47] & b[226])^(a[46] & b[227])^(a[45] & b[228])^(a[44] & b[229])^(a[43] & b[230])^(a[42] & b[231])^(a[41] & b[232])^(a[40] & b[233])^(a[39] & b[234])^(a[38] & b[235])^(a[37] & b[236])^(a[36] & b[237])^(a[35] & b[238])^(a[34] & b[239])^(a[33] & b[240])^(a[32] & b[241])^(a[31] & b[242])^(a[30] & b[243])^(a[29] & b[244])^(a[28] & b[245])^(a[27] & b[246])^(a[26] & b[247])^(a[25] & b[248])^(a[24] & b[249])^(a[23] & b[250])^(a[22] & b[251])^(a[21] & b[252])^(a[20] & b[253])^(a[19] & b[254])^(a[18] & b[255])^(a[17] & b[256])^(a[16] & b[257])^(a[15] & b[258])^(a[14] & b[259])^(a[13] & b[260])^(a[12] & b[261])^(a[11] & b[262])^(a[10] & b[263])^(a[9] & b[264])^(a[8] & b[265])^(a[7] & b[266])^(a[6] & b[267])^(a[5] & b[268])^(a[4] & b[269])^(a[3] & b[270])^(a[2] & b[271])^(a[1] & b[272])^(a[0] & b[273]);
assign y[274] = (a[274] & b[0])^(a[273] & b[1])^(a[272] & b[2])^(a[271] & b[3])^(a[270] & b[4])^(a[269] & b[5])^(a[268] & b[6])^(a[267] & b[7])^(a[266] & b[8])^(a[265] & b[9])^(a[264] & b[10])^(a[263] & b[11])^(a[262] & b[12])^(a[261] & b[13])^(a[260] & b[14])^(a[259] & b[15])^(a[258] & b[16])^(a[257] & b[17])^(a[256] & b[18])^(a[255] & b[19])^(a[254] & b[20])^(a[253] & b[21])^(a[252] & b[22])^(a[251] & b[23])^(a[250] & b[24])^(a[249] & b[25])^(a[248] & b[26])^(a[247] & b[27])^(a[246] & b[28])^(a[245] & b[29])^(a[244] & b[30])^(a[243] & b[31])^(a[242] & b[32])^(a[241] & b[33])^(a[240] & b[34])^(a[239] & b[35])^(a[238] & b[36])^(a[237] & b[37])^(a[236] & b[38])^(a[235] & b[39])^(a[234] & b[40])^(a[233] & b[41])^(a[232] & b[42])^(a[231] & b[43])^(a[230] & b[44])^(a[229] & b[45])^(a[228] & b[46])^(a[227] & b[47])^(a[226] & b[48])^(a[225] & b[49])^(a[224] & b[50])^(a[223] & b[51])^(a[222] & b[52])^(a[221] & b[53])^(a[220] & b[54])^(a[219] & b[55])^(a[218] & b[56])^(a[217] & b[57])^(a[216] & b[58])^(a[215] & b[59])^(a[214] & b[60])^(a[213] & b[61])^(a[212] & b[62])^(a[211] & b[63])^(a[210] & b[64])^(a[209] & b[65])^(a[208] & b[66])^(a[207] & b[67])^(a[206] & b[68])^(a[205] & b[69])^(a[204] & b[70])^(a[203] & b[71])^(a[202] & b[72])^(a[201] & b[73])^(a[200] & b[74])^(a[199] & b[75])^(a[198] & b[76])^(a[197] & b[77])^(a[196] & b[78])^(a[195] & b[79])^(a[194] & b[80])^(a[193] & b[81])^(a[192] & b[82])^(a[191] & b[83])^(a[190] & b[84])^(a[189] & b[85])^(a[188] & b[86])^(a[187] & b[87])^(a[186] & b[88])^(a[185] & b[89])^(a[184] & b[90])^(a[183] & b[91])^(a[182] & b[92])^(a[181] & b[93])^(a[180] & b[94])^(a[179] & b[95])^(a[178] & b[96])^(a[177] & b[97])^(a[176] & b[98])^(a[175] & b[99])^(a[174] & b[100])^(a[173] & b[101])^(a[172] & b[102])^(a[171] & b[103])^(a[170] & b[104])^(a[169] & b[105])^(a[168] & b[106])^(a[167] & b[107])^(a[166] & b[108])^(a[165] & b[109])^(a[164] & b[110])^(a[163] & b[111])^(a[162] & b[112])^(a[161] & b[113])^(a[160] & b[114])^(a[159] & b[115])^(a[158] & b[116])^(a[157] & b[117])^(a[156] & b[118])^(a[155] & b[119])^(a[154] & b[120])^(a[153] & b[121])^(a[152] & b[122])^(a[151] & b[123])^(a[150] & b[124])^(a[149] & b[125])^(a[148] & b[126])^(a[147] & b[127])^(a[146] & b[128])^(a[145] & b[129])^(a[144] & b[130])^(a[143] & b[131])^(a[142] & b[132])^(a[141] & b[133])^(a[140] & b[134])^(a[139] & b[135])^(a[138] & b[136])^(a[137] & b[137])^(a[136] & b[138])^(a[135] & b[139])^(a[134] & b[140])^(a[133] & b[141])^(a[132] & b[142])^(a[131] & b[143])^(a[130] & b[144])^(a[129] & b[145])^(a[128] & b[146])^(a[127] & b[147])^(a[126] & b[148])^(a[125] & b[149])^(a[124] & b[150])^(a[123] & b[151])^(a[122] & b[152])^(a[121] & b[153])^(a[120] & b[154])^(a[119] & b[155])^(a[118] & b[156])^(a[117] & b[157])^(a[116] & b[158])^(a[115] & b[159])^(a[114] & b[160])^(a[113] & b[161])^(a[112] & b[162])^(a[111] & b[163])^(a[110] & b[164])^(a[109] & b[165])^(a[108] & b[166])^(a[107] & b[167])^(a[106] & b[168])^(a[105] & b[169])^(a[104] & b[170])^(a[103] & b[171])^(a[102] & b[172])^(a[101] & b[173])^(a[100] & b[174])^(a[99] & b[175])^(a[98] & b[176])^(a[97] & b[177])^(a[96] & b[178])^(a[95] & b[179])^(a[94] & b[180])^(a[93] & b[181])^(a[92] & b[182])^(a[91] & b[183])^(a[90] & b[184])^(a[89] & b[185])^(a[88] & b[186])^(a[87] & b[187])^(a[86] & b[188])^(a[85] & b[189])^(a[84] & b[190])^(a[83] & b[191])^(a[82] & b[192])^(a[81] & b[193])^(a[80] & b[194])^(a[79] & b[195])^(a[78] & b[196])^(a[77] & b[197])^(a[76] & b[198])^(a[75] & b[199])^(a[74] & b[200])^(a[73] & b[201])^(a[72] & b[202])^(a[71] & b[203])^(a[70] & b[204])^(a[69] & b[205])^(a[68] & b[206])^(a[67] & b[207])^(a[66] & b[208])^(a[65] & b[209])^(a[64] & b[210])^(a[63] & b[211])^(a[62] & b[212])^(a[61] & b[213])^(a[60] & b[214])^(a[59] & b[215])^(a[58] & b[216])^(a[57] & b[217])^(a[56] & b[218])^(a[55] & b[219])^(a[54] & b[220])^(a[53] & b[221])^(a[52] & b[222])^(a[51] & b[223])^(a[50] & b[224])^(a[49] & b[225])^(a[48] & b[226])^(a[47] & b[227])^(a[46] & b[228])^(a[45] & b[229])^(a[44] & b[230])^(a[43] & b[231])^(a[42] & b[232])^(a[41] & b[233])^(a[40] & b[234])^(a[39] & b[235])^(a[38] & b[236])^(a[37] & b[237])^(a[36] & b[238])^(a[35] & b[239])^(a[34] & b[240])^(a[33] & b[241])^(a[32] & b[242])^(a[31] & b[243])^(a[30] & b[244])^(a[29] & b[245])^(a[28] & b[246])^(a[27] & b[247])^(a[26] & b[248])^(a[25] & b[249])^(a[24] & b[250])^(a[23] & b[251])^(a[22] & b[252])^(a[21] & b[253])^(a[20] & b[254])^(a[19] & b[255])^(a[18] & b[256])^(a[17] & b[257])^(a[16] & b[258])^(a[15] & b[259])^(a[14] & b[260])^(a[13] & b[261])^(a[12] & b[262])^(a[11] & b[263])^(a[10] & b[264])^(a[9] & b[265])^(a[8] & b[266])^(a[7] & b[267])^(a[6] & b[268])^(a[5] & b[269])^(a[4] & b[270])^(a[3] & b[271])^(a[2] & b[272])^(a[1] & b[273])^(a[0] & b[274]);
assign y[275] = (a[275] & b[0])^(a[274] & b[1])^(a[273] & b[2])^(a[272] & b[3])^(a[271] & b[4])^(a[270] & b[5])^(a[269] & b[6])^(a[268] & b[7])^(a[267] & b[8])^(a[266] & b[9])^(a[265] & b[10])^(a[264] & b[11])^(a[263] & b[12])^(a[262] & b[13])^(a[261] & b[14])^(a[260] & b[15])^(a[259] & b[16])^(a[258] & b[17])^(a[257] & b[18])^(a[256] & b[19])^(a[255] & b[20])^(a[254] & b[21])^(a[253] & b[22])^(a[252] & b[23])^(a[251] & b[24])^(a[250] & b[25])^(a[249] & b[26])^(a[248] & b[27])^(a[247] & b[28])^(a[246] & b[29])^(a[245] & b[30])^(a[244] & b[31])^(a[243] & b[32])^(a[242] & b[33])^(a[241] & b[34])^(a[240] & b[35])^(a[239] & b[36])^(a[238] & b[37])^(a[237] & b[38])^(a[236] & b[39])^(a[235] & b[40])^(a[234] & b[41])^(a[233] & b[42])^(a[232] & b[43])^(a[231] & b[44])^(a[230] & b[45])^(a[229] & b[46])^(a[228] & b[47])^(a[227] & b[48])^(a[226] & b[49])^(a[225] & b[50])^(a[224] & b[51])^(a[223] & b[52])^(a[222] & b[53])^(a[221] & b[54])^(a[220] & b[55])^(a[219] & b[56])^(a[218] & b[57])^(a[217] & b[58])^(a[216] & b[59])^(a[215] & b[60])^(a[214] & b[61])^(a[213] & b[62])^(a[212] & b[63])^(a[211] & b[64])^(a[210] & b[65])^(a[209] & b[66])^(a[208] & b[67])^(a[207] & b[68])^(a[206] & b[69])^(a[205] & b[70])^(a[204] & b[71])^(a[203] & b[72])^(a[202] & b[73])^(a[201] & b[74])^(a[200] & b[75])^(a[199] & b[76])^(a[198] & b[77])^(a[197] & b[78])^(a[196] & b[79])^(a[195] & b[80])^(a[194] & b[81])^(a[193] & b[82])^(a[192] & b[83])^(a[191] & b[84])^(a[190] & b[85])^(a[189] & b[86])^(a[188] & b[87])^(a[187] & b[88])^(a[186] & b[89])^(a[185] & b[90])^(a[184] & b[91])^(a[183] & b[92])^(a[182] & b[93])^(a[181] & b[94])^(a[180] & b[95])^(a[179] & b[96])^(a[178] & b[97])^(a[177] & b[98])^(a[176] & b[99])^(a[175] & b[100])^(a[174] & b[101])^(a[173] & b[102])^(a[172] & b[103])^(a[171] & b[104])^(a[170] & b[105])^(a[169] & b[106])^(a[168] & b[107])^(a[167] & b[108])^(a[166] & b[109])^(a[165] & b[110])^(a[164] & b[111])^(a[163] & b[112])^(a[162] & b[113])^(a[161] & b[114])^(a[160] & b[115])^(a[159] & b[116])^(a[158] & b[117])^(a[157] & b[118])^(a[156] & b[119])^(a[155] & b[120])^(a[154] & b[121])^(a[153] & b[122])^(a[152] & b[123])^(a[151] & b[124])^(a[150] & b[125])^(a[149] & b[126])^(a[148] & b[127])^(a[147] & b[128])^(a[146] & b[129])^(a[145] & b[130])^(a[144] & b[131])^(a[143] & b[132])^(a[142] & b[133])^(a[141] & b[134])^(a[140] & b[135])^(a[139] & b[136])^(a[138] & b[137])^(a[137] & b[138])^(a[136] & b[139])^(a[135] & b[140])^(a[134] & b[141])^(a[133] & b[142])^(a[132] & b[143])^(a[131] & b[144])^(a[130] & b[145])^(a[129] & b[146])^(a[128] & b[147])^(a[127] & b[148])^(a[126] & b[149])^(a[125] & b[150])^(a[124] & b[151])^(a[123] & b[152])^(a[122] & b[153])^(a[121] & b[154])^(a[120] & b[155])^(a[119] & b[156])^(a[118] & b[157])^(a[117] & b[158])^(a[116] & b[159])^(a[115] & b[160])^(a[114] & b[161])^(a[113] & b[162])^(a[112] & b[163])^(a[111] & b[164])^(a[110] & b[165])^(a[109] & b[166])^(a[108] & b[167])^(a[107] & b[168])^(a[106] & b[169])^(a[105] & b[170])^(a[104] & b[171])^(a[103] & b[172])^(a[102] & b[173])^(a[101] & b[174])^(a[100] & b[175])^(a[99] & b[176])^(a[98] & b[177])^(a[97] & b[178])^(a[96] & b[179])^(a[95] & b[180])^(a[94] & b[181])^(a[93] & b[182])^(a[92] & b[183])^(a[91] & b[184])^(a[90] & b[185])^(a[89] & b[186])^(a[88] & b[187])^(a[87] & b[188])^(a[86] & b[189])^(a[85] & b[190])^(a[84] & b[191])^(a[83] & b[192])^(a[82] & b[193])^(a[81] & b[194])^(a[80] & b[195])^(a[79] & b[196])^(a[78] & b[197])^(a[77] & b[198])^(a[76] & b[199])^(a[75] & b[200])^(a[74] & b[201])^(a[73] & b[202])^(a[72] & b[203])^(a[71] & b[204])^(a[70] & b[205])^(a[69] & b[206])^(a[68] & b[207])^(a[67] & b[208])^(a[66] & b[209])^(a[65] & b[210])^(a[64] & b[211])^(a[63] & b[212])^(a[62] & b[213])^(a[61] & b[214])^(a[60] & b[215])^(a[59] & b[216])^(a[58] & b[217])^(a[57] & b[218])^(a[56] & b[219])^(a[55] & b[220])^(a[54] & b[221])^(a[53] & b[222])^(a[52] & b[223])^(a[51] & b[224])^(a[50] & b[225])^(a[49] & b[226])^(a[48] & b[227])^(a[47] & b[228])^(a[46] & b[229])^(a[45] & b[230])^(a[44] & b[231])^(a[43] & b[232])^(a[42] & b[233])^(a[41] & b[234])^(a[40] & b[235])^(a[39] & b[236])^(a[38] & b[237])^(a[37] & b[238])^(a[36] & b[239])^(a[35] & b[240])^(a[34] & b[241])^(a[33] & b[242])^(a[32] & b[243])^(a[31] & b[244])^(a[30] & b[245])^(a[29] & b[246])^(a[28] & b[247])^(a[27] & b[248])^(a[26] & b[249])^(a[25] & b[250])^(a[24] & b[251])^(a[23] & b[252])^(a[22] & b[253])^(a[21] & b[254])^(a[20] & b[255])^(a[19] & b[256])^(a[18] & b[257])^(a[17] & b[258])^(a[16] & b[259])^(a[15] & b[260])^(a[14] & b[261])^(a[13] & b[262])^(a[12] & b[263])^(a[11] & b[264])^(a[10] & b[265])^(a[9] & b[266])^(a[8] & b[267])^(a[7] & b[268])^(a[6] & b[269])^(a[5] & b[270])^(a[4] & b[271])^(a[3] & b[272])^(a[2] & b[273])^(a[1] & b[274])^(a[0] & b[275]);
assign y[276] = (a[276] & b[0])^(a[275] & b[1])^(a[274] & b[2])^(a[273] & b[3])^(a[272] & b[4])^(a[271] & b[5])^(a[270] & b[6])^(a[269] & b[7])^(a[268] & b[8])^(a[267] & b[9])^(a[266] & b[10])^(a[265] & b[11])^(a[264] & b[12])^(a[263] & b[13])^(a[262] & b[14])^(a[261] & b[15])^(a[260] & b[16])^(a[259] & b[17])^(a[258] & b[18])^(a[257] & b[19])^(a[256] & b[20])^(a[255] & b[21])^(a[254] & b[22])^(a[253] & b[23])^(a[252] & b[24])^(a[251] & b[25])^(a[250] & b[26])^(a[249] & b[27])^(a[248] & b[28])^(a[247] & b[29])^(a[246] & b[30])^(a[245] & b[31])^(a[244] & b[32])^(a[243] & b[33])^(a[242] & b[34])^(a[241] & b[35])^(a[240] & b[36])^(a[239] & b[37])^(a[238] & b[38])^(a[237] & b[39])^(a[236] & b[40])^(a[235] & b[41])^(a[234] & b[42])^(a[233] & b[43])^(a[232] & b[44])^(a[231] & b[45])^(a[230] & b[46])^(a[229] & b[47])^(a[228] & b[48])^(a[227] & b[49])^(a[226] & b[50])^(a[225] & b[51])^(a[224] & b[52])^(a[223] & b[53])^(a[222] & b[54])^(a[221] & b[55])^(a[220] & b[56])^(a[219] & b[57])^(a[218] & b[58])^(a[217] & b[59])^(a[216] & b[60])^(a[215] & b[61])^(a[214] & b[62])^(a[213] & b[63])^(a[212] & b[64])^(a[211] & b[65])^(a[210] & b[66])^(a[209] & b[67])^(a[208] & b[68])^(a[207] & b[69])^(a[206] & b[70])^(a[205] & b[71])^(a[204] & b[72])^(a[203] & b[73])^(a[202] & b[74])^(a[201] & b[75])^(a[200] & b[76])^(a[199] & b[77])^(a[198] & b[78])^(a[197] & b[79])^(a[196] & b[80])^(a[195] & b[81])^(a[194] & b[82])^(a[193] & b[83])^(a[192] & b[84])^(a[191] & b[85])^(a[190] & b[86])^(a[189] & b[87])^(a[188] & b[88])^(a[187] & b[89])^(a[186] & b[90])^(a[185] & b[91])^(a[184] & b[92])^(a[183] & b[93])^(a[182] & b[94])^(a[181] & b[95])^(a[180] & b[96])^(a[179] & b[97])^(a[178] & b[98])^(a[177] & b[99])^(a[176] & b[100])^(a[175] & b[101])^(a[174] & b[102])^(a[173] & b[103])^(a[172] & b[104])^(a[171] & b[105])^(a[170] & b[106])^(a[169] & b[107])^(a[168] & b[108])^(a[167] & b[109])^(a[166] & b[110])^(a[165] & b[111])^(a[164] & b[112])^(a[163] & b[113])^(a[162] & b[114])^(a[161] & b[115])^(a[160] & b[116])^(a[159] & b[117])^(a[158] & b[118])^(a[157] & b[119])^(a[156] & b[120])^(a[155] & b[121])^(a[154] & b[122])^(a[153] & b[123])^(a[152] & b[124])^(a[151] & b[125])^(a[150] & b[126])^(a[149] & b[127])^(a[148] & b[128])^(a[147] & b[129])^(a[146] & b[130])^(a[145] & b[131])^(a[144] & b[132])^(a[143] & b[133])^(a[142] & b[134])^(a[141] & b[135])^(a[140] & b[136])^(a[139] & b[137])^(a[138] & b[138])^(a[137] & b[139])^(a[136] & b[140])^(a[135] & b[141])^(a[134] & b[142])^(a[133] & b[143])^(a[132] & b[144])^(a[131] & b[145])^(a[130] & b[146])^(a[129] & b[147])^(a[128] & b[148])^(a[127] & b[149])^(a[126] & b[150])^(a[125] & b[151])^(a[124] & b[152])^(a[123] & b[153])^(a[122] & b[154])^(a[121] & b[155])^(a[120] & b[156])^(a[119] & b[157])^(a[118] & b[158])^(a[117] & b[159])^(a[116] & b[160])^(a[115] & b[161])^(a[114] & b[162])^(a[113] & b[163])^(a[112] & b[164])^(a[111] & b[165])^(a[110] & b[166])^(a[109] & b[167])^(a[108] & b[168])^(a[107] & b[169])^(a[106] & b[170])^(a[105] & b[171])^(a[104] & b[172])^(a[103] & b[173])^(a[102] & b[174])^(a[101] & b[175])^(a[100] & b[176])^(a[99] & b[177])^(a[98] & b[178])^(a[97] & b[179])^(a[96] & b[180])^(a[95] & b[181])^(a[94] & b[182])^(a[93] & b[183])^(a[92] & b[184])^(a[91] & b[185])^(a[90] & b[186])^(a[89] & b[187])^(a[88] & b[188])^(a[87] & b[189])^(a[86] & b[190])^(a[85] & b[191])^(a[84] & b[192])^(a[83] & b[193])^(a[82] & b[194])^(a[81] & b[195])^(a[80] & b[196])^(a[79] & b[197])^(a[78] & b[198])^(a[77] & b[199])^(a[76] & b[200])^(a[75] & b[201])^(a[74] & b[202])^(a[73] & b[203])^(a[72] & b[204])^(a[71] & b[205])^(a[70] & b[206])^(a[69] & b[207])^(a[68] & b[208])^(a[67] & b[209])^(a[66] & b[210])^(a[65] & b[211])^(a[64] & b[212])^(a[63] & b[213])^(a[62] & b[214])^(a[61] & b[215])^(a[60] & b[216])^(a[59] & b[217])^(a[58] & b[218])^(a[57] & b[219])^(a[56] & b[220])^(a[55] & b[221])^(a[54] & b[222])^(a[53] & b[223])^(a[52] & b[224])^(a[51] & b[225])^(a[50] & b[226])^(a[49] & b[227])^(a[48] & b[228])^(a[47] & b[229])^(a[46] & b[230])^(a[45] & b[231])^(a[44] & b[232])^(a[43] & b[233])^(a[42] & b[234])^(a[41] & b[235])^(a[40] & b[236])^(a[39] & b[237])^(a[38] & b[238])^(a[37] & b[239])^(a[36] & b[240])^(a[35] & b[241])^(a[34] & b[242])^(a[33] & b[243])^(a[32] & b[244])^(a[31] & b[245])^(a[30] & b[246])^(a[29] & b[247])^(a[28] & b[248])^(a[27] & b[249])^(a[26] & b[250])^(a[25] & b[251])^(a[24] & b[252])^(a[23] & b[253])^(a[22] & b[254])^(a[21] & b[255])^(a[20] & b[256])^(a[19] & b[257])^(a[18] & b[258])^(a[17] & b[259])^(a[16] & b[260])^(a[15] & b[261])^(a[14] & b[262])^(a[13] & b[263])^(a[12] & b[264])^(a[11] & b[265])^(a[10] & b[266])^(a[9] & b[267])^(a[8] & b[268])^(a[7] & b[269])^(a[6] & b[270])^(a[5] & b[271])^(a[4] & b[272])^(a[3] & b[273])^(a[2] & b[274])^(a[1] & b[275])^(a[0] & b[276]);
assign y[277] = (a[277] & b[0])^(a[276] & b[1])^(a[275] & b[2])^(a[274] & b[3])^(a[273] & b[4])^(a[272] & b[5])^(a[271] & b[6])^(a[270] & b[7])^(a[269] & b[8])^(a[268] & b[9])^(a[267] & b[10])^(a[266] & b[11])^(a[265] & b[12])^(a[264] & b[13])^(a[263] & b[14])^(a[262] & b[15])^(a[261] & b[16])^(a[260] & b[17])^(a[259] & b[18])^(a[258] & b[19])^(a[257] & b[20])^(a[256] & b[21])^(a[255] & b[22])^(a[254] & b[23])^(a[253] & b[24])^(a[252] & b[25])^(a[251] & b[26])^(a[250] & b[27])^(a[249] & b[28])^(a[248] & b[29])^(a[247] & b[30])^(a[246] & b[31])^(a[245] & b[32])^(a[244] & b[33])^(a[243] & b[34])^(a[242] & b[35])^(a[241] & b[36])^(a[240] & b[37])^(a[239] & b[38])^(a[238] & b[39])^(a[237] & b[40])^(a[236] & b[41])^(a[235] & b[42])^(a[234] & b[43])^(a[233] & b[44])^(a[232] & b[45])^(a[231] & b[46])^(a[230] & b[47])^(a[229] & b[48])^(a[228] & b[49])^(a[227] & b[50])^(a[226] & b[51])^(a[225] & b[52])^(a[224] & b[53])^(a[223] & b[54])^(a[222] & b[55])^(a[221] & b[56])^(a[220] & b[57])^(a[219] & b[58])^(a[218] & b[59])^(a[217] & b[60])^(a[216] & b[61])^(a[215] & b[62])^(a[214] & b[63])^(a[213] & b[64])^(a[212] & b[65])^(a[211] & b[66])^(a[210] & b[67])^(a[209] & b[68])^(a[208] & b[69])^(a[207] & b[70])^(a[206] & b[71])^(a[205] & b[72])^(a[204] & b[73])^(a[203] & b[74])^(a[202] & b[75])^(a[201] & b[76])^(a[200] & b[77])^(a[199] & b[78])^(a[198] & b[79])^(a[197] & b[80])^(a[196] & b[81])^(a[195] & b[82])^(a[194] & b[83])^(a[193] & b[84])^(a[192] & b[85])^(a[191] & b[86])^(a[190] & b[87])^(a[189] & b[88])^(a[188] & b[89])^(a[187] & b[90])^(a[186] & b[91])^(a[185] & b[92])^(a[184] & b[93])^(a[183] & b[94])^(a[182] & b[95])^(a[181] & b[96])^(a[180] & b[97])^(a[179] & b[98])^(a[178] & b[99])^(a[177] & b[100])^(a[176] & b[101])^(a[175] & b[102])^(a[174] & b[103])^(a[173] & b[104])^(a[172] & b[105])^(a[171] & b[106])^(a[170] & b[107])^(a[169] & b[108])^(a[168] & b[109])^(a[167] & b[110])^(a[166] & b[111])^(a[165] & b[112])^(a[164] & b[113])^(a[163] & b[114])^(a[162] & b[115])^(a[161] & b[116])^(a[160] & b[117])^(a[159] & b[118])^(a[158] & b[119])^(a[157] & b[120])^(a[156] & b[121])^(a[155] & b[122])^(a[154] & b[123])^(a[153] & b[124])^(a[152] & b[125])^(a[151] & b[126])^(a[150] & b[127])^(a[149] & b[128])^(a[148] & b[129])^(a[147] & b[130])^(a[146] & b[131])^(a[145] & b[132])^(a[144] & b[133])^(a[143] & b[134])^(a[142] & b[135])^(a[141] & b[136])^(a[140] & b[137])^(a[139] & b[138])^(a[138] & b[139])^(a[137] & b[140])^(a[136] & b[141])^(a[135] & b[142])^(a[134] & b[143])^(a[133] & b[144])^(a[132] & b[145])^(a[131] & b[146])^(a[130] & b[147])^(a[129] & b[148])^(a[128] & b[149])^(a[127] & b[150])^(a[126] & b[151])^(a[125] & b[152])^(a[124] & b[153])^(a[123] & b[154])^(a[122] & b[155])^(a[121] & b[156])^(a[120] & b[157])^(a[119] & b[158])^(a[118] & b[159])^(a[117] & b[160])^(a[116] & b[161])^(a[115] & b[162])^(a[114] & b[163])^(a[113] & b[164])^(a[112] & b[165])^(a[111] & b[166])^(a[110] & b[167])^(a[109] & b[168])^(a[108] & b[169])^(a[107] & b[170])^(a[106] & b[171])^(a[105] & b[172])^(a[104] & b[173])^(a[103] & b[174])^(a[102] & b[175])^(a[101] & b[176])^(a[100] & b[177])^(a[99] & b[178])^(a[98] & b[179])^(a[97] & b[180])^(a[96] & b[181])^(a[95] & b[182])^(a[94] & b[183])^(a[93] & b[184])^(a[92] & b[185])^(a[91] & b[186])^(a[90] & b[187])^(a[89] & b[188])^(a[88] & b[189])^(a[87] & b[190])^(a[86] & b[191])^(a[85] & b[192])^(a[84] & b[193])^(a[83] & b[194])^(a[82] & b[195])^(a[81] & b[196])^(a[80] & b[197])^(a[79] & b[198])^(a[78] & b[199])^(a[77] & b[200])^(a[76] & b[201])^(a[75] & b[202])^(a[74] & b[203])^(a[73] & b[204])^(a[72] & b[205])^(a[71] & b[206])^(a[70] & b[207])^(a[69] & b[208])^(a[68] & b[209])^(a[67] & b[210])^(a[66] & b[211])^(a[65] & b[212])^(a[64] & b[213])^(a[63] & b[214])^(a[62] & b[215])^(a[61] & b[216])^(a[60] & b[217])^(a[59] & b[218])^(a[58] & b[219])^(a[57] & b[220])^(a[56] & b[221])^(a[55] & b[222])^(a[54] & b[223])^(a[53] & b[224])^(a[52] & b[225])^(a[51] & b[226])^(a[50] & b[227])^(a[49] & b[228])^(a[48] & b[229])^(a[47] & b[230])^(a[46] & b[231])^(a[45] & b[232])^(a[44] & b[233])^(a[43] & b[234])^(a[42] & b[235])^(a[41] & b[236])^(a[40] & b[237])^(a[39] & b[238])^(a[38] & b[239])^(a[37] & b[240])^(a[36] & b[241])^(a[35] & b[242])^(a[34] & b[243])^(a[33] & b[244])^(a[32] & b[245])^(a[31] & b[246])^(a[30] & b[247])^(a[29] & b[248])^(a[28] & b[249])^(a[27] & b[250])^(a[26] & b[251])^(a[25] & b[252])^(a[24] & b[253])^(a[23] & b[254])^(a[22] & b[255])^(a[21] & b[256])^(a[20] & b[257])^(a[19] & b[258])^(a[18] & b[259])^(a[17] & b[260])^(a[16] & b[261])^(a[15] & b[262])^(a[14] & b[263])^(a[13] & b[264])^(a[12] & b[265])^(a[11] & b[266])^(a[10] & b[267])^(a[9] & b[268])^(a[8] & b[269])^(a[7] & b[270])^(a[6] & b[271])^(a[5] & b[272])^(a[4] & b[273])^(a[3] & b[274])^(a[2] & b[275])^(a[1] & b[276])^(a[0] & b[277]);
assign y[278] = (a[278] & b[0])^(a[277] & b[1])^(a[276] & b[2])^(a[275] & b[3])^(a[274] & b[4])^(a[273] & b[5])^(a[272] & b[6])^(a[271] & b[7])^(a[270] & b[8])^(a[269] & b[9])^(a[268] & b[10])^(a[267] & b[11])^(a[266] & b[12])^(a[265] & b[13])^(a[264] & b[14])^(a[263] & b[15])^(a[262] & b[16])^(a[261] & b[17])^(a[260] & b[18])^(a[259] & b[19])^(a[258] & b[20])^(a[257] & b[21])^(a[256] & b[22])^(a[255] & b[23])^(a[254] & b[24])^(a[253] & b[25])^(a[252] & b[26])^(a[251] & b[27])^(a[250] & b[28])^(a[249] & b[29])^(a[248] & b[30])^(a[247] & b[31])^(a[246] & b[32])^(a[245] & b[33])^(a[244] & b[34])^(a[243] & b[35])^(a[242] & b[36])^(a[241] & b[37])^(a[240] & b[38])^(a[239] & b[39])^(a[238] & b[40])^(a[237] & b[41])^(a[236] & b[42])^(a[235] & b[43])^(a[234] & b[44])^(a[233] & b[45])^(a[232] & b[46])^(a[231] & b[47])^(a[230] & b[48])^(a[229] & b[49])^(a[228] & b[50])^(a[227] & b[51])^(a[226] & b[52])^(a[225] & b[53])^(a[224] & b[54])^(a[223] & b[55])^(a[222] & b[56])^(a[221] & b[57])^(a[220] & b[58])^(a[219] & b[59])^(a[218] & b[60])^(a[217] & b[61])^(a[216] & b[62])^(a[215] & b[63])^(a[214] & b[64])^(a[213] & b[65])^(a[212] & b[66])^(a[211] & b[67])^(a[210] & b[68])^(a[209] & b[69])^(a[208] & b[70])^(a[207] & b[71])^(a[206] & b[72])^(a[205] & b[73])^(a[204] & b[74])^(a[203] & b[75])^(a[202] & b[76])^(a[201] & b[77])^(a[200] & b[78])^(a[199] & b[79])^(a[198] & b[80])^(a[197] & b[81])^(a[196] & b[82])^(a[195] & b[83])^(a[194] & b[84])^(a[193] & b[85])^(a[192] & b[86])^(a[191] & b[87])^(a[190] & b[88])^(a[189] & b[89])^(a[188] & b[90])^(a[187] & b[91])^(a[186] & b[92])^(a[185] & b[93])^(a[184] & b[94])^(a[183] & b[95])^(a[182] & b[96])^(a[181] & b[97])^(a[180] & b[98])^(a[179] & b[99])^(a[178] & b[100])^(a[177] & b[101])^(a[176] & b[102])^(a[175] & b[103])^(a[174] & b[104])^(a[173] & b[105])^(a[172] & b[106])^(a[171] & b[107])^(a[170] & b[108])^(a[169] & b[109])^(a[168] & b[110])^(a[167] & b[111])^(a[166] & b[112])^(a[165] & b[113])^(a[164] & b[114])^(a[163] & b[115])^(a[162] & b[116])^(a[161] & b[117])^(a[160] & b[118])^(a[159] & b[119])^(a[158] & b[120])^(a[157] & b[121])^(a[156] & b[122])^(a[155] & b[123])^(a[154] & b[124])^(a[153] & b[125])^(a[152] & b[126])^(a[151] & b[127])^(a[150] & b[128])^(a[149] & b[129])^(a[148] & b[130])^(a[147] & b[131])^(a[146] & b[132])^(a[145] & b[133])^(a[144] & b[134])^(a[143] & b[135])^(a[142] & b[136])^(a[141] & b[137])^(a[140] & b[138])^(a[139] & b[139])^(a[138] & b[140])^(a[137] & b[141])^(a[136] & b[142])^(a[135] & b[143])^(a[134] & b[144])^(a[133] & b[145])^(a[132] & b[146])^(a[131] & b[147])^(a[130] & b[148])^(a[129] & b[149])^(a[128] & b[150])^(a[127] & b[151])^(a[126] & b[152])^(a[125] & b[153])^(a[124] & b[154])^(a[123] & b[155])^(a[122] & b[156])^(a[121] & b[157])^(a[120] & b[158])^(a[119] & b[159])^(a[118] & b[160])^(a[117] & b[161])^(a[116] & b[162])^(a[115] & b[163])^(a[114] & b[164])^(a[113] & b[165])^(a[112] & b[166])^(a[111] & b[167])^(a[110] & b[168])^(a[109] & b[169])^(a[108] & b[170])^(a[107] & b[171])^(a[106] & b[172])^(a[105] & b[173])^(a[104] & b[174])^(a[103] & b[175])^(a[102] & b[176])^(a[101] & b[177])^(a[100] & b[178])^(a[99] & b[179])^(a[98] & b[180])^(a[97] & b[181])^(a[96] & b[182])^(a[95] & b[183])^(a[94] & b[184])^(a[93] & b[185])^(a[92] & b[186])^(a[91] & b[187])^(a[90] & b[188])^(a[89] & b[189])^(a[88] & b[190])^(a[87] & b[191])^(a[86] & b[192])^(a[85] & b[193])^(a[84] & b[194])^(a[83] & b[195])^(a[82] & b[196])^(a[81] & b[197])^(a[80] & b[198])^(a[79] & b[199])^(a[78] & b[200])^(a[77] & b[201])^(a[76] & b[202])^(a[75] & b[203])^(a[74] & b[204])^(a[73] & b[205])^(a[72] & b[206])^(a[71] & b[207])^(a[70] & b[208])^(a[69] & b[209])^(a[68] & b[210])^(a[67] & b[211])^(a[66] & b[212])^(a[65] & b[213])^(a[64] & b[214])^(a[63] & b[215])^(a[62] & b[216])^(a[61] & b[217])^(a[60] & b[218])^(a[59] & b[219])^(a[58] & b[220])^(a[57] & b[221])^(a[56] & b[222])^(a[55] & b[223])^(a[54] & b[224])^(a[53] & b[225])^(a[52] & b[226])^(a[51] & b[227])^(a[50] & b[228])^(a[49] & b[229])^(a[48] & b[230])^(a[47] & b[231])^(a[46] & b[232])^(a[45] & b[233])^(a[44] & b[234])^(a[43] & b[235])^(a[42] & b[236])^(a[41] & b[237])^(a[40] & b[238])^(a[39] & b[239])^(a[38] & b[240])^(a[37] & b[241])^(a[36] & b[242])^(a[35] & b[243])^(a[34] & b[244])^(a[33] & b[245])^(a[32] & b[246])^(a[31] & b[247])^(a[30] & b[248])^(a[29] & b[249])^(a[28] & b[250])^(a[27] & b[251])^(a[26] & b[252])^(a[25] & b[253])^(a[24] & b[254])^(a[23] & b[255])^(a[22] & b[256])^(a[21] & b[257])^(a[20] & b[258])^(a[19] & b[259])^(a[18] & b[260])^(a[17] & b[261])^(a[16] & b[262])^(a[15] & b[263])^(a[14] & b[264])^(a[13] & b[265])^(a[12] & b[266])^(a[11] & b[267])^(a[10] & b[268])^(a[9] & b[269])^(a[8] & b[270])^(a[7] & b[271])^(a[6] & b[272])^(a[5] & b[273])^(a[4] & b[274])^(a[3] & b[275])^(a[2] & b[276])^(a[1] & b[277])^(a[0] & b[278]);
assign y[279] = (a[279] & b[0])^(a[278] & b[1])^(a[277] & b[2])^(a[276] & b[3])^(a[275] & b[4])^(a[274] & b[5])^(a[273] & b[6])^(a[272] & b[7])^(a[271] & b[8])^(a[270] & b[9])^(a[269] & b[10])^(a[268] & b[11])^(a[267] & b[12])^(a[266] & b[13])^(a[265] & b[14])^(a[264] & b[15])^(a[263] & b[16])^(a[262] & b[17])^(a[261] & b[18])^(a[260] & b[19])^(a[259] & b[20])^(a[258] & b[21])^(a[257] & b[22])^(a[256] & b[23])^(a[255] & b[24])^(a[254] & b[25])^(a[253] & b[26])^(a[252] & b[27])^(a[251] & b[28])^(a[250] & b[29])^(a[249] & b[30])^(a[248] & b[31])^(a[247] & b[32])^(a[246] & b[33])^(a[245] & b[34])^(a[244] & b[35])^(a[243] & b[36])^(a[242] & b[37])^(a[241] & b[38])^(a[240] & b[39])^(a[239] & b[40])^(a[238] & b[41])^(a[237] & b[42])^(a[236] & b[43])^(a[235] & b[44])^(a[234] & b[45])^(a[233] & b[46])^(a[232] & b[47])^(a[231] & b[48])^(a[230] & b[49])^(a[229] & b[50])^(a[228] & b[51])^(a[227] & b[52])^(a[226] & b[53])^(a[225] & b[54])^(a[224] & b[55])^(a[223] & b[56])^(a[222] & b[57])^(a[221] & b[58])^(a[220] & b[59])^(a[219] & b[60])^(a[218] & b[61])^(a[217] & b[62])^(a[216] & b[63])^(a[215] & b[64])^(a[214] & b[65])^(a[213] & b[66])^(a[212] & b[67])^(a[211] & b[68])^(a[210] & b[69])^(a[209] & b[70])^(a[208] & b[71])^(a[207] & b[72])^(a[206] & b[73])^(a[205] & b[74])^(a[204] & b[75])^(a[203] & b[76])^(a[202] & b[77])^(a[201] & b[78])^(a[200] & b[79])^(a[199] & b[80])^(a[198] & b[81])^(a[197] & b[82])^(a[196] & b[83])^(a[195] & b[84])^(a[194] & b[85])^(a[193] & b[86])^(a[192] & b[87])^(a[191] & b[88])^(a[190] & b[89])^(a[189] & b[90])^(a[188] & b[91])^(a[187] & b[92])^(a[186] & b[93])^(a[185] & b[94])^(a[184] & b[95])^(a[183] & b[96])^(a[182] & b[97])^(a[181] & b[98])^(a[180] & b[99])^(a[179] & b[100])^(a[178] & b[101])^(a[177] & b[102])^(a[176] & b[103])^(a[175] & b[104])^(a[174] & b[105])^(a[173] & b[106])^(a[172] & b[107])^(a[171] & b[108])^(a[170] & b[109])^(a[169] & b[110])^(a[168] & b[111])^(a[167] & b[112])^(a[166] & b[113])^(a[165] & b[114])^(a[164] & b[115])^(a[163] & b[116])^(a[162] & b[117])^(a[161] & b[118])^(a[160] & b[119])^(a[159] & b[120])^(a[158] & b[121])^(a[157] & b[122])^(a[156] & b[123])^(a[155] & b[124])^(a[154] & b[125])^(a[153] & b[126])^(a[152] & b[127])^(a[151] & b[128])^(a[150] & b[129])^(a[149] & b[130])^(a[148] & b[131])^(a[147] & b[132])^(a[146] & b[133])^(a[145] & b[134])^(a[144] & b[135])^(a[143] & b[136])^(a[142] & b[137])^(a[141] & b[138])^(a[140] & b[139])^(a[139] & b[140])^(a[138] & b[141])^(a[137] & b[142])^(a[136] & b[143])^(a[135] & b[144])^(a[134] & b[145])^(a[133] & b[146])^(a[132] & b[147])^(a[131] & b[148])^(a[130] & b[149])^(a[129] & b[150])^(a[128] & b[151])^(a[127] & b[152])^(a[126] & b[153])^(a[125] & b[154])^(a[124] & b[155])^(a[123] & b[156])^(a[122] & b[157])^(a[121] & b[158])^(a[120] & b[159])^(a[119] & b[160])^(a[118] & b[161])^(a[117] & b[162])^(a[116] & b[163])^(a[115] & b[164])^(a[114] & b[165])^(a[113] & b[166])^(a[112] & b[167])^(a[111] & b[168])^(a[110] & b[169])^(a[109] & b[170])^(a[108] & b[171])^(a[107] & b[172])^(a[106] & b[173])^(a[105] & b[174])^(a[104] & b[175])^(a[103] & b[176])^(a[102] & b[177])^(a[101] & b[178])^(a[100] & b[179])^(a[99] & b[180])^(a[98] & b[181])^(a[97] & b[182])^(a[96] & b[183])^(a[95] & b[184])^(a[94] & b[185])^(a[93] & b[186])^(a[92] & b[187])^(a[91] & b[188])^(a[90] & b[189])^(a[89] & b[190])^(a[88] & b[191])^(a[87] & b[192])^(a[86] & b[193])^(a[85] & b[194])^(a[84] & b[195])^(a[83] & b[196])^(a[82] & b[197])^(a[81] & b[198])^(a[80] & b[199])^(a[79] & b[200])^(a[78] & b[201])^(a[77] & b[202])^(a[76] & b[203])^(a[75] & b[204])^(a[74] & b[205])^(a[73] & b[206])^(a[72] & b[207])^(a[71] & b[208])^(a[70] & b[209])^(a[69] & b[210])^(a[68] & b[211])^(a[67] & b[212])^(a[66] & b[213])^(a[65] & b[214])^(a[64] & b[215])^(a[63] & b[216])^(a[62] & b[217])^(a[61] & b[218])^(a[60] & b[219])^(a[59] & b[220])^(a[58] & b[221])^(a[57] & b[222])^(a[56] & b[223])^(a[55] & b[224])^(a[54] & b[225])^(a[53] & b[226])^(a[52] & b[227])^(a[51] & b[228])^(a[50] & b[229])^(a[49] & b[230])^(a[48] & b[231])^(a[47] & b[232])^(a[46] & b[233])^(a[45] & b[234])^(a[44] & b[235])^(a[43] & b[236])^(a[42] & b[237])^(a[41] & b[238])^(a[40] & b[239])^(a[39] & b[240])^(a[38] & b[241])^(a[37] & b[242])^(a[36] & b[243])^(a[35] & b[244])^(a[34] & b[245])^(a[33] & b[246])^(a[32] & b[247])^(a[31] & b[248])^(a[30] & b[249])^(a[29] & b[250])^(a[28] & b[251])^(a[27] & b[252])^(a[26] & b[253])^(a[25] & b[254])^(a[24] & b[255])^(a[23] & b[256])^(a[22] & b[257])^(a[21] & b[258])^(a[20] & b[259])^(a[19] & b[260])^(a[18] & b[261])^(a[17] & b[262])^(a[16] & b[263])^(a[15] & b[264])^(a[14] & b[265])^(a[13] & b[266])^(a[12] & b[267])^(a[11] & b[268])^(a[10] & b[269])^(a[9] & b[270])^(a[8] & b[271])^(a[7] & b[272])^(a[6] & b[273])^(a[5] & b[274])^(a[4] & b[275])^(a[3] & b[276])^(a[2] & b[277])^(a[1] & b[278])^(a[0] & b[279]);
assign y[280] = (a[280] & b[0])^(a[279] & b[1])^(a[278] & b[2])^(a[277] & b[3])^(a[276] & b[4])^(a[275] & b[5])^(a[274] & b[6])^(a[273] & b[7])^(a[272] & b[8])^(a[271] & b[9])^(a[270] & b[10])^(a[269] & b[11])^(a[268] & b[12])^(a[267] & b[13])^(a[266] & b[14])^(a[265] & b[15])^(a[264] & b[16])^(a[263] & b[17])^(a[262] & b[18])^(a[261] & b[19])^(a[260] & b[20])^(a[259] & b[21])^(a[258] & b[22])^(a[257] & b[23])^(a[256] & b[24])^(a[255] & b[25])^(a[254] & b[26])^(a[253] & b[27])^(a[252] & b[28])^(a[251] & b[29])^(a[250] & b[30])^(a[249] & b[31])^(a[248] & b[32])^(a[247] & b[33])^(a[246] & b[34])^(a[245] & b[35])^(a[244] & b[36])^(a[243] & b[37])^(a[242] & b[38])^(a[241] & b[39])^(a[240] & b[40])^(a[239] & b[41])^(a[238] & b[42])^(a[237] & b[43])^(a[236] & b[44])^(a[235] & b[45])^(a[234] & b[46])^(a[233] & b[47])^(a[232] & b[48])^(a[231] & b[49])^(a[230] & b[50])^(a[229] & b[51])^(a[228] & b[52])^(a[227] & b[53])^(a[226] & b[54])^(a[225] & b[55])^(a[224] & b[56])^(a[223] & b[57])^(a[222] & b[58])^(a[221] & b[59])^(a[220] & b[60])^(a[219] & b[61])^(a[218] & b[62])^(a[217] & b[63])^(a[216] & b[64])^(a[215] & b[65])^(a[214] & b[66])^(a[213] & b[67])^(a[212] & b[68])^(a[211] & b[69])^(a[210] & b[70])^(a[209] & b[71])^(a[208] & b[72])^(a[207] & b[73])^(a[206] & b[74])^(a[205] & b[75])^(a[204] & b[76])^(a[203] & b[77])^(a[202] & b[78])^(a[201] & b[79])^(a[200] & b[80])^(a[199] & b[81])^(a[198] & b[82])^(a[197] & b[83])^(a[196] & b[84])^(a[195] & b[85])^(a[194] & b[86])^(a[193] & b[87])^(a[192] & b[88])^(a[191] & b[89])^(a[190] & b[90])^(a[189] & b[91])^(a[188] & b[92])^(a[187] & b[93])^(a[186] & b[94])^(a[185] & b[95])^(a[184] & b[96])^(a[183] & b[97])^(a[182] & b[98])^(a[181] & b[99])^(a[180] & b[100])^(a[179] & b[101])^(a[178] & b[102])^(a[177] & b[103])^(a[176] & b[104])^(a[175] & b[105])^(a[174] & b[106])^(a[173] & b[107])^(a[172] & b[108])^(a[171] & b[109])^(a[170] & b[110])^(a[169] & b[111])^(a[168] & b[112])^(a[167] & b[113])^(a[166] & b[114])^(a[165] & b[115])^(a[164] & b[116])^(a[163] & b[117])^(a[162] & b[118])^(a[161] & b[119])^(a[160] & b[120])^(a[159] & b[121])^(a[158] & b[122])^(a[157] & b[123])^(a[156] & b[124])^(a[155] & b[125])^(a[154] & b[126])^(a[153] & b[127])^(a[152] & b[128])^(a[151] & b[129])^(a[150] & b[130])^(a[149] & b[131])^(a[148] & b[132])^(a[147] & b[133])^(a[146] & b[134])^(a[145] & b[135])^(a[144] & b[136])^(a[143] & b[137])^(a[142] & b[138])^(a[141] & b[139])^(a[140] & b[140])^(a[139] & b[141])^(a[138] & b[142])^(a[137] & b[143])^(a[136] & b[144])^(a[135] & b[145])^(a[134] & b[146])^(a[133] & b[147])^(a[132] & b[148])^(a[131] & b[149])^(a[130] & b[150])^(a[129] & b[151])^(a[128] & b[152])^(a[127] & b[153])^(a[126] & b[154])^(a[125] & b[155])^(a[124] & b[156])^(a[123] & b[157])^(a[122] & b[158])^(a[121] & b[159])^(a[120] & b[160])^(a[119] & b[161])^(a[118] & b[162])^(a[117] & b[163])^(a[116] & b[164])^(a[115] & b[165])^(a[114] & b[166])^(a[113] & b[167])^(a[112] & b[168])^(a[111] & b[169])^(a[110] & b[170])^(a[109] & b[171])^(a[108] & b[172])^(a[107] & b[173])^(a[106] & b[174])^(a[105] & b[175])^(a[104] & b[176])^(a[103] & b[177])^(a[102] & b[178])^(a[101] & b[179])^(a[100] & b[180])^(a[99] & b[181])^(a[98] & b[182])^(a[97] & b[183])^(a[96] & b[184])^(a[95] & b[185])^(a[94] & b[186])^(a[93] & b[187])^(a[92] & b[188])^(a[91] & b[189])^(a[90] & b[190])^(a[89] & b[191])^(a[88] & b[192])^(a[87] & b[193])^(a[86] & b[194])^(a[85] & b[195])^(a[84] & b[196])^(a[83] & b[197])^(a[82] & b[198])^(a[81] & b[199])^(a[80] & b[200])^(a[79] & b[201])^(a[78] & b[202])^(a[77] & b[203])^(a[76] & b[204])^(a[75] & b[205])^(a[74] & b[206])^(a[73] & b[207])^(a[72] & b[208])^(a[71] & b[209])^(a[70] & b[210])^(a[69] & b[211])^(a[68] & b[212])^(a[67] & b[213])^(a[66] & b[214])^(a[65] & b[215])^(a[64] & b[216])^(a[63] & b[217])^(a[62] & b[218])^(a[61] & b[219])^(a[60] & b[220])^(a[59] & b[221])^(a[58] & b[222])^(a[57] & b[223])^(a[56] & b[224])^(a[55] & b[225])^(a[54] & b[226])^(a[53] & b[227])^(a[52] & b[228])^(a[51] & b[229])^(a[50] & b[230])^(a[49] & b[231])^(a[48] & b[232])^(a[47] & b[233])^(a[46] & b[234])^(a[45] & b[235])^(a[44] & b[236])^(a[43] & b[237])^(a[42] & b[238])^(a[41] & b[239])^(a[40] & b[240])^(a[39] & b[241])^(a[38] & b[242])^(a[37] & b[243])^(a[36] & b[244])^(a[35] & b[245])^(a[34] & b[246])^(a[33] & b[247])^(a[32] & b[248])^(a[31] & b[249])^(a[30] & b[250])^(a[29] & b[251])^(a[28] & b[252])^(a[27] & b[253])^(a[26] & b[254])^(a[25] & b[255])^(a[24] & b[256])^(a[23] & b[257])^(a[22] & b[258])^(a[21] & b[259])^(a[20] & b[260])^(a[19] & b[261])^(a[18] & b[262])^(a[17] & b[263])^(a[16] & b[264])^(a[15] & b[265])^(a[14] & b[266])^(a[13] & b[267])^(a[12] & b[268])^(a[11] & b[269])^(a[10] & b[270])^(a[9] & b[271])^(a[8] & b[272])^(a[7] & b[273])^(a[6] & b[274])^(a[5] & b[275])^(a[4] & b[276])^(a[3] & b[277])^(a[2] & b[278])^(a[1] & b[279])^(a[0] & b[280]);
assign y[281] = (a[281] & b[0])^(a[280] & b[1])^(a[279] & b[2])^(a[278] & b[3])^(a[277] & b[4])^(a[276] & b[5])^(a[275] & b[6])^(a[274] & b[7])^(a[273] & b[8])^(a[272] & b[9])^(a[271] & b[10])^(a[270] & b[11])^(a[269] & b[12])^(a[268] & b[13])^(a[267] & b[14])^(a[266] & b[15])^(a[265] & b[16])^(a[264] & b[17])^(a[263] & b[18])^(a[262] & b[19])^(a[261] & b[20])^(a[260] & b[21])^(a[259] & b[22])^(a[258] & b[23])^(a[257] & b[24])^(a[256] & b[25])^(a[255] & b[26])^(a[254] & b[27])^(a[253] & b[28])^(a[252] & b[29])^(a[251] & b[30])^(a[250] & b[31])^(a[249] & b[32])^(a[248] & b[33])^(a[247] & b[34])^(a[246] & b[35])^(a[245] & b[36])^(a[244] & b[37])^(a[243] & b[38])^(a[242] & b[39])^(a[241] & b[40])^(a[240] & b[41])^(a[239] & b[42])^(a[238] & b[43])^(a[237] & b[44])^(a[236] & b[45])^(a[235] & b[46])^(a[234] & b[47])^(a[233] & b[48])^(a[232] & b[49])^(a[231] & b[50])^(a[230] & b[51])^(a[229] & b[52])^(a[228] & b[53])^(a[227] & b[54])^(a[226] & b[55])^(a[225] & b[56])^(a[224] & b[57])^(a[223] & b[58])^(a[222] & b[59])^(a[221] & b[60])^(a[220] & b[61])^(a[219] & b[62])^(a[218] & b[63])^(a[217] & b[64])^(a[216] & b[65])^(a[215] & b[66])^(a[214] & b[67])^(a[213] & b[68])^(a[212] & b[69])^(a[211] & b[70])^(a[210] & b[71])^(a[209] & b[72])^(a[208] & b[73])^(a[207] & b[74])^(a[206] & b[75])^(a[205] & b[76])^(a[204] & b[77])^(a[203] & b[78])^(a[202] & b[79])^(a[201] & b[80])^(a[200] & b[81])^(a[199] & b[82])^(a[198] & b[83])^(a[197] & b[84])^(a[196] & b[85])^(a[195] & b[86])^(a[194] & b[87])^(a[193] & b[88])^(a[192] & b[89])^(a[191] & b[90])^(a[190] & b[91])^(a[189] & b[92])^(a[188] & b[93])^(a[187] & b[94])^(a[186] & b[95])^(a[185] & b[96])^(a[184] & b[97])^(a[183] & b[98])^(a[182] & b[99])^(a[181] & b[100])^(a[180] & b[101])^(a[179] & b[102])^(a[178] & b[103])^(a[177] & b[104])^(a[176] & b[105])^(a[175] & b[106])^(a[174] & b[107])^(a[173] & b[108])^(a[172] & b[109])^(a[171] & b[110])^(a[170] & b[111])^(a[169] & b[112])^(a[168] & b[113])^(a[167] & b[114])^(a[166] & b[115])^(a[165] & b[116])^(a[164] & b[117])^(a[163] & b[118])^(a[162] & b[119])^(a[161] & b[120])^(a[160] & b[121])^(a[159] & b[122])^(a[158] & b[123])^(a[157] & b[124])^(a[156] & b[125])^(a[155] & b[126])^(a[154] & b[127])^(a[153] & b[128])^(a[152] & b[129])^(a[151] & b[130])^(a[150] & b[131])^(a[149] & b[132])^(a[148] & b[133])^(a[147] & b[134])^(a[146] & b[135])^(a[145] & b[136])^(a[144] & b[137])^(a[143] & b[138])^(a[142] & b[139])^(a[141] & b[140])^(a[140] & b[141])^(a[139] & b[142])^(a[138] & b[143])^(a[137] & b[144])^(a[136] & b[145])^(a[135] & b[146])^(a[134] & b[147])^(a[133] & b[148])^(a[132] & b[149])^(a[131] & b[150])^(a[130] & b[151])^(a[129] & b[152])^(a[128] & b[153])^(a[127] & b[154])^(a[126] & b[155])^(a[125] & b[156])^(a[124] & b[157])^(a[123] & b[158])^(a[122] & b[159])^(a[121] & b[160])^(a[120] & b[161])^(a[119] & b[162])^(a[118] & b[163])^(a[117] & b[164])^(a[116] & b[165])^(a[115] & b[166])^(a[114] & b[167])^(a[113] & b[168])^(a[112] & b[169])^(a[111] & b[170])^(a[110] & b[171])^(a[109] & b[172])^(a[108] & b[173])^(a[107] & b[174])^(a[106] & b[175])^(a[105] & b[176])^(a[104] & b[177])^(a[103] & b[178])^(a[102] & b[179])^(a[101] & b[180])^(a[100] & b[181])^(a[99] & b[182])^(a[98] & b[183])^(a[97] & b[184])^(a[96] & b[185])^(a[95] & b[186])^(a[94] & b[187])^(a[93] & b[188])^(a[92] & b[189])^(a[91] & b[190])^(a[90] & b[191])^(a[89] & b[192])^(a[88] & b[193])^(a[87] & b[194])^(a[86] & b[195])^(a[85] & b[196])^(a[84] & b[197])^(a[83] & b[198])^(a[82] & b[199])^(a[81] & b[200])^(a[80] & b[201])^(a[79] & b[202])^(a[78] & b[203])^(a[77] & b[204])^(a[76] & b[205])^(a[75] & b[206])^(a[74] & b[207])^(a[73] & b[208])^(a[72] & b[209])^(a[71] & b[210])^(a[70] & b[211])^(a[69] & b[212])^(a[68] & b[213])^(a[67] & b[214])^(a[66] & b[215])^(a[65] & b[216])^(a[64] & b[217])^(a[63] & b[218])^(a[62] & b[219])^(a[61] & b[220])^(a[60] & b[221])^(a[59] & b[222])^(a[58] & b[223])^(a[57] & b[224])^(a[56] & b[225])^(a[55] & b[226])^(a[54] & b[227])^(a[53] & b[228])^(a[52] & b[229])^(a[51] & b[230])^(a[50] & b[231])^(a[49] & b[232])^(a[48] & b[233])^(a[47] & b[234])^(a[46] & b[235])^(a[45] & b[236])^(a[44] & b[237])^(a[43] & b[238])^(a[42] & b[239])^(a[41] & b[240])^(a[40] & b[241])^(a[39] & b[242])^(a[38] & b[243])^(a[37] & b[244])^(a[36] & b[245])^(a[35] & b[246])^(a[34] & b[247])^(a[33] & b[248])^(a[32] & b[249])^(a[31] & b[250])^(a[30] & b[251])^(a[29] & b[252])^(a[28] & b[253])^(a[27] & b[254])^(a[26] & b[255])^(a[25] & b[256])^(a[24] & b[257])^(a[23] & b[258])^(a[22] & b[259])^(a[21] & b[260])^(a[20] & b[261])^(a[19] & b[262])^(a[18] & b[263])^(a[17] & b[264])^(a[16] & b[265])^(a[15] & b[266])^(a[14] & b[267])^(a[13] & b[268])^(a[12] & b[269])^(a[11] & b[270])^(a[10] & b[271])^(a[9] & b[272])^(a[8] & b[273])^(a[7] & b[274])^(a[6] & b[275])^(a[5] & b[276])^(a[4] & b[277])^(a[3] & b[278])^(a[2] & b[279])^(a[1] & b[280])^(a[0] & b[281]);
assign y[282] = (a[282] & b[0])^(a[281] & b[1])^(a[280] & b[2])^(a[279] & b[3])^(a[278] & b[4])^(a[277] & b[5])^(a[276] & b[6])^(a[275] & b[7])^(a[274] & b[8])^(a[273] & b[9])^(a[272] & b[10])^(a[271] & b[11])^(a[270] & b[12])^(a[269] & b[13])^(a[268] & b[14])^(a[267] & b[15])^(a[266] & b[16])^(a[265] & b[17])^(a[264] & b[18])^(a[263] & b[19])^(a[262] & b[20])^(a[261] & b[21])^(a[260] & b[22])^(a[259] & b[23])^(a[258] & b[24])^(a[257] & b[25])^(a[256] & b[26])^(a[255] & b[27])^(a[254] & b[28])^(a[253] & b[29])^(a[252] & b[30])^(a[251] & b[31])^(a[250] & b[32])^(a[249] & b[33])^(a[248] & b[34])^(a[247] & b[35])^(a[246] & b[36])^(a[245] & b[37])^(a[244] & b[38])^(a[243] & b[39])^(a[242] & b[40])^(a[241] & b[41])^(a[240] & b[42])^(a[239] & b[43])^(a[238] & b[44])^(a[237] & b[45])^(a[236] & b[46])^(a[235] & b[47])^(a[234] & b[48])^(a[233] & b[49])^(a[232] & b[50])^(a[231] & b[51])^(a[230] & b[52])^(a[229] & b[53])^(a[228] & b[54])^(a[227] & b[55])^(a[226] & b[56])^(a[225] & b[57])^(a[224] & b[58])^(a[223] & b[59])^(a[222] & b[60])^(a[221] & b[61])^(a[220] & b[62])^(a[219] & b[63])^(a[218] & b[64])^(a[217] & b[65])^(a[216] & b[66])^(a[215] & b[67])^(a[214] & b[68])^(a[213] & b[69])^(a[212] & b[70])^(a[211] & b[71])^(a[210] & b[72])^(a[209] & b[73])^(a[208] & b[74])^(a[207] & b[75])^(a[206] & b[76])^(a[205] & b[77])^(a[204] & b[78])^(a[203] & b[79])^(a[202] & b[80])^(a[201] & b[81])^(a[200] & b[82])^(a[199] & b[83])^(a[198] & b[84])^(a[197] & b[85])^(a[196] & b[86])^(a[195] & b[87])^(a[194] & b[88])^(a[193] & b[89])^(a[192] & b[90])^(a[191] & b[91])^(a[190] & b[92])^(a[189] & b[93])^(a[188] & b[94])^(a[187] & b[95])^(a[186] & b[96])^(a[185] & b[97])^(a[184] & b[98])^(a[183] & b[99])^(a[182] & b[100])^(a[181] & b[101])^(a[180] & b[102])^(a[179] & b[103])^(a[178] & b[104])^(a[177] & b[105])^(a[176] & b[106])^(a[175] & b[107])^(a[174] & b[108])^(a[173] & b[109])^(a[172] & b[110])^(a[171] & b[111])^(a[170] & b[112])^(a[169] & b[113])^(a[168] & b[114])^(a[167] & b[115])^(a[166] & b[116])^(a[165] & b[117])^(a[164] & b[118])^(a[163] & b[119])^(a[162] & b[120])^(a[161] & b[121])^(a[160] & b[122])^(a[159] & b[123])^(a[158] & b[124])^(a[157] & b[125])^(a[156] & b[126])^(a[155] & b[127])^(a[154] & b[128])^(a[153] & b[129])^(a[152] & b[130])^(a[151] & b[131])^(a[150] & b[132])^(a[149] & b[133])^(a[148] & b[134])^(a[147] & b[135])^(a[146] & b[136])^(a[145] & b[137])^(a[144] & b[138])^(a[143] & b[139])^(a[142] & b[140])^(a[141] & b[141])^(a[140] & b[142])^(a[139] & b[143])^(a[138] & b[144])^(a[137] & b[145])^(a[136] & b[146])^(a[135] & b[147])^(a[134] & b[148])^(a[133] & b[149])^(a[132] & b[150])^(a[131] & b[151])^(a[130] & b[152])^(a[129] & b[153])^(a[128] & b[154])^(a[127] & b[155])^(a[126] & b[156])^(a[125] & b[157])^(a[124] & b[158])^(a[123] & b[159])^(a[122] & b[160])^(a[121] & b[161])^(a[120] & b[162])^(a[119] & b[163])^(a[118] & b[164])^(a[117] & b[165])^(a[116] & b[166])^(a[115] & b[167])^(a[114] & b[168])^(a[113] & b[169])^(a[112] & b[170])^(a[111] & b[171])^(a[110] & b[172])^(a[109] & b[173])^(a[108] & b[174])^(a[107] & b[175])^(a[106] & b[176])^(a[105] & b[177])^(a[104] & b[178])^(a[103] & b[179])^(a[102] & b[180])^(a[101] & b[181])^(a[100] & b[182])^(a[99] & b[183])^(a[98] & b[184])^(a[97] & b[185])^(a[96] & b[186])^(a[95] & b[187])^(a[94] & b[188])^(a[93] & b[189])^(a[92] & b[190])^(a[91] & b[191])^(a[90] & b[192])^(a[89] & b[193])^(a[88] & b[194])^(a[87] & b[195])^(a[86] & b[196])^(a[85] & b[197])^(a[84] & b[198])^(a[83] & b[199])^(a[82] & b[200])^(a[81] & b[201])^(a[80] & b[202])^(a[79] & b[203])^(a[78] & b[204])^(a[77] & b[205])^(a[76] & b[206])^(a[75] & b[207])^(a[74] & b[208])^(a[73] & b[209])^(a[72] & b[210])^(a[71] & b[211])^(a[70] & b[212])^(a[69] & b[213])^(a[68] & b[214])^(a[67] & b[215])^(a[66] & b[216])^(a[65] & b[217])^(a[64] & b[218])^(a[63] & b[219])^(a[62] & b[220])^(a[61] & b[221])^(a[60] & b[222])^(a[59] & b[223])^(a[58] & b[224])^(a[57] & b[225])^(a[56] & b[226])^(a[55] & b[227])^(a[54] & b[228])^(a[53] & b[229])^(a[52] & b[230])^(a[51] & b[231])^(a[50] & b[232])^(a[49] & b[233])^(a[48] & b[234])^(a[47] & b[235])^(a[46] & b[236])^(a[45] & b[237])^(a[44] & b[238])^(a[43] & b[239])^(a[42] & b[240])^(a[41] & b[241])^(a[40] & b[242])^(a[39] & b[243])^(a[38] & b[244])^(a[37] & b[245])^(a[36] & b[246])^(a[35] & b[247])^(a[34] & b[248])^(a[33] & b[249])^(a[32] & b[250])^(a[31] & b[251])^(a[30] & b[252])^(a[29] & b[253])^(a[28] & b[254])^(a[27] & b[255])^(a[26] & b[256])^(a[25] & b[257])^(a[24] & b[258])^(a[23] & b[259])^(a[22] & b[260])^(a[21] & b[261])^(a[20] & b[262])^(a[19] & b[263])^(a[18] & b[264])^(a[17] & b[265])^(a[16] & b[266])^(a[15] & b[267])^(a[14] & b[268])^(a[13] & b[269])^(a[12] & b[270])^(a[11] & b[271])^(a[10] & b[272])^(a[9] & b[273])^(a[8] & b[274])^(a[7] & b[275])^(a[6] & b[276])^(a[5] & b[277])^(a[4] & b[278])^(a[3] & b[279])^(a[2] & b[280])^(a[1] & b[281])^(a[0] & b[282]);
assign y[283] = (a[283] & b[0])^(a[282] & b[1])^(a[281] & b[2])^(a[280] & b[3])^(a[279] & b[4])^(a[278] & b[5])^(a[277] & b[6])^(a[276] & b[7])^(a[275] & b[8])^(a[274] & b[9])^(a[273] & b[10])^(a[272] & b[11])^(a[271] & b[12])^(a[270] & b[13])^(a[269] & b[14])^(a[268] & b[15])^(a[267] & b[16])^(a[266] & b[17])^(a[265] & b[18])^(a[264] & b[19])^(a[263] & b[20])^(a[262] & b[21])^(a[261] & b[22])^(a[260] & b[23])^(a[259] & b[24])^(a[258] & b[25])^(a[257] & b[26])^(a[256] & b[27])^(a[255] & b[28])^(a[254] & b[29])^(a[253] & b[30])^(a[252] & b[31])^(a[251] & b[32])^(a[250] & b[33])^(a[249] & b[34])^(a[248] & b[35])^(a[247] & b[36])^(a[246] & b[37])^(a[245] & b[38])^(a[244] & b[39])^(a[243] & b[40])^(a[242] & b[41])^(a[241] & b[42])^(a[240] & b[43])^(a[239] & b[44])^(a[238] & b[45])^(a[237] & b[46])^(a[236] & b[47])^(a[235] & b[48])^(a[234] & b[49])^(a[233] & b[50])^(a[232] & b[51])^(a[231] & b[52])^(a[230] & b[53])^(a[229] & b[54])^(a[228] & b[55])^(a[227] & b[56])^(a[226] & b[57])^(a[225] & b[58])^(a[224] & b[59])^(a[223] & b[60])^(a[222] & b[61])^(a[221] & b[62])^(a[220] & b[63])^(a[219] & b[64])^(a[218] & b[65])^(a[217] & b[66])^(a[216] & b[67])^(a[215] & b[68])^(a[214] & b[69])^(a[213] & b[70])^(a[212] & b[71])^(a[211] & b[72])^(a[210] & b[73])^(a[209] & b[74])^(a[208] & b[75])^(a[207] & b[76])^(a[206] & b[77])^(a[205] & b[78])^(a[204] & b[79])^(a[203] & b[80])^(a[202] & b[81])^(a[201] & b[82])^(a[200] & b[83])^(a[199] & b[84])^(a[198] & b[85])^(a[197] & b[86])^(a[196] & b[87])^(a[195] & b[88])^(a[194] & b[89])^(a[193] & b[90])^(a[192] & b[91])^(a[191] & b[92])^(a[190] & b[93])^(a[189] & b[94])^(a[188] & b[95])^(a[187] & b[96])^(a[186] & b[97])^(a[185] & b[98])^(a[184] & b[99])^(a[183] & b[100])^(a[182] & b[101])^(a[181] & b[102])^(a[180] & b[103])^(a[179] & b[104])^(a[178] & b[105])^(a[177] & b[106])^(a[176] & b[107])^(a[175] & b[108])^(a[174] & b[109])^(a[173] & b[110])^(a[172] & b[111])^(a[171] & b[112])^(a[170] & b[113])^(a[169] & b[114])^(a[168] & b[115])^(a[167] & b[116])^(a[166] & b[117])^(a[165] & b[118])^(a[164] & b[119])^(a[163] & b[120])^(a[162] & b[121])^(a[161] & b[122])^(a[160] & b[123])^(a[159] & b[124])^(a[158] & b[125])^(a[157] & b[126])^(a[156] & b[127])^(a[155] & b[128])^(a[154] & b[129])^(a[153] & b[130])^(a[152] & b[131])^(a[151] & b[132])^(a[150] & b[133])^(a[149] & b[134])^(a[148] & b[135])^(a[147] & b[136])^(a[146] & b[137])^(a[145] & b[138])^(a[144] & b[139])^(a[143] & b[140])^(a[142] & b[141])^(a[141] & b[142])^(a[140] & b[143])^(a[139] & b[144])^(a[138] & b[145])^(a[137] & b[146])^(a[136] & b[147])^(a[135] & b[148])^(a[134] & b[149])^(a[133] & b[150])^(a[132] & b[151])^(a[131] & b[152])^(a[130] & b[153])^(a[129] & b[154])^(a[128] & b[155])^(a[127] & b[156])^(a[126] & b[157])^(a[125] & b[158])^(a[124] & b[159])^(a[123] & b[160])^(a[122] & b[161])^(a[121] & b[162])^(a[120] & b[163])^(a[119] & b[164])^(a[118] & b[165])^(a[117] & b[166])^(a[116] & b[167])^(a[115] & b[168])^(a[114] & b[169])^(a[113] & b[170])^(a[112] & b[171])^(a[111] & b[172])^(a[110] & b[173])^(a[109] & b[174])^(a[108] & b[175])^(a[107] & b[176])^(a[106] & b[177])^(a[105] & b[178])^(a[104] & b[179])^(a[103] & b[180])^(a[102] & b[181])^(a[101] & b[182])^(a[100] & b[183])^(a[99] & b[184])^(a[98] & b[185])^(a[97] & b[186])^(a[96] & b[187])^(a[95] & b[188])^(a[94] & b[189])^(a[93] & b[190])^(a[92] & b[191])^(a[91] & b[192])^(a[90] & b[193])^(a[89] & b[194])^(a[88] & b[195])^(a[87] & b[196])^(a[86] & b[197])^(a[85] & b[198])^(a[84] & b[199])^(a[83] & b[200])^(a[82] & b[201])^(a[81] & b[202])^(a[80] & b[203])^(a[79] & b[204])^(a[78] & b[205])^(a[77] & b[206])^(a[76] & b[207])^(a[75] & b[208])^(a[74] & b[209])^(a[73] & b[210])^(a[72] & b[211])^(a[71] & b[212])^(a[70] & b[213])^(a[69] & b[214])^(a[68] & b[215])^(a[67] & b[216])^(a[66] & b[217])^(a[65] & b[218])^(a[64] & b[219])^(a[63] & b[220])^(a[62] & b[221])^(a[61] & b[222])^(a[60] & b[223])^(a[59] & b[224])^(a[58] & b[225])^(a[57] & b[226])^(a[56] & b[227])^(a[55] & b[228])^(a[54] & b[229])^(a[53] & b[230])^(a[52] & b[231])^(a[51] & b[232])^(a[50] & b[233])^(a[49] & b[234])^(a[48] & b[235])^(a[47] & b[236])^(a[46] & b[237])^(a[45] & b[238])^(a[44] & b[239])^(a[43] & b[240])^(a[42] & b[241])^(a[41] & b[242])^(a[40] & b[243])^(a[39] & b[244])^(a[38] & b[245])^(a[37] & b[246])^(a[36] & b[247])^(a[35] & b[248])^(a[34] & b[249])^(a[33] & b[250])^(a[32] & b[251])^(a[31] & b[252])^(a[30] & b[253])^(a[29] & b[254])^(a[28] & b[255])^(a[27] & b[256])^(a[26] & b[257])^(a[25] & b[258])^(a[24] & b[259])^(a[23] & b[260])^(a[22] & b[261])^(a[21] & b[262])^(a[20] & b[263])^(a[19] & b[264])^(a[18] & b[265])^(a[17] & b[266])^(a[16] & b[267])^(a[15] & b[268])^(a[14] & b[269])^(a[13] & b[270])^(a[12] & b[271])^(a[11] & b[272])^(a[10] & b[273])^(a[9] & b[274])^(a[8] & b[275])^(a[7] & b[276])^(a[6] & b[277])^(a[5] & b[278])^(a[4] & b[279])^(a[3] & b[280])^(a[2] & b[281])^(a[1] & b[282])^(a[0] & b[283]);
assign y[284] = (a[284] & b[0])^(a[283] & b[1])^(a[282] & b[2])^(a[281] & b[3])^(a[280] & b[4])^(a[279] & b[5])^(a[278] & b[6])^(a[277] & b[7])^(a[276] & b[8])^(a[275] & b[9])^(a[274] & b[10])^(a[273] & b[11])^(a[272] & b[12])^(a[271] & b[13])^(a[270] & b[14])^(a[269] & b[15])^(a[268] & b[16])^(a[267] & b[17])^(a[266] & b[18])^(a[265] & b[19])^(a[264] & b[20])^(a[263] & b[21])^(a[262] & b[22])^(a[261] & b[23])^(a[260] & b[24])^(a[259] & b[25])^(a[258] & b[26])^(a[257] & b[27])^(a[256] & b[28])^(a[255] & b[29])^(a[254] & b[30])^(a[253] & b[31])^(a[252] & b[32])^(a[251] & b[33])^(a[250] & b[34])^(a[249] & b[35])^(a[248] & b[36])^(a[247] & b[37])^(a[246] & b[38])^(a[245] & b[39])^(a[244] & b[40])^(a[243] & b[41])^(a[242] & b[42])^(a[241] & b[43])^(a[240] & b[44])^(a[239] & b[45])^(a[238] & b[46])^(a[237] & b[47])^(a[236] & b[48])^(a[235] & b[49])^(a[234] & b[50])^(a[233] & b[51])^(a[232] & b[52])^(a[231] & b[53])^(a[230] & b[54])^(a[229] & b[55])^(a[228] & b[56])^(a[227] & b[57])^(a[226] & b[58])^(a[225] & b[59])^(a[224] & b[60])^(a[223] & b[61])^(a[222] & b[62])^(a[221] & b[63])^(a[220] & b[64])^(a[219] & b[65])^(a[218] & b[66])^(a[217] & b[67])^(a[216] & b[68])^(a[215] & b[69])^(a[214] & b[70])^(a[213] & b[71])^(a[212] & b[72])^(a[211] & b[73])^(a[210] & b[74])^(a[209] & b[75])^(a[208] & b[76])^(a[207] & b[77])^(a[206] & b[78])^(a[205] & b[79])^(a[204] & b[80])^(a[203] & b[81])^(a[202] & b[82])^(a[201] & b[83])^(a[200] & b[84])^(a[199] & b[85])^(a[198] & b[86])^(a[197] & b[87])^(a[196] & b[88])^(a[195] & b[89])^(a[194] & b[90])^(a[193] & b[91])^(a[192] & b[92])^(a[191] & b[93])^(a[190] & b[94])^(a[189] & b[95])^(a[188] & b[96])^(a[187] & b[97])^(a[186] & b[98])^(a[185] & b[99])^(a[184] & b[100])^(a[183] & b[101])^(a[182] & b[102])^(a[181] & b[103])^(a[180] & b[104])^(a[179] & b[105])^(a[178] & b[106])^(a[177] & b[107])^(a[176] & b[108])^(a[175] & b[109])^(a[174] & b[110])^(a[173] & b[111])^(a[172] & b[112])^(a[171] & b[113])^(a[170] & b[114])^(a[169] & b[115])^(a[168] & b[116])^(a[167] & b[117])^(a[166] & b[118])^(a[165] & b[119])^(a[164] & b[120])^(a[163] & b[121])^(a[162] & b[122])^(a[161] & b[123])^(a[160] & b[124])^(a[159] & b[125])^(a[158] & b[126])^(a[157] & b[127])^(a[156] & b[128])^(a[155] & b[129])^(a[154] & b[130])^(a[153] & b[131])^(a[152] & b[132])^(a[151] & b[133])^(a[150] & b[134])^(a[149] & b[135])^(a[148] & b[136])^(a[147] & b[137])^(a[146] & b[138])^(a[145] & b[139])^(a[144] & b[140])^(a[143] & b[141])^(a[142] & b[142])^(a[141] & b[143])^(a[140] & b[144])^(a[139] & b[145])^(a[138] & b[146])^(a[137] & b[147])^(a[136] & b[148])^(a[135] & b[149])^(a[134] & b[150])^(a[133] & b[151])^(a[132] & b[152])^(a[131] & b[153])^(a[130] & b[154])^(a[129] & b[155])^(a[128] & b[156])^(a[127] & b[157])^(a[126] & b[158])^(a[125] & b[159])^(a[124] & b[160])^(a[123] & b[161])^(a[122] & b[162])^(a[121] & b[163])^(a[120] & b[164])^(a[119] & b[165])^(a[118] & b[166])^(a[117] & b[167])^(a[116] & b[168])^(a[115] & b[169])^(a[114] & b[170])^(a[113] & b[171])^(a[112] & b[172])^(a[111] & b[173])^(a[110] & b[174])^(a[109] & b[175])^(a[108] & b[176])^(a[107] & b[177])^(a[106] & b[178])^(a[105] & b[179])^(a[104] & b[180])^(a[103] & b[181])^(a[102] & b[182])^(a[101] & b[183])^(a[100] & b[184])^(a[99] & b[185])^(a[98] & b[186])^(a[97] & b[187])^(a[96] & b[188])^(a[95] & b[189])^(a[94] & b[190])^(a[93] & b[191])^(a[92] & b[192])^(a[91] & b[193])^(a[90] & b[194])^(a[89] & b[195])^(a[88] & b[196])^(a[87] & b[197])^(a[86] & b[198])^(a[85] & b[199])^(a[84] & b[200])^(a[83] & b[201])^(a[82] & b[202])^(a[81] & b[203])^(a[80] & b[204])^(a[79] & b[205])^(a[78] & b[206])^(a[77] & b[207])^(a[76] & b[208])^(a[75] & b[209])^(a[74] & b[210])^(a[73] & b[211])^(a[72] & b[212])^(a[71] & b[213])^(a[70] & b[214])^(a[69] & b[215])^(a[68] & b[216])^(a[67] & b[217])^(a[66] & b[218])^(a[65] & b[219])^(a[64] & b[220])^(a[63] & b[221])^(a[62] & b[222])^(a[61] & b[223])^(a[60] & b[224])^(a[59] & b[225])^(a[58] & b[226])^(a[57] & b[227])^(a[56] & b[228])^(a[55] & b[229])^(a[54] & b[230])^(a[53] & b[231])^(a[52] & b[232])^(a[51] & b[233])^(a[50] & b[234])^(a[49] & b[235])^(a[48] & b[236])^(a[47] & b[237])^(a[46] & b[238])^(a[45] & b[239])^(a[44] & b[240])^(a[43] & b[241])^(a[42] & b[242])^(a[41] & b[243])^(a[40] & b[244])^(a[39] & b[245])^(a[38] & b[246])^(a[37] & b[247])^(a[36] & b[248])^(a[35] & b[249])^(a[34] & b[250])^(a[33] & b[251])^(a[32] & b[252])^(a[31] & b[253])^(a[30] & b[254])^(a[29] & b[255])^(a[28] & b[256])^(a[27] & b[257])^(a[26] & b[258])^(a[25] & b[259])^(a[24] & b[260])^(a[23] & b[261])^(a[22] & b[262])^(a[21] & b[263])^(a[20] & b[264])^(a[19] & b[265])^(a[18] & b[266])^(a[17] & b[267])^(a[16] & b[268])^(a[15] & b[269])^(a[14] & b[270])^(a[13] & b[271])^(a[12] & b[272])^(a[11] & b[273])^(a[10] & b[274])^(a[9] & b[275])^(a[8] & b[276])^(a[7] & b[277])^(a[6] & b[278])^(a[5] & b[279])^(a[4] & b[280])^(a[3] & b[281])^(a[2] & b[282])^(a[1] & b[283])^(a[0] & b[284]);
assign y[285] = (a[285] & b[0])^(a[284] & b[1])^(a[283] & b[2])^(a[282] & b[3])^(a[281] & b[4])^(a[280] & b[5])^(a[279] & b[6])^(a[278] & b[7])^(a[277] & b[8])^(a[276] & b[9])^(a[275] & b[10])^(a[274] & b[11])^(a[273] & b[12])^(a[272] & b[13])^(a[271] & b[14])^(a[270] & b[15])^(a[269] & b[16])^(a[268] & b[17])^(a[267] & b[18])^(a[266] & b[19])^(a[265] & b[20])^(a[264] & b[21])^(a[263] & b[22])^(a[262] & b[23])^(a[261] & b[24])^(a[260] & b[25])^(a[259] & b[26])^(a[258] & b[27])^(a[257] & b[28])^(a[256] & b[29])^(a[255] & b[30])^(a[254] & b[31])^(a[253] & b[32])^(a[252] & b[33])^(a[251] & b[34])^(a[250] & b[35])^(a[249] & b[36])^(a[248] & b[37])^(a[247] & b[38])^(a[246] & b[39])^(a[245] & b[40])^(a[244] & b[41])^(a[243] & b[42])^(a[242] & b[43])^(a[241] & b[44])^(a[240] & b[45])^(a[239] & b[46])^(a[238] & b[47])^(a[237] & b[48])^(a[236] & b[49])^(a[235] & b[50])^(a[234] & b[51])^(a[233] & b[52])^(a[232] & b[53])^(a[231] & b[54])^(a[230] & b[55])^(a[229] & b[56])^(a[228] & b[57])^(a[227] & b[58])^(a[226] & b[59])^(a[225] & b[60])^(a[224] & b[61])^(a[223] & b[62])^(a[222] & b[63])^(a[221] & b[64])^(a[220] & b[65])^(a[219] & b[66])^(a[218] & b[67])^(a[217] & b[68])^(a[216] & b[69])^(a[215] & b[70])^(a[214] & b[71])^(a[213] & b[72])^(a[212] & b[73])^(a[211] & b[74])^(a[210] & b[75])^(a[209] & b[76])^(a[208] & b[77])^(a[207] & b[78])^(a[206] & b[79])^(a[205] & b[80])^(a[204] & b[81])^(a[203] & b[82])^(a[202] & b[83])^(a[201] & b[84])^(a[200] & b[85])^(a[199] & b[86])^(a[198] & b[87])^(a[197] & b[88])^(a[196] & b[89])^(a[195] & b[90])^(a[194] & b[91])^(a[193] & b[92])^(a[192] & b[93])^(a[191] & b[94])^(a[190] & b[95])^(a[189] & b[96])^(a[188] & b[97])^(a[187] & b[98])^(a[186] & b[99])^(a[185] & b[100])^(a[184] & b[101])^(a[183] & b[102])^(a[182] & b[103])^(a[181] & b[104])^(a[180] & b[105])^(a[179] & b[106])^(a[178] & b[107])^(a[177] & b[108])^(a[176] & b[109])^(a[175] & b[110])^(a[174] & b[111])^(a[173] & b[112])^(a[172] & b[113])^(a[171] & b[114])^(a[170] & b[115])^(a[169] & b[116])^(a[168] & b[117])^(a[167] & b[118])^(a[166] & b[119])^(a[165] & b[120])^(a[164] & b[121])^(a[163] & b[122])^(a[162] & b[123])^(a[161] & b[124])^(a[160] & b[125])^(a[159] & b[126])^(a[158] & b[127])^(a[157] & b[128])^(a[156] & b[129])^(a[155] & b[130])^(a[154] & b[131])^(a[153] & b[132])^(a[152] & b[133])^(a[151] & b[134])^(a[150] & b[135])^(a[149] & b[136])^(a[148] & b[137])^(a[147] & b[138])^(a[146] & b[139])^(a[145] & b[140])^(a[144] & b[141])^(a[143] & b[142])^(a[142] & b[143])^(a[141] & b[144])^(a[140] & b[145])^(a[139] & b[146])^(a[138] & b[147])^(a[137] & b[148])^(a[136] & b[149])^(a[135] & b[150])^(a[134] & b[151])^(a[133] & b[152])^(a[132] & b[153])^(a[131] & b[154])^(a[130] & b[155])^(a[129] & b[156])^(a[128] & b[157])^(a[127] & b[158])^(a[126] & b[159])^(a[125] & b[160])^(a[124] & b[161])^(a[123] & b[162])^(a[122] & b[163])^(a[121] & b[164])^(a[120] & b[165])^(a[119] & b[166])^(a[118] & b[167])^(a[117] & b[168])^(a[116] & b[169])^(a[115] & b[170])^(a[114] & b[171])^(a[113] & b[172])^(a[112] & b[173])^(a[111] & b[174])^(a[110] & b[175])^(a[109] & b[176])^(a[108] & b[177])^(a[107] & b[178])^(a[106] & b[179])^(a[105] & b[180])^(a[104] & b[181])^(a[103] & b[182])^(a[102] & b[183])^(a[101] & b[184])^(a[100] & b[185])^(a[99] & b[186])^(a[98] & b[187])^(a[97] & b[188])^(a[96] & b[189])^(a[95] & b[190])^(a[94] & b[191])^(a[93] & b[192])^(a[92] & b[193])^(a[91] & b[194])^(a[90] & b[195])^(a[89] & b[196])^(a[88] & b[197])^(a[87] & b[198])^(a[86] & b[199])^(a[85] & b[200])^(a[84] & b[201])^(a[83] & b[202])^(a[82] & b[203])^(a[81] & b[204])^(a[80] & b[205])^(a[79] & b[206])^(a[78] & b[207])^(a[77] & b[208])^(a[76] & b[209])^(a[75] & b[210])^(a[74] & b[211])^(a[73] & b[212])^(a[72] & b[213])^(a[71] & b[214])^(a[70] & b[215])^(a[69] & b[216])^(a[68] & b[217])^(a[67] & b[218])^(a[66] & b[219])^(a[65] & b[220])^(a[64] & b[221])^(a[63] & b[222])^(a[62] & b[223])^(a[61] & b[224])^(a[60] & b[225])^(a[59] & b[226])^(a[58] & b[227])^(a[57] & b[228])^(a[56] & b[229])^(a[55] & b[230])^(a[54] & b[231])^(a[53] & b[232])^(a[52] & b[233])^(a[51] & b[234])^(a[50] & b[235])^(a[49] & b[236])^(a[48] & b[237])^(a[47] & b[238])^(a[46] & b[239])^(a[45] & b[240])^(a[44] & b[241])^(a[43] & b[242])^(a[42] & b[243])^(a[41] & b[244])^(a[40] & b[245])^(a[39] & b[246])^(a[38] & b[247])^(a[37] & b[248])^(a[36] & b[249])^(a[35] & b[250])^(a[34] & b[251])^(a[33] & b[252])^(a[32] & b[253])^(a[31] & b[254])^(a[30] & b[255])^(a[29] & b[256])^(a[28] & b[257])^(a[27] & b[258])^(a[26] & b[259])^(a[25] & b[260])^(a[24] & b[261])^(a[23] & b[262])^(a[22] & b[263])^(a[21] & b[264])^(a[20] & b[265])^(a[19] & b[266])^(a[18] & b[267])^(a[17] & b[268])^(a[16] & b[269])^(a[15] & b[270])^(a[14] & b[271])^(a[13] & b[272])^(a[12] & b[273])^(a[11] & b[274])^(a[10] & b[275])^(a[9] & b[276])^(a[8] & b[277])^(a[7] & b[278])^(a[6] & b[279])^(a[5] & b[280])^(a[4] & b[281])^(a[3] & b[282])^(a[2] & b[283])^(a[1] & b[284])^(a[0] & b[285]);
assign y[286] = (a[286] & b[0])^(a[285] & b[1])^(a[284] & b[2])^(a[283] & b[3])^(a[282] & b[4])^(a[281] & b[5])^(a[280] & b[6])^(a[279] & b[7])^(a[278] & b[8])^(a[277] & b[9])^(a[276] & b[10])^(a[275] & b[11])^(a[274] & b[12])^(a[273] & b[13])^(a[272] & b[14])^(a[271] & b[15])^(a[270] & b[16])^(a[269] & b[17])^(a[268] & b[18])^(a[267] & b[19])^(a[266] & b[20])^(a[265] & b[21])^(a[264] & b[22])^(a[263] & b[23])^(a[262] & b[24])^(a[261] & b[25])^(a[260] & b[26])^(a[259] & b[27])^(a[258] & b[28])^(a[257] & b[29])^(a[256] & b[30])^(a[255] & b[31])^(a[254] & b[32])^(a[253] & b[33])^(a[252] & b[34])^(a[251] & b[35])^(a[250] & b[36])^(a[249] & b[37])^(a[248] & b[38])^(a[247] & b[39])^(a[246] & b[40])^(a[245] & b[41])^(a[244] & b[42])^(a[243] & b[43])^(a[242] & b[44])^(a[241] & b[45])^(a[240] & b[46])^(a[239] & b[47])^(a[238] & b[48])^(a[237] & b[49])^(a[236] & b[50])^(a[235] & b[51])^(a[234] & b[52])^(a[233] & b[53])^(a[232] & b[54])^(a[231] & b[55])^(a[230] & b[56])^(a[229] & b[57])^(a[228] & b[58])^(a[227] & b[59])^(a[226] & b[60])^(a[225] & b[61])^(a[224] & b[62])^(a[223] & b[63])^(a[222] & b[64])^(a[221] & b[65])^(a[220] & b[66])^(a[219] & b[67])^(a[218] & b[68])^(a[217] & b[69])^(a[216] & b[70])^(a[215] & b[71])^(a[214] & b[72])^(a[213] & b[73])^(a[212] & b[74])^(a[211] & b[75])^(a[210] & b[76])^(a[209] & b[77])^(a[208] & b[78])^(a[207] & b[79])^(a[206] & b[80])^(a[205] & b[81])^(a[204] & b[82])^(a[203] & b[83])^(a[202] & b[84])^(a[201] & b[85])^(a[200] & b[86])^(a[199] & b[87])^(a[198] & b[88])^(a[197] & b[89])^(a[196] & b[90])^(a[195] & b[91])^(a[194] & b[92])^(a[193] & b[93])^(a[192] & b[94])^(a[191] & b[95])^(a[190] & b[96])^(a[189] & b[97])^(a[188] & b[98])^(a[187] & b[99])^(a[186] & b[100])^(a[185] & b[101])^(a[184] & b[102])^(a[183] & b[103])^(a[182] & b[104])^(a[181] & b[105])^(a[180] & b[106])^(a[179] & b[107])^(a[178] & b[108])^(a[177] & b[109])^(a[176] & b[110])^(a[175] & b[111])^(a[174] & b[112])^(a[173] & b[113])^(a[172] & b[114])^(a[171] & b[115])^(a[170] & b[116])^(a[169] & b[117])^(a[168] & b[118])^(a[167] & b[119])^(a[166] & b[120])^(a[165] & b[121])^(a[164] & b[122])^(a[163] & b[123])^(a[162] & b[124])^(a[161] & b[125])^(a[160] & b[126])^(a[159] & b[127])^(a[158] & b[128])^(a[157] & b[129])^(a[156] & b[130])^(a[155] & b[131])^(a[154] & b[132])^(a[153] & b[133])^(a[152] & b[134])^(a[151] & b[135])^(a[150] & b[136])^(a[149] & b[137])^(a[148] & b[138])^(a[147] & b[139])^(a[146] & b[140])^(a[145] & b[141])^(a[144] & b[142])^(a[143] & b[143])^(a[142] & b[144])^(a[141] & b[145])^(a[140] & b[146])^(a[139] & b[147])^(a[138] & b[148])^(a[137] & b[149])^(a[136] & b[150])^(a[135] & b[151])^(a[134] & b[152])^(a[133] & b[153])^(a[132] & b[154])^(a[131] & b[155])^(a[130] & b[156])^(a[129] & b[157])^(a[128] & b[158])^(a[127] & b[159])^(a[126] & b[160])^(a[125] & b[161])^(a[124] & b[162])^(a[123] & b[163])^(a[122] & b[164])^(a[121] & b[165])^(a[120] & b[166])^(a[119] & b[167])^(a[118] & b[168])^(a[117] & b[169])^(a[116] & b[170])^(a[115] & b[171])^(a[114] & b[172])^(a[113] & b[173])^(a[112] & b[174])^(a[111] & b[175])^(a[110] & b[176])^(a[109] & b[177])^(a[108] & b[178])^(a[107] & b[179])^(a[106] & b[180])^(a[105] & b[181])^(a[104] & b[182])^(a[103] & b[183])^(a[102] & b[184])^(a[101] & b[185])^(a[100] & b[186])^(a[99] & b[187])^(a[98] & b[188])^(a[97] & b[189])^(a[96] & b[190])^(a[95] & b[191])^(a[94] & b[192])^(a[93] & b[193])^(a[92] & b[194])^(a[91] & b[195])^(a[90] & b[196])^(a[89] & b[197])^(a[88] & b[198])^(a[87] & b[199])^(a[86] & b[200])^(a[85] & b[201])^(a[84] & b[202])^(a[83] & b[203])^(a[82] & b[204])^(a[81] & b[205])^(a[80] & b[206])^(a[79] & b[207])^(a[78] & b[208])^(a[77] & b[209])^(a[76] & b[210])^(a[75] & b[211])^(a[74] & b[212])^(a[73] & b[213])^(a[72] & b[214])^(a[71] & b[215])^(a[70] & b[216])^(a[69] & b[217])^(a[68] & b[218])^(a[67] & b[219])^(a[66] & b[220])^(a[65] & b[221])^(a[64] & b[222])^(a[63] & b[223])^(a[62] & b[224])^(a[61] & b[225])^(a[60] & b[226])^(a[59] & b[227])^(a[58] & b[228])^(a[57] & b[229])^(a[56] & b[230])^(a[55] & b[231])^(a[54] & b[232])^(a[53] & b[233])^(a[52] & b[234])^(a[51] & b[235])^(a[50] & b[236])^(a[49] & b[237])^(a[48] & b[238])^(a[47] & b[239])^(a[46] & b[240])^(a[45] & b[241])^(a[44] & b[242])^(a[43] & b[243])^(a[42] & b[244])^(a[41] & b[245])^(a[40] & b[246])^(a[39] & b[247])^(a[38] & b[248])^(a[37] & b[249])^(a[36] & b[250])^(a[35] & b[251])^(a[34] & b[252])^(a[33] & b[253])^(a[32] & b[254])^(a[31] & b[255])^(a[30] & b[256])^(a[29] & b[257])^(a[28] & b[258])^(a[27] & b[259])^(a[26] & b[260])^(a[25] & b[261])^(a[24] & b[262])^(a[23] & b[263])^(a[22] & b[264])^(a[21] & b[265])^(a[20] & b[266])^(a[19] & b[267])^(a[18] & b[268])^(a[17] & b[269])^(a[16] & b[270])^(a[15] & b[271])^(a[14] & b[272])^(a[13] & b[273])^(a[12] & b[274])^(a[11] & b[275])^(a[10] & b[276])^(a[9] & b[277])^(a[8] & b[278])^(a[7] & b[279])^(a[6] & b[280])^(a[5] & b[281])^(a[4] & b[282])^(a[3] & b[283])^(a[2] & b[284])^(a[1] & b[285])^(a[0] & b[286]);
assign y[287] = (a[287] & b[0])^(a[286] & b[1])^(a[285] & b[2])^(a[284] & b[3])^(a[283] & b[4])^(a[282] & b[5])^(a[281] & b[6])^(a[280] & b[7])^(a[279] & b[8])^(a[278] & b[9])^(a[277] & b[10])^(a[276] & b[11])^(a[275] & b[12])^(a[274] & b[13])^(a[273] & b[14])^(a[272] & b[15])^(a[271] & b[16])^(a[270] & b[17])^(a[269] & b[18])^(a[268] & b[19])^(a[267] & b[20])^(a[266] & b[21])^(a[265] & b[22])^(a[264] & b[23])^(a[263] & b[24])^(a[262] & b[25])^(a[261] & b[26])^(a[260] & b[27])^(a[259] & b[28])^(a[258] & b[29])^(a[257] & b[30])^(a[256] & b[31])^(a[255] & b[32])^(a[254] & b[33])^(a[253] & b[34])^(a[252] & b[35])^(a[251] & b[36])^(a[250] & b[37])^(a[249] & b[38])^(a[248] & b[39])^(a[247] & b[40])^(a[246] & b[41])^(a[245] & b[42])^(a[244] & b[43])^(a[243] & b[44])^(a[242] & b[45])^(a[241] & b[46])^(a[240] & b[47])^(a[239] & b[48])^(a[238] & b[49])^(a[237] & b[50])^(a[236] & b[51])^(a[235] & b[52])^(a[234] & b[53])^(a[233] & b[54])^(a[232] & b[55])^(a[231] & b[56])^(a[230] & b[57])^(a[229] & b[58])^(a[228] & b[59])^(a[227] & b[60])^(a[226] & b[61])^(a[225] & b[62])^(a[224] & b[63])^(a[223] & b[64])^(a[222] & b[65])^(a[221] & b[66])^(a[220] & b[67])^(a[219] & b[68])^(a[218] & b[69])^(a[217] & b[70])^(a[216] & b[71])^(a[215] & b[72])^(a[214] & b[73])^(a[213] & b[74])^(a[212] & b[75])^(a[211] & b[76])^(a[210] & b[77])^(a[209] & b[78])^(a[208] & b[79])^(a[207] & b[80])^(a[206] & b[81])^(a[205] & b[82])^(a[204] & b[83])^(a[203] & b[84])^(a[202] & b[85])^(a[201] & b[86])^(a[200] & b[87])^(a[199] & b[88])^(a[198] & b[89])^(a[197] & b[90])^(a[196] & b[91])^(a[195] & b[92])^(a[194] & b[93])^(a[193] & b[94])^(a[192] & b[95])^(a[191] & b[96])^(a[190] & b[97])^(a[189] & b[98])^(a[188] & b[99])^(a[187] & b[100])^(a[186] & b[101])^(a[185] & b[102])^(a[184] & b[103])^(a[183] & b[104])^(a[182] & b[105])^(a[181] & b[106])^(a[180] & b[107])^(a[179] & b[108])^(a[178] & b[109])^(a[177] & b[110])^(a[176] & b[111])^(a[175] & b[112])^(a[174] & b[113])^(a[173] & b[114])^(a[172] & b[115])^(a[171] & b[116])^(a[170] & b[117])^(a[169] & b[118])^(a[168] & b[119])^(a[167] & b[120])^(a[166] & b[121])^(a[165] & b[122])^(a[164] & b[123])^(a[163] & b[124])^(a[162] & b[125])^(a[161] & b[126])^(a[160] & b[127])^(a[159] & b[128])^(a[158] & b[129])^(a[157] & b[130])^(a[156] & b[131])^(a[155] & b[132])^(a[154] & b[133])^(a[153] & b[134])^(a[152] & b[135])^(a[151] & b[136])^(a[150] & b[137])^(a[149] & b[138])^(a[148] & b[139])^(a[147] & b[140])^(a[146] & b[141])^(a[145] & b[142])^(a[144] & b[143])^(a[143] & b[144])^(a[142] & b[145])^(a[141] & b[146])^(a[140] & b[147])^(a[139] & b[148])^(a[138] & b[149])^(a[137] & b[150])^(a[136] & b[151])^(a[135] & b[152])^(a[134] & b[153])^(a[133] & b[154])^(a[132] & b[155])^(a[131] & b[156])^(a[130] & b[157])^(a[129] & b[158])^(a[128] & b[159])^(a[127] & b[160])^(a[126] & b[161])^(a[125] & b[162])^(a[124] & b[163])^(a[123] & b[164])^(a[122] & b[165])^(a[121] & b[166])^(a[120] & b[167])^(a[119] & b[168])^(a[118] & b[169])^(a[117] & b[170])^(a[116] & b[171])^(a[115] & b[172])^(a[114] & b[173])^(a[113] & b[174])^(a[112] & b[175])^(a[111] & b[176])^(a[110] & b[177])^(a[109] & b[178])^(a[108] & b[179])^(a[107] & b[180])^(a[106] & b[181])^(a[105] & b[182])^(a[104] & b[183])^(a[103] & b[184])^(a[102] & b[185])^(a[101] & b[186])^(a[100] & b[187])^(a[99] & b[188])^(a[98] & b[189])^(a[97] & b[190])^(a[96] & b[191])^(a[95] & b[192])^(a[94] & b[193])^(a[93] & b[194])^(a[92] & b[195])^(a[91] & b[196])^(a[90] & b[197])^(a[89] & b[198])^(a[88] & b[199])^(a[87] & b[200])^(a[86] & b[201])^(a[85] & b[202])^(a[84] & b[203])^(a[83] & b[204])^(a[82] & b[205])^(a[81] & b[206])^(a[80] & b[207])^(a[79] & b[208])^(a[78] & b[209])^(a[77] & b[210])^(a[76] & b[211])^(a[75] & b[212])^(a[74] & b[213])^(a[73] & b[214])^(a[72] & b[215])^(a[71] & b[216])^(a[70] & b[217])^(a[69] & b[218])^(a[68] & b[219])^(a[67] & b[220])^(a[66] & b[221])^(a[65] & b[222])^(a[64] & b[223])^(a[63] & b[224])^(a[62] & b[225])^(a[61] & b[226])^(a[60] & b[227])^(a[59] & b[228])^(a[58] & b[229])^(a[57] & b[230])^(a[56] & b[231])^(a[55] & b[232])^(a[54] & b[233])^(a[53] & b[234])^(a[52] & b[235])^(a[51] & b[236])^(a[50] & b[237])^(a[49] & b[238])^(a[48] & b[239])^(a[47] & b[240])^(a[46] & b[241])^(a[45] & b[242])^(a[44] & b[243])^(a[43] & b[244])^(a[42] & b[245])^(a[41] & b[246])^(a[40] & b[247])^(a[39] & b[248])^(a[38] & b[249])^(a[37] & b[250])^(a[36] & b[251])^(a[35] & b[252])^(a[34] & b[253])^(a[33] & b[254])^(a[32] & b[255])^(a[31] & b[256])^(a[30] & b[257])^(a[29] & b[258])^(a[28] & b[259])^(a[27] & b[260])^(a[26] & b[261])^(a[25] & b[262])^(a[24] & b[263])^(a[23] & b[264])^(a[22] & b[265])^(a[21] & b[266])^(a[20] & b[267])^(a[19] & b[268])^(a[18] & b[269])^(a[17] & b[270])^(a[16] & b[271])^(a[15] & b[272])^(a[14] & b[273])^(a[13] & b[274])^(a[12] & b[275])^(a[11] & b[276])^(a[10] & b[277])^(a[9] & b[278])^(a[8] & b[279])^(a[7] & b[280])^(a[6] & b[281])^(a[5] & b[282])^(a[4] & b[283])^(a[3] & b[284])^(a[2] & b[285])^(a[1] & b[286])^(a[0] & b[287]);
assign y[288] = (a[288] & b[0])^(a[287] & b[1])^(a[286] & b[2])^(a[285] & b[3])^(a[284] & b[4])^(a[283] & b[5])^(a[282] & b[6])^(a[281] & b[7])^(a[280] & b[8])^(a[279] & b[9])^(a[278] & b[10])^(a[277] & b[11])^(a[276] & b[12])^(a[275] & b[13])^(a[274] & b[14])^(a[273] & b[15])^(a[272] & b[16])^(a[271] & b[17])^(a[270] & b[18])^(a[269] & b[19])^(a[268] & b[20])^(a[267] & b[21])^(a[266] & b[22])^(a[265] & b[23])^(a[264] & b[24])^(a[263] & b[25])^(a[262] & b[26])^(a[261] & b[27])^(a[260] & b[28])^(a[259] & b[29])^(a[258] & b[30])^(a[257] & b[31])^(a[256] & b[32])^(a[255] & b[33])^(a[254] & b[34])^(a[253] & b[35])^(a[252] & b[36])^(a[251] & b[37])^(a[250] & b[38])^(a[249] & b[39])^(a[248] & b[40])^(a[247] & b[41])^(a[246] & b[42])^(a[245] & b[43])^(a[244] & b[44])^(a[243] & b[45])^(a[242] & b[46])^(a[241] & b[47])^(a[240] & b[48])^(a[239] & b[49])^(a[238] & b[50])^(a[237] & b[51])^(a[236] & b[52])^(a[235] & b[53])^(a[234] & b[54])^(a[233] & b[55])^(a[232] & b[56])^(a[231] & b[57])^(a[230] & b[58])^(a[229] & b[59])^(a[228] & b[60])^(a[227] & b[61])^(a[226] & b[62])^(a[225] & b[63])^(a[224] & b[64])^(a[223] & b[65])^(a[222] & b[66])^(a[221] & b[67])^(a[220] & b[68])^(a[219] & b[69])^(a[218] & b[70])^(a[217] & b[71])^(a[216] & b[72])^(a[215] & b[73])^(a[214] & b[74])^(a[213] & b[75])^(a[212] & b[76])^(a[211] & b[77])^(a[210] & b[78])^(a[209] & b[79])^(a[208] & b[80])^(a[207] & b[81])^(a[206] & b[82])^(a[205] & b[83])^(a[204] & b[84])^(a[203] & b[85])^(a[202] & b[86])^(a[201] & b[87])^(a[200] & b[88])^(a[199] & b[89])^(a[198] & b[90])^(a[197] & b[91])^(a[196] & b[92])^(a[195] & b[93])^(a[194] & b[94])^(a[193] & b[95])^(a[192] & b[96])^(a[191] & b[97])^(a[190] & b[98])^(a[189] & b[99])^(a[188] & b[100])^(a[187] & b[101])^(a[186] & b[102])^(a[185] & b[103])^(a[184] & b[104])^(a[183] & b[105])^(a[182] & b[106])^(a[181] & b[107])^(a[180] & b[108])^(a[179] & b[109])^(a[178] & b[110])^(a[177] & b[111])^(a[176] & b[112])^(a[175] & b[113])^(a[174] & b[114])^(a[173] & b[115])^(a[172] & b[116])^(a[171] & b[117])^(a[170] & b[118])^(a[169] & b[119])^(a[168] & b[120])^(a[167] & b[121])^(a[166] & b[122])^(a[165] & b[123])^(a[164] & b[124])^(a[163] & b[125])^(a[162] & b[126])^(a[161] & b[127])^(a[160] & b[128])^(a[159] & b[129])^(a[158] & b[130])^(a[157] & b[131])^(a[156] & b[132])^(a[155] & b[133])^(a[154] & b[134])^(a[153] & b[135])^(a[152] & b[136])^(a[151] & b[137])^(a[150] & b[138])^(a[149] & b[139])^(a[148] & b[140])^(a[147] & b[141])^(a[146] & b[142])^(a[145] & b[143])^(a[144] & b[144])^(a[143] & b[145])^(a[142] & b[146])^(a[141] & b[147])^(a[140] & b[148])^(a[139] & b[149])^(a[138] & b[150])^(a[137] & b[151])^(a[136] & b[152])^(a[135] & b[153])^(a[134] & b[154])^(a[133] & b[155])^(a[132] & b[156])^(a[131] & b[157])^(a[130] & b[158])^(a[129] & b[159])^(a[128] & b[160])^(a[127] & b[161])^(a[126] & b[162])^(a[125] & b[163])^(a[124] & b[164])^(a[123] & b[165])^(a[122] & b[166])^(a[121] & b[167])^(a[120] & b[168])^(a[119] & b[169])^(a[118] & b[170])^(a[117] & b[171])^(a[116] & b[172])^(a[115] & b[173])^(a[114] & b[174])^(a[113] & b[175])^(a[112] & b[176])^(a[111] & b[177])^(a[110] & b[178])^(a[109] & b[179])^(a[108] & b[180])^(a[107] & b[181])^(a[106] & b[182])^(a[105] & b[183])^(a[104] & b[184])^(a[103] & b[185])^(a[102] & b[186])^(a[101] & b[187])^(a[100] & b[188])^(a[99] & b[189])^(a[98] & b[190])^(a[97] & b[191])^(a[96] & b[192])^(a[95] & b[193])^(a[94] & b[194])^(a[93] & b[195])^(a[92] & b[196])^(a[91] & b[197])^(a[90] & b[198])^(a[89] & b[199])^(a[88] & b[200])^(a[87] & b[201])^(a[86] & b[202])^(a[85] & b[203])^(a[84] & b[204])^(a[83] & b[205])^(a[82] & b[206])^(a[81] & b[207])^(a[80] & b[208])^(a[79] & b[209])^(a[78] & b[210])^(a[77] & b[211])^(a[76] & b[212])^(a[75] & b[213])^(a[74] & b[214])^(a[73] & b[215])^(a[72] & b[216])^(a[71] & b[217])^(a[70] & b[218])^(a[69] & b[219])^(a[68] & b[220])^(a[67] & b[221])^(a[66] & b[222])^(a[65] & b[223])^(a[64] & b[224])^(a[63] & b[225])^(a[62] & b[226])^(a[61] & b[227])^(a[60] & b[228])^(a[59] & b[229])^(a[58] & b[230])^(a[57] & b[231])^(a[56] & b[232])^(a[55] & b[233])^(a[54] & b[234])^(a[53] & b[235])^(a[52] & b[236])^(a[51] & b[237])^(a[50] & b[238])^(a[49] & b[239])^(a[48] & b[240])^(a[47] & b[241])^(a[46] & b[242])^(a[45] & b[243])^(a[44] & b[244])^(a[43] & b[245])^(a[42] & b[246])^(a[41] & b[247])^(a[40] & b[248])^(a[39] & b[249])^(a[38] & b[250])^(a[37] & b[251])^(a[36] & b[252])^(a[35] & b[253])^(a[34] & b[254])^(a[33] & b[255])^(a[32] & b[256])^(a[31] & b[257])^(a[30] & b[258])^(a[29] & b[259])^(a[28] & b[260])^(a[27] & b[261])^(a[26] & b[262])^(a[25] & b[263])^(a[24] & b[264])^(a[23] & b[265])^(a[22] & b[266])^(a[21] & b[267])^(a[20] & b[268])^(a[19] & b[269])^(a[18] & b[270])^(a[17] & b[271])^(a[16] & b[272])^(a[15] & b[273])^(a[14] & b[274])^(a[13] & b[275])^(a[12] & b[276])^(a[11] & b[277])^(a[10] & b[278])^(a[9] & b[279])^(a[8] & b[280])^(a[7] & b[281])^(a[6] & b[282])^(a[5] & b[283])^(a[4] & b[284])^(a[3] & b[285])^(a[2] & b[286])^(a[1] & b[287])^(a[0] & b[288]);
assign y[289] = (a[289] & b[0])^(a[288] & b[1])^(a[287] & b[2])^(a[286] & b[3])^(a[285] & b[4])^(a[284] & b[5])^(a[283] & b[6])^(a[282] & b[7])^(a[281] & b[8])^(a[280] & b[9])^(a[279] & b[10])^(a[278] & b[11])^(a[277] & b[12])^(a[276] & b[13])^(a[275] & b[14])^(a[274] & b[15])^(a[273] & b[16])^(a[272] & b[17])^(a[271] & b[18])^(a[270] & b[19])^(a[269] & b[20])^(a[268] & b[21])^(a[267] & b[22])^(a[266] & b[23])^(a[265] & b[24])^(a[264] & b[25])^(a[263] & b[26])^(a[262] & b[27])^(a[261] & b[28])^(a[260] & b[29])^(a[259] & b[30])^(a[258] & b[31])^(a[257] & b[32])^(a[256] & b[33])^(a[255] & b[34])^(a[254] & b[35])^(a[253] & b[36])^(a[252] & b[37])^(a[251] & b[38])^(a[250] & b[39])^(a[249] & b[40])^(a[248] & b[41])^(a[247] & b[42])^(a[246] & b[43])^(a[245] & b[44])^(a[244] & b[45])^(a[243] & b[46])^(a[242] & b[47])^(a[241] & b[48])^(a[240] & b[49])^(a[239] & b[50])^(a[238] & b[51])^(a[237] & b[52])^(a[236] & b[53])^(a[235] & b[54])^(a[234] & b[55])^(a[233] & b[56])^(a[232] & b[57])^(a[231] & b[58])^(a[230] & b[59])^(a[229] & b[60])^(a[228] & b[61])^(a[227] & b[62])^(a[226] & b[63])^(a[225] & b[64])^(a[224] & b[65])^(a[223] & b[66])^(a[222] & b[67])^(a[221] & b[68])^(a[220] & b[69])^(a[219] & b[70])^(a[218] & b[71])^(a[217] & b[72])^(a[216] & b[73])^(a[215] & b[74])^(a[214] & b[75])^(a[213] & b[76])^(a[212] & b[77])^(a[211] & b[78])^(a[210] & b[79])^(a[209] & b[80])^(a[208] & b[81])^(a[207] & b[82])^(a[206] & b[83])^(a[205] & b[84])^(a[204] & b[85])^(a[203] & b[86])^(a[202] & b[87])^(a[201] & b[88])^(a[200] & b[89])^(a[199] & b[90])^(a[198] & b[91])^(a[197] & b[92])^(a[196] & b[93])^(a[195] & b[94])^(a[194] & b[95])^(a[193] & b[96])^(a[192] & b[97])^(a[191] & b[98])^(a[190] & b[99])^(a[189] & b[100])^(a[188] & b[101])^(a[187] & b[102])^(a[186] & b[103])^(a[185] & b[104])^(a[184] & b[105])^(a[183] & b[106])^(a[182] & b[107])^(a[181] & b[108])^(a[180] & b[109])^(a[179] & b[110])^(a[178] & b[111])^(a[177] & b[112])^(a[176] & b[113])^(a[175] & b[114])^(a[174] & b[115])^(a[173] & b[116])^(a[172] & b[117])^(a[171] & b[118])^(a[170] & b[119])^(a[169] & b[120])^(a[168] & b[121])^(a[167] & b[122])^(a[166] & b[123])^(a[165] & b[124])^(a[164] & b[125])^(a[163] & b[126])^(a[162] & b[127])^(a[161] & b[128])^(a[160] & b[129])^(a[159] & b[130])^(a[158] & b[131])^(a[157] & b[132])^(a[156] & b[133])^(a[155] & b[134])^(a[154] & b[135])^(a[153] & b[136])^(a[152] & b[137])^(a[151] & b[138])^(a[150] & b[139])^(a[149] & b[140])^(a[148] & b[141])^(a[147] & b[142])^(a[146] & b[143])^(a[145] & b[144])^(a[144] & b[145])^(a[143] & b[146])^(a[142] & b[147])^(a[141] & b[148])^(a[140] & b[149])^(a[139] & b[150])^(a[138] & b[151])^(a[137] & b[152])^(a[136] & b[153])^(a[135] & b[154])^(a[134] & b[155])^(a[133] & b[156])^(a[132] & b[157])^(a[131] & b[158])^(a[130] & b[159])^(a[129] & b[160])^(a[128] & b[161])^(a[127] & b[162])^(a[126] & b[163])^(a[125] & b[164])^(a[124] & b[165])^(a[123] & b[166])^(a[122] & b[167])^(a[121] & b[168])^(a[120] & b[169])^(a[119] & b[170])^(a[118] & b[171])^(a[117] & b[172])^(a[116] & b[173])^(a[115] & b[174])^(a[114] & b[175])^(a[113] & b[176])^(a[112] & b[177])^(a[111] & b[178])^(a[110] & b[179])^(a[109] & b[180])^(a[108] & b[181])^(a[107] & b[182])^(a[106] & b[183])^(a[105] & b[184])^(a[104] & b[185])^(a[103] & b[186])^(a[102] & b[187])^(a[101] & b[188])^(a[100] & b[189])^(a[99] & b[190])^(a[98] & b[191])^(a[97] & b[192])^(a[96] & b[193])^(a[95] & b[194])^(a[94] & b[195])^(a[93] & b[196])^(a[92] & b[197])^(a[91] & b[198])^(a[90] & b[199])^(a[89] & b[200])^(a[88] & b[201])^(a[87] & b[202])^(a[86] & b[203])^(a[85] & b[204])^(a[84] & b[205])^(a[83] & b[206])^(a[82] & b[207])^(a[81] & b[208])^(a[80] & b[209])^(a[79] & b[210])^(a[78] & b[211])^(a[77] & b[212])^(a[76] & b[213])^(a[75] & b[214])^(a[74] & b[215])^(a[73] & b[216])^(a[72] & b[217])^(a[71] & b[218])^(a[70] & b[219])^(a[69] & b[220])^(a[68] & b[221])^(a[67] & b[222])^(a[66] & b[223])^(a[65] & b[224])^(a[64] & b[225])^(a[63] & b[226])^(a[62] & b[227])^(a[61] & b[228])^(a[60] & b[229])^(a[59] & b[230])^(a[58] & b[231])^(a[57] & b[232])^(a[56] & b[233])^(a[55] & b[234])^(a[54] & b[235])^(a[53] & b[236])^(a[52] & b[237])^(a[51] & b[238])^(a[50] & b[239])^(a[49] & b[240])^(a[48] & b[241])^(a[47] & b[242])^(a[46] & b[243])^(a[45] & b[244])^(a[44] & b[245])^(a[43] & b[246])^(a[42] & b[247])^(a[41] & b[248])^(a[40] & b[249])^(a[39] & b[250])^(a[38] & b[251])^(a[37] & b[252])^(a[36] & b[253])^(a[35] & b[254])^(a[34] & b[255])^(a[33] & b[256])^(a[32] & b[257])^(a[31] & b[258])^(a[30] & b[259])^(a[29] & b[260])^(a[28] & b[261])^(a[27] & b[262])^(a[26] & b[263])^(a[25] & b[264])^(a[24] & b[265])^(a[23] & b[266])^(a[22] & b[267])^(a[21] & b[268])^(a[20] & b[269])^(a[19] & b[270])^(a[18] & b[271])^(a[17] & b[272])^(a[16] & b[273])^(a[15] & b[274])^(a[14] & b[275])^(a[13] & b[276])^(a[12] & b[277])^(a[11] & b[278])^(a[10] & b[279])^(a[9] & b[280])^(a[8] & b[281])^(a[7] & b[282])^(a[6] & b[283])^(a[5] & b[284])^(a[4] & b[285])^(a[3] & b[286])^(a[2] & b[287])^(a[1] & b[288])^(a[0] & b[289]);
assign y[290] = (a[290] & b[0])^(a[289] & b[1])^(a[288] & b[2])^(a[287] & b[3])^(a[286] & b[4])^(a[285] & b[5])^(a[284] & b[6])^(a[283] & b[7])^(a[282] & b[8])^(a[281] & b[9])^(a[280] & b[10])^(a[279] & b[11])^(a[278] & b[12])^(a[277] & b[13])^(a[276] & b[14])^(a[275] & b[15])^(a[274] & b[16])^(a[273] & b[17])^(a[272] & b[18])^(a[271] & b[19])^(a[270] & b[20])^(a[269] & b[21])^(a[268] & b[22])^(a[267] & b[23])^(a[266] & b[24])^(a[265] & b[25])^(a[264] & b[26])^(a[263] & b[27])^(a[262] & b[28])^(a[261] & b[29])^(a[260] & b[30])^(a[259] & b[31])^(a[258] & b[32])^(a[257] & b[33])^(a[256] & b[34])^(a[255] & b[35])^(a[254] & b[36])^(a[253] & b[37])^(a[252] & b[38])^(a[251] & b[39])^(a[250] & b[40])^(a[249] & b[41])^(a[248] & b[42])^(a[247] & b[43])^(a[246] & b[44])^(a[245] & b[45])^(a[244] & b[46])^(a[243] & b[47])^(a[242] & b[48])^(a[241] & b[49])^(a[240] & b[50])^(a[239] & b[51])^(a[238] & b[52])^(a[237] & b[53])^(a[236] & b[54])^(a[235] & b[55])^(a[234] & b[56])^(a[233] & b[57])^(a[232] & b[58])^(a[231] & b[59])^(a[230] & b[60])^(a[229] & b[61])^(a[228] & b[62])^(a[227] & b[63])^(a[226] & b[64])^(a[225] & b[65])^(a[224] & b[66])^(a[223] & b[67])^(a[222] & b[68])^(a[221] & b[69])^(a[220] & b[70])^(a[219] & b[71])^(a[218] & b[72])^(a[217] & b[73])^(a[216] & b[74])^(a[215] & b[75])^(a[214] & b[76])^(a[213] & b[77])^(a[212] & b[78])^(a[211] & b[79])^(a[210] & b[80])^(a[209] & b[81])^(a[208] & b[82])^(a[207] & b[83])^(a[206] & b[84])^(a[205] & b[85])^(a[204] & b[86])^(a[203] & b[87])^(a[202] & b[88])^(a[201] & b[89])^(a[200] & b[90])^(a[199] & b[91])^(a[198] & b[92])^(a[197] & b[93])^(a[196] & b[94])^(a[195] & b[95])^(a[194] & b[96])^(a[193] & b[97])^(a[192] & b[98])^(a[191] & b[99])^(a[190] & b[100])^(a[189] & b[101])^(a[188] & b[102])^(a[187] & b[103])^(a[186] & b[104])^(a[185] & b[105])^(a[184] & b[106])^(a[183] & b[107])^(a[182] & b[108])^(a[181] & b[109])^(a[180] & b[110])^(a[179] & b[111])^(a[178] & b[112])^(a[177] & b[113])^(a[176] & b[114])^(a[175] & b[115])^(a[174] & b[116])^(a[173] & b[117])^(a[172] & b[118])^(a[171] & b[119])^(a[170] & b[120])^(a[169] & b[121])^(a[168] & b[122])^(a[167] & b[123])^(a[166] & b[124])^(a[165] & b[125])^(a[164] & b[126])^(a[163] & b[127])^(a[162] & b[128])^(a[161] & b[129])^(a[160] & b[130])^(a[159] & b[131])^(a[158] & b[132])^(a[157] & b[133])^(a[156] & b[134])^(a[155] & b[135])^(a[154] & b[136])^(a[153] & b[137])^(a[152] & b[138])^(a[151] & b[139])^(a[150] & b[140])^(a[149] & b[141])^(a[148] & b[142])^(a[147] & b[143])^(a[146] & b[144])^(a[145] & b[145])^(a[144] & b[146])^(a[143] & b[147])^(a[142] & b[148])^(a[141] & b[149])^(a[140] & b[150])^(a[139] & b[151])^(a[138] & b[152])^(a[137] & b[153])^(a[136] & b[154])^(a[135] & b[155])^(a[134] & b[156])^(a[133] & b[157])^(a[132] & b[158])^(a[131] & b[159])^(a[130] & b[160])^(a[129] & b[161])^(a[128] & b[162])^(a[127] & b[163])^(a[126] & b[164])^(a[125] & b[165])^(a[124] & b[166])^(a[123] & b[167])^(a[122] & b[168])^(a[121] & b[169])^(a[120] & b[170])^(a[119] & b[171])^(a[118] & b[172])^(a[117] & b[173])^(a[116] & b[174])^(a[115] & b[175])^(a[114] & b[176])^(a[113] & b[177])^(a[112] & b[178])^(a[111] & b[179])^(a[110] & b[180])^(a[109] & b[181])^(a[108] & b[182])^(a[107] & b[183])^(a[106] & b[184])^(a[105] & b[185])^(a[104] & b[186])^(a[103] & b[187])^(a[102] & b[188])^(a[101] & b[189])^(a[100] & b[190])^(a[99] & b[191])^(a[98] & b[192])^(a[97] & b[193])^(a[96] & b[194])^(a[95] & b[195])^(a[94] & b[196])^(a[93] & b[197])^(a[92] & b[198])^(a[91] & b[199])^(a[90] & b[200])^(a[89] & b[201])^(a[88] & b[202])^(a[87] & b[203])^(a[86] & b[204])^(a[85] & b[205])^(a[84] & b[206])^(a[83] & b[207])^(a[82] & b[208])^(a[81] & b[209])^(a[80] & b[210])^(a[79] & b[211])^(a[78] & b[212])^(a[77] & b[213])^(a[76] & b[214])^(a[75] & b[215])^(a[74] & b[216])^(a[73] & b[217])^(a[72] & b[218])^(a[71] & b[219])^(a[70] & b[220])^(a[69] & b[221])^(a[68] & b[222])^(a[67] & b[223])^(a[66] & b[224])^(a[65] & b[225])^(a[64] & b[226])^(a[63] & b[227])^(a[62] & b[228])^(a[61] & b[229])^(a[60] & b[230])^(a[59] & b[231])^(a[58] & b[232])^(a[57] & b[233])^(a[56] & b[234])^(a[55] & b[235])^(a[54] & b[236])^(a[53] & b[237])^(a[52] & b[238])^(a[51] & b[239])^(a[50] & b[240])^(a[49] & b[241])^(a[48] & b[242])^(a[47] & b[243])^(a[46] & b[244])^(a[45] & b[245])^(a[44] & b[246])^(a[43] & b[247])^(a[42] & b[248])^(a[41] & b[249])^(a[40] & b[250])^(a[39] & b[251])^(a[38] & b[252])^(a[37] & b[253])^(a[36] & b[254])^(a[35] & b[255])^(a[34] & b[256])^(a[33] & b[257])^(a[32] & b[258])^(a[31] & b[259])^(a[30] & b[260])^(a[29] & b[261])^(a[28] & b[262])^(a[27] & b[263])^(a[26] & b[264])^(a[25] & b[265])^(a[24] & b[266])^(a[23] & b[267])^(a[22] & b[268])^(a[21] & b[269])^(a[20] & b[270])^(a[19] & b[271])^(a[18] & b[272])^(a[17] & b[273])^(a[16] & b[274])^(a[15] & b[275])^(a[14] & b[276])^(a[13] & b[277])^(a[12] & b[278])^(a[11] & b[279])^(a[10] & b[280])^(a[9] & b[281])^(a[8] & b[282])^(a[7] & b[283])^(a[6] & b[284])^(a[5] & b[285])^(a[4] & b[286])^(a[3] & b[287])^(a[2] & b[288])^(a[1] & b[289])^(a[0] & b[290]);
assign y[291] = (a[291] & b[0])^(a[290] & b[1])^(a[289] & b[2])^(a[288] & b[3])^(a[287] & b[4])^(a[286] & b[5])^(a[285] & b[6])^(a[284] & b[7])^(a[283] & b[8])^(a[282] & b[9])^(a[281] & b[10])^(a[280] & b[11])^(a[279] & b[12])^(a[278] & b[13])^(a[277] & b[14])^(a[276] & b[15])^(a[275] & b[16])^(a[274] & b[17])^(a[273] & b[18])^(a[272] & b[19])^(a[271] & b[20])^(a[270] & b[21])^(a[269] & b[22])^(a[268] & b[23])^(a[267] & b[24])^(a[266] & b[25])^(a[265] & b[26])^(a[264] & b[27])^(a[263] & b[28])^(a[262] & b[29])^(a[261] & b[30])^(a[260] & b[31])^(a[259] & b[32])^(a[258] & b[33])^(a[257] & b[34])^(a[256] & b[35])^(a[255] & b[36])^(a[254] & b[37])^(a[253] & b[38])^(a[252] & b[39])^(a[251] & b[40])^(a[250] & b[41])^(a[249] & b[42])^(a[248] & b[43])^(a[247] & b[44])^(a[246] & b[45])^(a[245] & b[46])^(a[244] & b[47])^(a[243] & b[48])^(a[242] & b[49])^(a[241] & b[50])^(a[240] & b[51])^(a[239] & b[52])^(a[238] & b[53])^(a[237] & b[54])^(a[236] & b[55])^(a[235] & b[56])^(a[234] & b[57])^(a[233] & b[58])^(a[232] & b[59])^(a[231] & b[60])^(a[230] & b[61])^(a[229] & b[62])^(a[228] & b[63])^(a[227] & b[64])^(a[226] & b[65])^(a[225] & b[66])^(a[224] & b[67])^(a[223] & b[68])^(a[222] & b[69])^(a[221] & b[70])^(a[220] & b[71])^(a[219] & b[72])^(a[218] & b[73])^(a[217] & b[74])^(a[216] & b[75])^(a[215] & b[76])^(a[214] & b[77])^(a[213] & b[78])^(a[212] & b[79])^(a[211] & b[80])^(a[210] & b[81])^(a[209] & b[82])^(a[208] & b[83])^(a[207] & b[84])^(a[206] & b[85])^(a[205] & b[86])^(a[204] & b[87])^(a[203] & b[88])^(a[202] & b[89])^(a[201] & b[90])^(a[200] & b[91])^(a[199] & b[92])^(a[198] & b[93])^(a[197] & b[94])^(a[196] & b[95])^(a[195] & b[96])^(a[194] & b[97])^(a[193] & b[98])^(a[192] & b[99])^(a[191] & b[100])^(a[190] & b[101])^(a[189] & b[102])^(a[188] & b[103])^(a[187] & b[104])^(a[186] & b[105])^(a[185] & b[106])^(a[184] & b[107])^(a[183] & b[108])^(a[182] & b[109])^(a[181] & b[110])^(a[180] & b[111])^(a[179] & b[112])^(a[178] & b[113])^(a[177] & b[114])^(a[176] & b[115])^(a[175] & b[116])^(a[174] & b[117])^(a[173] & b[118])^(a[172] & b[119])^(a[171] & b[120])^(a[170] & b[121])^(a[169] & b[122])^(a[168] & b[123])^(a[167] & b[124])^(a[166] & b[125])^(a[165] & b[126])^(a[164] & b[127])^(a[163] & b[128])^(a[162] & b[129])^(a[161] & b[130])^(a[160] & b[131])^(a[159] & b[132])^(a[158] & b[133])^(a[157] & b[134])^(a[156] & b[135])^(a[155] & b[136])^(a[154] & b[137])^(a[153] & b[138])^(a[152] & b[139])^(a[151] & b[140])^(a[150] & b[141])^(a[149] & b[142])^(a[148] & b[143])^(a[147] & b[144])^(a[146] & b[145])^(a[145] & b[146])^(a[144] & b[147])^(a[143] & b[148])^(a[142] & b[149])^(a[141] & b[150])^(a[140] & b[151])^(a[139] & b[152])^(a[138] & b[153])^(a[137] & b[154])^(a[136] & b[155])^(a[135] & b[156])^(a[134] & b[157])^(a[133] & b[158])^(a[132] & b[159])^(a[131] & b[160])^(a[130] & b[161])^(a[129] & b[162])^(a[128] & b[163])^(a[127] & b[164])^(a[126] & b[165])^(a[125] & b[166])^(a[124] & b[167])^(a[123] & b[168])^(a[122] & b[169])^(a[121] & b[170])^(a[120] & b[171])^(a[119] & b[172])^(a[118] & b[173])^(a[117] & b[174])^(a[116] & b[175])^(a[115] & b[176])^(a[114] & b[177])^(a[113] & b[178])^(a[112] & b[179])^(a[111] & b[180])^(a[110] & b[181])^(a[109] & b[182])^(a[108] & b[183])^(a[107] & b[184])^(a[106] & b[185])^(a[105] & b[186])^(a[104] & b[187])^(a[103] & b[188])^(a[102] & b[189])^(a[101] & b[190])^(a[100] & b[191])^(a[99] & b[192])^(a[98] & b[193])^(a[97] & b[194])^(a[96] & b[195])^(a[95] & b[196])^(a[94] & b[197])^(a[93] & b[198])^(a[92] & b[199])^(a[91] & b[200])^(a[90] & b[201])^(a[89] & b[202])^(a[88] & b[203])^(a[87] & b[204])^(a[86] & b[205])^(a[85] & b[206])^(a[84] & b[207])^(a[83] & b[208])^(a[82] & b[209])^(a[81] & b[210])^(a[80] & b[211])^(a[79] & b[212])^(a[78] & b[213])^(a[77] & b[214])^(a[76] & b[215])^(a[75] & b[216])^(a[74] & b[217])^(a[73] & b[218])^(a[72] & b[219])^(a[71] & b[220])^(a[70] & b[221])^(a[69] & b[222])^(a[68] & b[223])^(a[67] & b[224])^(a[66] & b[225])^(a[65] & b[226])^(a[64] & b[227])^(a[63] & b[228])^(a[62] & b[229])^(a[61] & b[230])^(a[60] & b[231])^(a[59] & b[232])^(a[58] & b[233])^(a[57] & b[234])^(a[56] & b[235])^(a[55] & b[236])^(a[54] & b[237])^(a[53] & b[238])^(a[52] & b[239])^(a[51] & b[240])^(a[50] & b[241])^(a[49] & b[242])^(a[48] & b[243])^(a[47] & b[244])^(a[46] & b[245])^(a[45] & b[246])^(a[44] & b[247])^(a[43] & b[248])^(a[42] & b[249])^(a[41] & b[250])^(a[40] & b[251])^(a[39] & b[252])^(a[38] & b[253])^(a[37] & b[254])^(a[36] & b[255])^(a[35] & b[256])^(a[34] & b[257])^(a[33] & b[258])^(a[32] & b[259])^(a[31] & b[260])^(a[30] & b[261])^(a[29] & b[262])^(a[28] & b[263])^(a[27] & b[264])^(a[26] & b[265])^(a[25] & b[266])^(a[24] & b[267])^(a[23] & b[268])^(a[22] & b[269])^(a[21] & b[270])^(a[20] & b[271])^(a[19] & b[272])^(a[18] & b[273])^(a[17] & b[274])^(a[16] & b[275])^(a[15] & b[276])^(a[14] & b[277])^(a[13] & b[278])^(a[12] & b[279])^(a[11] & b[280])^(a[10] & b[281])^(a[9] & b[282])^(a[8] & b[283])^(a[7] & b[284])^(a[6] & b[285])^(a[5] & b[286])^(a[4] & b[287])^(a[3] & b[288])^(a[2] & b[289])^(a[1] & b[290])^(a[0] & b[291]);
assign y[292] = (a[292] & b[0])^(a[291] & b[1])^(a[290] & b[2])^(a[289] & b[3])^(a[288] & b[4])^(a[287] & b[5])^(a[286] & b[6])^(a[285] & b[7])^(a[284] & b[8])^(a[283] & b[9])^(a[282] & b[10])^(a[281] & b[11])^(a[280] & b[12])^(a[279] & b[13])^(a[278] & b[14])^(a[277] & b[15])^(a[276] & b[16])^(a[275] & b[17])^(a[274] & b[18])^(a[273] & b[19])^(a[272] & b[20])^(a[271] & b[21])^(a[270] & b[22])^(a[269] & b[23])^(a[268] & b[24])^(a[267] & b[25])^(a[266] & b[26])^(a[265] & b[27])^(a[264] & b[28])^(a[263] & b[29])^(a[262] & b[30])^(a[261] & b[31])^(a[260] & b[32])^(a[259] & b[33])^(a[258] & b[34])^(a[257] & b[35])^(a[256] & b[36])^(a[255] & b[37])^(a[254] & b[38])^(a[253] & b[39])^(a[252] & b[40])^(a[251] & b[41])^(a[250] & b[42])^(a[249] & b[43])^(a[248] & b[44])^(a[247] & b[45])^(a[246] & b[46])^(a[245] & b[47])^(a[244] & b[48])^(a[243] & b[49])^(a[242] & b[50])^(a[241] & b[51])^(a[240] & b[52])^(a[239] & b[53])^(a[238] & b[54])^(a[237] & b[55])^(a[236] & b[56])^(a[235] & b[57])^(a[234] & b[58])^(a[233] & b[59])^(a[232] & b[60])^(a[231] & b[61])^(a[230] & b[62])^(a[229] & b[63])^(a[228] & b[64])^(a[227] & b[65])^(a[226] & b[66])^(a[225] & b[67])^(a[224] & b[68])^(a[223] & b[69])^(a[222] & b[70])^(a[221] & b[71])^(a[220] & b[72])^(a[219] & b[73])^(a[218] & b[74])^(a[217] & b[75])^(a[216] & b[76])^(a[215] & b[77])^(a[214] & b[78])^(a[213] & b[79])^(a[212] & b[80])^(a[211] & b[81])^(a[210] & b[82])^(a[209] & b[83])^(a[208] & b[84])^(a[207] & b[85])^(a[206] & b[86])^(a[205] & b[87])^(a[204] & b[88])^(a[203] & b[89])^(a[202] & b[90])^(a[201] & b[91])^(a[200] & b[92])^(a[199] & b[93])^(a[198] & b[94])^(a[197] & b[95])^(a[196] & b[96])^(a[195] & b[97])^(a[194] & b[98])^(a[193] & b[99])^(a[192] & b[100])^(a[191] & b[101])^(a[190] & b[102])^(a[189] & b[103])^(a[188] & b[104])^(a[187] & b[105])^(a[186] & b[106])^(a[185] & b[107])^(a[184] & b[108])^(a[183] & b[109])^(a[182] & b[110])^(a[181] & b[111])^(a[180] & b[112])^(a[179] & b[113])^(a[178] & b[114])^(a[177] & b[115])^(a[176] & b[116])^(a[175] & b[117])^(a[174] & b[118])^(a[173] & b[119])^(a[172] & b[120])^(a[171] & b[121])^(a[170] & b[122])^(a[169] & b[123])^(a[168] & b[124])^(a[167] & b[125])^(a[166] & b[126])^(a[165] & b[127])^(a[164] & b[128])^(a[163] & b[129])^(a[162] & b[130])^(a[161] & b[131])^(a[160] & b[132])^(a[159] & b[133])^(a[158] & b[134])^(a[157] & b[135])^(a[156] & b[136])^(a[155] & b[137])^(a[154] & b[138])^(a[153] & b[139])^(a[152] & b[140])^(a[151] & b[141])^(a[150] & b[142])^(a[149] & b[143])^(a[148] & b[144])^(a[147] & b[145])^(a[146] & b[146])^(a[145] & b[147])^(a[144] & b[148])^(a[143] & b[149])^(a[142] & b[150])^(a[141] & b[151])^(a[140] & b[152])^(a[139] & b[153])^(a[138] & b[154])^(a[137] & b[155])^(a[136] & b[156])^(a[135] & b[157])^(a[134] & b[158])^(a[133] & b[159])^(a[132] & b[160])^(a[131] & b[161])^(a[130] & b[162])^(a[129] & b[163])^(a[128] & b[164])^(a[127] & b[165])^(a[126] & b[166])^(a[125] & b[167])^(a[124] & b[168])^(a[123] & b[169])^(a[122] & b[170])^(a[121] & b[171])^(a[120] & b[172])^(a[119] & b[173])^(a[118] & b[174])^(a[117] & b[175])^(a[116] & b[176])^(a[115] & b[177])^(a[114] & b[178])^(a[113] & b[179])^(a[112] & b[180])^(a[111] & b[181])^(a[110] & b[182])^(a[109] & b[183])^(a[108] & b[184])^(a[107] & b[185])^(a[106] & b[186])^(a[105] & b[187])^(a[104] & b[188])^(a[103] & b[189])^(a[102] & b[190])^(a[101] & b[191])^(a[100] & b[192])^(a[99] & b[193])^(a[98] & b[194])^(a[97] & b[195])^(a[96] & b[196])^(a[95] & b[197])^(a[94] & b[198])^(a[93] & b[199])^(a[92] & b[200])^(a[91] & b[201])^(a[90] & b[202])^(a[89] & b[203])^(a[88] & b[204])^(a[87] & b[205])^(a[86] & b[206])^(a[85] & b[207])^(a[84] & b[208])^(a[83] & b[209])^(a[82] & b[210])^(a[81] & b[211])^(a[80] & b[212])^(a[79] & b[213])^(a[78] & b[214])^(a[77] & b[215])^(a[76] & b[216])^(a[75] & b[217])^(a[74] & b[218])^(a[73] & b[219])^(a[72] & b[220])^(a[71] & b[221])^(a[70] & b[222])^(a[69] & b[223])^(a[68] & b[224])^(a[67] & b[225])^(a[66] & b[226])^(a[65] & b[227])^(a[64] & b[228])^(a[63] & b[229])^(a[62] & b[230])^(a[61] & b[231])^(a[60] & b[232])^(a[59] & b[233])^(a[58] & b[234])^(a[57] & b[235])^(a[56] & b[236])^(a[55] & b[237])^(a[54] & b[238])^(a[53] & b[239])^(a[52] & b[240])^(a[51] & b[241])^(a[50] & b[242])^(a[49] & b[243])^(a[48] & b[244])^(a[47] & b[245])^(a[46] & b[246])^(a[45] & b[247])^(a[44] & b[248])^(a[43] & b[249])^(a[42] & b[250])^(a[41] & b[251])^(a[40] & b[252])^(a[39] & b[253])^(a[38] & b[254])^(a[37] & b[255])^(a[36] & b[256])^(a[35] & b[257])^(a[34] & b[258])^(a[33] & b[259])^(a[32] & b[260])^(a[31] & b[261])^(a[30] & b[262])^(a[29] & b[263])^(a[28] & b[264])^(a[27] & b[265])^(a[26] & b[266])^(a[25] & b[267])^(a[24] & b[268])^(a[23] & b[269])^(a[22] & b[270])^(a[21] & b[271])^(a[20] & b[272])^(a[19] & b[273])^(a[18] & b[274])^(a[17] & b[275])^(a[16] & b[276])^(a[15] & b[277])^(a[14] & b[278])^(a[13] & b[279])^(a[12] & b[280])^(a[11] & b[281])^(a[10] & b[282])^(a[9] & b[283])^(a[8] & b[284])^(a[7] & b[285])^(a[6] & b[286])^(a[5] & b[287])^(a[4] & b[288])^(a[3] & b[289])^(a[2] & b[290])^(a[1] & b[291])^(a[0] & b[292]);
assign y[293] = (a[293] & b[0])^(a[292] & b[1])^(a[291] & b[2])^(a[290] & b[3])^(a[289] & b[4])^(a[288] & b[5])^(a[287] & b[6])^(a[286] & b[7])^(a[285] & b[8])^(a[284] & b[9])^(a[283] & b[10])^(a[282] & b[11])^(a[281] & b[12])^(a[280] & b[13])^(a[279] & b[14])^(a[278] & b[15])^(a[277] & b[16])^(a[276] & b[17])^(a[275] & b[18])^(a[274] & b[19])^(a[273] & b[20])^(a[272] & b[21])^(a[271] & b[22])^(a[270] & b[23])^(a[269] & b[24])^(a[268] & b[25])^(a[267] & b[26])^(a[266] & b[27])^(a[265] & b[28])^(a[264] & b[29])^(a[263] & b[30])^(a[262] & b[31])^(a[261] & b[32])^(a[260] & b[33])^(a[259] & b[34])^(a[258] & b[35])^(a[257] & b[36])^(a[256] & b[37])^(a[255] & b[38])^(a[254] & b[39])^(a[253] & b[40])^(a[252] & b[41])^(a[251] & b[42])^(a[250] & b[43])^(a[249] & b[44])^(a[248] & b[45])^(a[247] & b[46])^(a[246] & b[47])^(a[245] & b[48])^(a[244] & b[49])^(a[243] & b[50])^(a[242] & b[51])^(a[241] & b[52])^(a[240] & b[53])^(a[239] & b[54])^(a[238] & b[55])^(a[237] & b[56])^(a[236] & b[57])^(a[235] & b[58])^(a[234] & b[59])^(a[233] & b[60])^(a[232] & b[61])^(a[231] & b[62])^(a[230] & b[63])^(a[229] & b[64])^(a[228] & b[65])^(a[227] & b[66])^(a[226] & b[67])^(a[225] & b[68])^(a[224] & b[69])^(a[223] & b[70])^(a[222] & b[71])^(a[221] & b[72])^(a[220] & b[73])^(a[219] & b[74])^(a[218] & b[75])^(a[217] & b[76])^(a[216] & b[77])^(a[215] & b[78])^(a[214] & b[79])^(a[213] & b[80])^(a[212] & b[81])^(a[211] & b[82])^(a[210] & b[83])^(a[209] & b[84])^(a[208] & b[85])^(a[207] & b[86])^(a[206] & b[87])^(a[205] & b[88])^(a[204] & b[89])^(a[203] & b[90])^(a[202] & b[91])^(a[201] & b[92])^(a[200] & b[93])^(a[199] & b[94])^(a[198] & b[95])^(a[197] & b[96])^(a[196] & b[97])^(a[195] & b[98])^(a[194] & b[99])^(a[193] & b[100])^(a[192] & b[101])^(a[191] & b[102])^(a[190] & b[103])^(a[189] & b[104])^(a[188] & b[105])^(a[187] & b[106])^(a[186] & b[107])^(a[185] & b[108])^(a[184] & b[109])^(a[183] & b[110])^(a[182] & b[111])^(a[181] & b[112])^(a[180] & b[113])^(a[179] & b[114])^(a[178] & b[115])^(a[177] & b[116])^(a[176] & b[117])^(a[175] & b[118])^(a[174] & b[119])^(a[173] & b[120])^(a[172] & b[121])^(a[171] & b[122])^(a[170] & b[123])^(a[169] & b[124])^(a[168] & b[125])^(a[167] & b[126])^(a[166] & b[127])^(a[165] & b[128])^(a[164] & b[129])^(a[163] & b[130])^(a[162] & b[131])^(a[161] & b[132])^(a[160] & b[133])^(a[159] & b[134])^(a[158] & b[135])^(a[157] & b[136])^(a[156] & b[137])^(a[155] & b[138])^(a[154] & b[139])^(a[153] & b[140])^(a[152] & b[141])^(a[151] & b[142])^(a[150] & b[143])^(a[149] & b[144])^(a[148] & b[145])^(a[147] & b[146])^(a[146] & b[147])^(a[145] & b[148])^(a[144] & b[149])^(a[143] & b[150])^(a[142] & b[151])^(a[141] & b[152])^(a[140] & b[153])^(a[139] & b[154])^(a[138] & b[155])^(a[137] & b[156])^(a[136] & b[157])^(a[135] & b[158])^(a[134] & b[159])^(a[133] & b[160])^(a[132] & b[161])^(a[131] & b[162])^(a[130] & b[163])^(a[129] & b[164])^(a[128] & b[165])^(a[127] & b[166])^(a[126] & b[167])^(a[125] & b[168])^(a[124] & b[169])^(a[123] & b[170])^(a[122] & b[171])^(a[121] & b[172])^(a[120] & b[173])^(a[119] & b[174])^(a[118] & b[175])^(a[117] & b[176])^(a[116] & b[177])^(a[115] & b[178])^(a[114] & b[179])^(a[113] & b[180])^(a[112] & b[181])^(a[111] & b[182])^(a[110] & b[183])^(a[109] & b[184])^(a[108] & b[185])^(a[107] & b[186])^(a[106] & b[187])^(a[105] & b[188])^(a[104] & b[189])^(a[103] & b[190])^(a[102] & b[191])^(a[101] & b[192])^(a[100] & b[193])^(a[99] & b[194])^(a[98] & b[195])^(a[97] & b[196])^(a[96] & b[197])^(a[95] & b[198])^(a[94] & b[199])^(a[93] & b[200])^(a[92] & b[201])^(a[91] & b[202])^(a[90] & b[203])^(a[89] & b[204])^(a[88] & b[205])^(a[87] & b[206])^(a[86] & b[207])^(a[85] & b[208])^(a[84] & b[209])^(a[83] & b[210])^(a[82] & b[211])^(a[81] & b[212])^(a[80] & b[213])^(a[79] & b[214])^(a[78] & b[215])^(a[77] & b[216])^(a[76] & b[217])^(a[75] & b[218])^(a[74] & b[219])^(a[73] & b[220])^(a[72] & b[221])^(a[71] & b[222])^(a[70] & b[223])^(a[69] & b[224])^(a[68] & b[225])^(a[67] & b[226])^(a[66] & b[227])^(a[65] & b[228])^(a[64] & b[229])^(a[63] & b[230])^(a[62] & b[231])^(a[61] & b[232])^(a[60] & b[233])^(a[59] & b[234])^(a[58] & b[235])^(a[57] & b[236])^(a[56] & b[237])^(a[55] & b[238])^(a[54] & b[239])^(a[53] & b[240])^(a[52] & b[241])^(a[51] & b[242])^(a[50] & b[243])^(a[49] & b[244])^(a[48] & b[245])^(a[47] & b[246])^(a[46] & b[247])^(a[45] & b[248])^(a[44] & b[249])^(a[43] & b[250])^(a[42] & b[251])^(a[41] & b[252])^(a[40] & b[253])^(a[39] & b[254])^(a[38] & b[255])^(a[37] & b[256])^(a[36] & b[257])^(a[35] & b[258])^(a[34] & b[259])^(a[33] & b[260])^(a[32] & b[261])^(a[31] & b[262])^(a[30] & b[263])^(a[29] & b[264])^(a[28] & b[265])^(a[27] & b[266])^(a[26] & b[267])^(a[25] & b[268])^(a[24] & b[269])^(a[23] & b[270])^(a[22] & b[271])^(a[21] & b[272])^(a[20] & b[273])^(a[19] & b[274])^(a[18] & b[275])^(a[17] & b[276])^(a[16] & b[277])^(a[15] & b[278])^(a[14] & b[279])^(a[13] & b[280])^(a[12] & b[281])^(a[11] & b[282])^(a[10] & b[283])^(a[9] & b[284])^(a[8] & b[285])^(a[7] & b[286])^(a[6] & b[287])^(a[5] & b[288])^(a[4] & b[289])^(a[3] & b[290])^(a[2] & b[291])^(a[1] & b[292])^(a[0] & b[293]);
assign y[294] = (a[294] & b[0])^(a[293] & b[1])^(a[292] & b[2])^(a[291] & b[3])^(a[290] & b[4])^(a[289] & b[5])^(a[288] & b[6])^(a[287] & b[7])^(a[286] & b[8])^(a[285] & b[9])^(a[284] & b[10])^(a[283] & b[11])^(a[282] & b[12])^(a[281] & b[13])^(a[280] & b[14])^(a[279] & b[15])^(a[278] & b[16])^(a[277] & b[17])^(a[276] & b[18])^(a[275] & b[19])^(a[274] & b[20])^(a[273] & b[21])^(a[272] & b[22])^(a[271] & b[23])^(a[270] & b[24])^(a[269] & b[25])^(a[268] & b[26])^(a[267] & b[27])^(a[266] & b[28])^(a[265] & b[29])^(a[264] & b[30])^(a[263] & b[31])^(a[262] & b[32])^(a[261] & b[33])^(a[260] & b[34])^(a[259] & b[35])^(a[258] & b[36])^(a[257] & b[37])^(a[256] & b[38])^(a[255] & b[39])^(a[254] & b[40])^(a[253] & b[41])^(a[252] & b[42])^(a[251] & b[43])^(a[250] & b[44])^(a[249] & b[45])^(a[248] & b[46])^(a[247] & b[47])^(a[246] & b[48])^(a[245] & b[49])^(a[244] & b[50])^(a[243] & b[51])^(a[242] & b[52])^(a[241] & b[53])^(a[240] & b[54])^(a[239] & b[55])^(a[238] & b[56])^(a[237] & b[57])^(a[236] & b[58])^(a[235] & b[59])^(a[234] & b[60])^(a[233] & b[61])^(a[232] & b[62])^(a[231] & b[63])^(a[230] & b[64])^(a[229] & b[65])^(a[228] & b[66])^(a[227] & b[67])^(a[226] & b[68])^(a[225] & b[69])^(a[224] & b[70])^(a[223] & b[71])^(a[222] & b[72])^(a[221] & b[73])^(a[220] & b[74])^(a[219] & b[75])^(a[218] & b[76])^(a[217] & b[77])^(a[216] & b[78])^(a[215] & b[79])^(a[214] & b[80])^(a[213] & b[81])^(a[212] & b[82])^(a[211] & b[83])^(a[210] & b[84])^(a[209] & b[85])^(a[208] & b[86])^(a[207] & b[87])^(a[206] & b[88])^(a[205] & b[89])^(a[204] & b[90])^(a[203] & b[91])^(a[202] & b[92])^(a[201] & b[93])^(a[200] & b[94])^(a[199] & b[95])^(a[198] & b[96])^(a[197] & b[97])^(a[196] & b[98])^(a[195] & b[99])^(a[194] & b[100])^(a[193] & b[101])^(a[192] & b[102])^(a[191] & b[103])^(a[190] & b[104])^(a[189] & b[105])^(a[188] & b[106])^(a[187] & b[107])^(a[186] & b[108])^(a[185] & b[109])^(a[184] & b[110])^(a[183] & b[111])^(a[182] & b[112])^(a[181] & b[113])^(a[180] & b[114])^(a[179] & b[115])^(a[178] & b[116])^(a[177] & b[117])^(a[176] & b[118])^(a[175] & b[119])^(a[174] & b[120])^(a[173] & b[121])^(a[172] & b[122])^(a[171] & b[123])^(a[170] & b[124])^(a[169] & b[125])^(a[168] & b[126])^(a[167] & b[127])^(a[166] & b[128])^(a[165] & b[129])^(a[164] & b[130])^(a[163] & b[131])^(a[162] & b[132])^(a[161] & b[133])^(a[160] & b[134])^(a[159] & b[135])^(a[158] & b[136])^(a[157] & b[137])^(a[156] & b[138])^(a[155] & b[139])^(a[154] & b[140])^(a[153] & b[141])^(a[152] & b[142])^(a[151] & b[143])^(a[150] & b[144])^(a[149] & b[145])^(a[148] & b[146])^(a[147] & b[147])^(a[146] & b[148])^(a[145] & b[149])^(a[144] & b[150])^(a[143] & b[151])^(a[142] & b[152])^(a[141] & b[153])^(a[140] & b[154])^(a[139] & b[155])^(a[138] & b[156])^(a[137] & b[157])^(a[136] & b[158])^(a[135] & b[159])^(a[134] & b[160])^(a[133] & b[161])^(a[132] & b[162])^(a[131] & b[163])^(a[130] & b[164])^(a[129] & b[165])^(a[128] & b[166])^(a[127] & b[167])^(a[126] & b[168])^(a[125] & b[169])^(a[124] & b[170])^(a[123] & b[171])^(a[122] & b[172])^(a[121] & b[173])^(a[120] & b[174])^(a[119] & b[175])^(a[118] & b[176])^(a[117] & b[177])^(a[116] & b[178])^(a[115] & b[179])^(a[114] & b[180])^(a[113] & b[181])^(a[112] & b[182])^(a[111] & b[183])^(a[110] & b[184])^(a[109] & b[185])^(a[108] & b[186])^(a[107] & b[187])^(a[106] & b[188])^(a[105] & b[189])^(a[104] & b[190])^(a[103] & b[191])^(a[102] & b[192])^(a[101] & b[193])^(a[100] & b[194])^(a[99] & b[195])^(a[98] & b[196])^(a[97] & b[197])^(a[96] & b[198])^(a[95] & b[199])^(a[94] & b[200])^(a[93] & b[201])^(a[92] & b[202])^(a[91] & b[203])^(a[90] & b[204])^(a[89] & b[205])^(a[88] & b[206])^(a[87] & b[207])^(a[86] & b[208])^(a[85] & b[209])^(a[84] & b[210])^(a[83] & b[211])^(a[82] & b[212])^(a[81] & b[213])^(a[80] & b[214])^(a[79] & b[215])^(a[78] & b[216])^(a[77] & b[217])^(a[76] & b[218])^(a[75] & b[219])^(a[74] & b[220])^(a[73] & b[221])^(a[72] & b[222])^(a[71] & b[223])^(a[70] & b[224])^(a[69] & b[225])^(a[68] & b[226])^(a[67] & b[227])^(a[66] & b[228])^(a[65] & b[229])^(a[64] & b[230])^(a[63] & b[231])^(a[62] & b[232])^(a[61] & b[233])^(a[60] & b[234])^(a[59] & b[235])^(a[58] & b[236])^(a[57] & b[237])^(a[56] & b[238])^(a[55] & b[239])^(a[54] & b[240])^(a[53] & b[241])^(a[52] & b[242])^(a[51] & b[243])^(a[50] & b[244])^(a[49] & b[245])^(a[48] & b[246])^(a[47] & b[247])^(a[46] & b[248])^(a[45] & b[249])^(a[44] & b[250])^(a[43] & b[251])^(a[42] & b[252])^(a[41] & b[253])^(a[40] & b[254])^(a[39] & b[255])^(a[38] & b[256])^(a[37] & b[257])^(a[36] & b[258])^(a[35] & b[259])^(a[34] & b[260])^(a[33] & b[261])^(a[32] & b[262])^(a[31] & b[263])^(a[30] & b[264])^(a[29] & b[265])^(a[28] & b[266])^(a[27] & b[267])^(a[26] & b[268])^(a[25] & b[269])^(a[24] & b[270])^(a[23] & b[271])^(a[22] & b[272])^(a[21] & b[273])^(a[20] & b[274])^(a[19] & b[275])^(a[18] & b[276])^(a[17] & b[277])^(a[16] & b[278])^(a[15] & b[279])^(a[14] & b[280])^(a[13] & b[281])^(a[12] & b[282])^(a[11] & b[283])^(a[10] & b[284])^(a[9] & b[285])^(a[8] & b[286])^(a[7] & b[287])^(a[6] & b[288])^(a[5] & b[289])^(a[4] & b[290])^(a[3] & b[291])^(a[2] & b[292])^(a[1] & b[293])^(a[0] & b[294]);
assign y[295] = (a[295] & b[0])^(a[294] & b[1])^(a[293] & b[2])^(a[292] & b[3])^(a[291] & b[4])^(a[290] & b[5])^(a[289] & b[6])^(a[288] & b[7])^(a[287] & b[8])^(a[286] & b[9])^(a[285] & b[10])^(a[284] & b[11])^(a[283] & b[12])^(a[282] & b[13])^(a[281] & b[14])^(a[280] & b[15])^(a[279] & b[16])^(a[278] & b[17])^(a[277] & b[18])^(a[276] & b[19])^(a[275] & b[20])^(a[274] & b[21])^(a[273] & b[22])^(a[272] & b[23])^(a[271] & b[24])^(a[270] & b[25])^(a[269] & b[26])^(a[268] & b[27])^(a[267] & b[28])^(a[266] & b[29])^(a[265] & b[30])^(a[264] & b[31])^(a[263] & b[32])^(a[262] & b[33])^(a[261] & b[34])^(a[260] & b[35])^(a[259] & b[36])^(a[258] & b[37])^(a[257] & b[38])^(a[256] & b[39])^(a[255] & b[40])^(a[254] & b[41])^(a[253] & b[42])^(a[252] & b[43])^(a[251] & b[44])^(a[250] & b[45])^(a[249] & b[46])^(a[248] & b[47])^(a[247] & b[48])^(a[246] & b[49])^(a[245] & b[50])^(a[244] & b[51])^(a[243] & b[52])^(a[242] & b[53])^(a[241] & b[54])^(a[240] & b[55])^(a[239] & b[56])^(a[238] & b[57])^(a[237] & b[58])^(a[236] & b[59])^(a[235] & b[60])^(a[234] & b[61])^(a[233] & b[62])^(a[232] & b[63])^(a[231] & b[64])^(a[230] & b[65])^(a[229] & b[66])^(a[228] & b[67])^(a[227] & b[68])^(a[226] & b[69])^(a[225] & b[70])^(a[224] & b[71])^(a[223] & b[72])^(a[222] & b[73])^(a[221] & b[74])^(a[220] & b[75])^(a[219] & b[76])^(a[218] & b[77])^(a[217] & b[78])^(a[216] & b[79])^(a[215] & b[80])^(a[214] & b[81])^(a[213] & b[82])^(a[212] & b[83])^(a[211] & b[84])^(a[210] & b[85])^(a[209] & b[86])^(a[208] & b[87])^(a[207] & b[88])^(a[206] & b[89])^(a[205] & b[90])^(a[204] & b[91])^(a[203] & b[92])^(a[202] & b[93])^(a[201] & b[94])^(a[200] & b[95])^(a[199] & b[96])^(a[198] & b[97])^(a[197] & b[98])^(a[196] & b[99])^(a[195] & b[100])^(a[194] & b[101])^(a[193] & b[102])^(a[192] & b[103])^(a[191] & b[104])^(a[190] & b[105])^(a[189] & b[106])^(a[188] & b[107])^(a[187] & b[108])^(a[186] & b[109])^(a[185] & b[110])^(a[184] & b[111])^(a[183] & b[112])^(a[182] & b[113])^(a[181] & b[114])^(a[180] & b[115])^(a[179] & b[116])^(a[178] & b[117])^(a[177] & b[118])^(a[176] & b[119])^(a[175] & b[120])^(a[174] & b[121])^(a[173] & b[122])^(a[172] & b[123])^(a[171] & b[124])^(a[170] & b[125])^(a[169] & b[126])^(a[168] & b[127])^(a[167] & b[128])^(a[166] & b[129])^(a[165] & b[130])^(a[164] & b[131])^(a[163] & b[132])^(a[162] & b[133])^(a[161] & b[134])^(a[160] & b[135])^(a[159] & b[136])^(a[158] & b[137])^(a[157] & b[138])^(a[156] & b[139])^(a[155] & b[140])^(a[154] & b[141])^(a[153] & b[142])^(a[152] & b[143])^(a[151] & b[144])^(a[150] & b[145])^(a[149] & b[146])^(a[148] & b[147])^(a[147] & b[148])^(a[146] & b[149])^(a[145] & b[150])^(a[144] & b[151])^(a[143] & b[152])^(a[142] & b[153])^(a[141] & b[154])^(a[140] & b[155])^(a[139] & b[156])^(a[138] & b[157])^(a[137] & b[158])^(a[136] & b[159])^(a[135] & b[160])^(a[134] & b[161])^(a[133] & b[162])^(a[132] & b[163])^(a[131] & b[164])^(a[130] & b[165])^(a[129] & b[166])^(a[128] & b[167])^(a[127] & b[168])^(a[126] & b[169])^(a[125] & b[170])^(a[124] & b[171])^(a[123] & b[172])^(a[122] & b[173])^(a[121] & b[174])^(a[120] & b[175])^(a[119] & b[176])^(a[118] & b[177])^(a[117] & b[178])^(a[116] & b[179])^(a[115] & b[180])^(a[114] & b[181])^(a[113] & b[182])^(a[112] & b[183])^(a[111] & b[184])^(a[110] & b[185])^(a[109] & b[186])^(a[108] & b[187])^(a[107] & b[188])^(a[106] & b[189])^(a[105] & b[190])^(a[104] & b[191])^(a[103] & b[192])^(a[102] & b[193])^(a[101] & b[194])^(a[100] & b[195])^(a[99] & b[196])^(a[98] & b[197])^(a[97] & b[198])^(a[96] & b[199])^(a[95] & b[200])^(a[94] & b[201])^(a[93] & b[202])^(a[92] & b[203])^(a[91] & b[204])^(a[90] & b[205])^(a[89] & b[206])^(a[88] & b[207])^(a[87] & b[208])^(a[86] & b[209])^(a[85] & b[210])^(a[84] & b[211])^(a[83] & b[212])^(a[82] & b[213])^(a[81] & b[214])^(a[80] & b[215])^(a[79] & b[216])^(a[78] & b[217])^(a[77] & b[218])^(a[76] & b[219])^(a[75] & b[220])^(a[74] & b[221])^(a[73] & b[222])^(a[72] & b[223])^(a[71] & b[224])^(a[70] & b[225])^(a[69] & b[226])^(a[68] & b[227])^(a[67] & b[228])^(a[66] & b[229])^(a[65] & b[230])^(a[64] & b[231])^(a[63] & b[232])^(a[62] & b[233])^(a[61] & b[234])^(a[60] & b[235])^(a[59] & b[236])^(a[58] & b[237])^(a[57] & b[238])^(a[56] & b[239])^(a[55] & b[240])^(a[54] & b[241])^(a[53] & b[242])^(a[52] & b[243])^(a[51] & b[244])^(a[50] & b[245])^(a[49] & b[246])^(a[48] & b[247])^(a[47] & b[248])^(a[46] & b[249])^(a[45] & b[250])^(a[44] & b[251])^(a[43] & b[252])^(a[42] & b[253])^(a[41] & b[254])^(a[40] & b[255])^(a[39] & b[256])^(a[38] & b[257])^(a[37] & b[258])^(a[36] & b[259])^(a[35] & b[260])^(a[34] & b[261])^(a[33] & b[262])^(a[32] & b[263])^(a[31] & b[264])^(a[30] & b[265])^(a[29] & b[266])^(a[28] & b[267])^(a[27] & b[268])^(a[26] & b[269])^(a[25] & b[270])^(a[24] & b[271])^(a[23] & b[272])^(a[22] & b[273])^(a[21] & b[274])^(a[20] & b[275])^(a[19] & b[276])^(a[18] & b[277])^(a[17] & b[278])^(a[16] & b[279])^(a[15] & b[280])^(a[14] & b[281])^(a[13] & b[282])^(a[12] & b[283])^(a[11] & b[284])^(a[10] & b[285])^(a[9] & b[286])^(a[8] & b[287])^(a[7] & b[288])^(a[6] & b[289])^(a[5] & b[290])^(a[4] & b[291])^(a[3] & b[292])^(a[2] & b[293])^(a[1] & b[294])^(a[0] & b[295]);
assign y[296] = (a[296] & b[0])^(a[295] & b[1])^(a[294] & b[2])^(a[293] & b[3])^(a[292] & b[4])^(a[291] & b[5])^(a[290] & b[6])^(a[289] & b[7])^(a[288] & b[8])^(a[287] & b[9])^(a[286] & b[10])^(a[285] & b[11])^(a[284] & b[12])^(a[283] & b[13])^(a[282] & b[14])^(a[281] & b[15])^(a[280] & b[16])^(a[279] & b[17])^(a[278] & b[18])^(a[277] & b[19])^(a[276] & b[20])^(a[275] & b[21])^(a[274] & b[22])^(a[273] & b[23])^(a[272] & b[24])^(a[271] & b[25])^(a[270] & b[26])^(a[269] & b[27])^(a[268] & b[28])^(a[267] & b[29])^(a[266] & b[30])^(a[265] & b[31])^(a[264] & b[32])^(a[263] & b[33])^(a[262] & b[34])^(a[261] & b[35])^(a[260] & b[36])^(a[259] & b[37])^(a[258] & b[38])^(a[257] & b[39])^(a[256] & b[40])^(a[255] & b[41])^(a[254] & b[42])^(a[253] & b[43])^(a[252] & b[44])^(a[251] & b[45])^(a[250] & b[46])^(a[249] & b[47])^(a[248] & b[48])^(a[247] & b[49])^(a[246] & b[50])^(a[245] & b[51])^(a[244] & b[52])^(a[243] & b[53])^(a[242] & b[54])^(a[241] & b[55])^(a[240] & b[56])^(a[239] & b[57])^(a[238] & b[58])^(a[237] & b[59])^(a[236] & b[60])^(a[235] & b[61])^(a[234] & b[62])^(a[233] & b[63])^(a[232] & b[64])^(a[231] & b[65])^(a[230] & b[66])^(a[229] & b[67])^(a[228] & b[68])^(a[227] & b[69])^(a[226] & b[70])^(a[225] & b[71])^(a[224] & b[72])^(a[223] & b[73])^(a[222] & b[74])^(a[221] & b[75])^(a[220] & b[76])^(a[219] & b[77])^(a[218] & b[78])^(a[217] & b[79])^(a[216] & b[80])^(a[215] & b[81])^(a[214] & b[82])^(a[213] & b[83])^(a[212] & b[84])^(a[211] & b[85])^(a[210] & b[86])^(a[209] & b[87])^(a[208] & b[88])^(a[207] & b[89])^(a[206] & b[90])^(a[205] & b[91])^(a[204] & b[92])^(a[203] & b[93])^(a[202] & b[94])^(a[201] & b[95])^(a[200] & b[96])^(a[199] & b[97])^(a[198] & b[98])^(a[197] & b[99])^(a[196] & b[100])^(a[195] & b[101])^(a[194] & b[102])^(a[193] & b[103])^(a[192] & b[104])^(a[191] & b[105])^(a[190] & b[106])^(a[189] & b[107])^(a[188] & b[108])^(a[187] & b[109])^(a[186] & b[110])^(a[185] & b[111])^(a[184] & b[112])^(a[183] & b[113])^(a[182] & b[114])^(a[181] & b[115])^(a[180] & b[116])^(a[179] & b[117])^(a[178] & b[118])^(a[177] & b[119])^(a[176] & b[120])^(a[175] & b[121])^(a[174] & b[122])^(a[173] & b[123])^(a[172] & b[124])^(a[171] & b[125])^(a[170] & b[126])^(a[169] & b[127])^(a[168] & b[128])^(a[167] & b[129])^(a[166] & b[130])^(a[165] & b[131])^(a[164] & b[132])^(a[163] & b[133])^(a[162] & b[134])^(a[161] & b[135])^(a[160] & b[136])^(a[159] & b[137])^(a[158] & b[138])^(a[157] & b[139])^(a[156] & b[140])^(a[155] & b[141])^(a[154] & b[142])^(a[153] & b[143])^(a[152] & b[144])^(a[151] & b[145])^(a[150] & b[146])^(a[149] & b[147])^(a[148] & b[148])^(a[147] & b[149])^(a[146] & b[150])^(a[145] & b[151])^(a[144] & b[152])^(a[143] & b[153])^(a[142] & b[154])^(a[141] & b[155])^(a[140] & b[156])^(a[139] & b[157])^(a[138] & b[158])^(a[137] & b[159])^(a[136] & b[160])^(a[135] & b[161])^(a[134] & b[162])^(a[133] & b[163])^(a[132] & b[164])^(a[131] & b[165])^(a[130] & b[166])^(a[129] & b[167])^(a[128] & b[168])^(a[127] & b[169])^(a[126] & b[170])^(a[125] & b[171])^(a[124] & b[172])^(a[123] & b[173])^(a[122] & b[174])^(a[121] & b[175])^(a[120] & b[176])^(a[119] & b[177])^(a[118] & b[178])^(a[117] & b[179])^(a[116] & b[180])^(a[115] & b[181])^(a[114] & b[182])^(a[113] & b[183])^(a[112] & b[184])^(a[111] & b[185])^(a[110] & b[186])^(a[109] & b[187])^(a[108] & b[188])^(a[107] & b[189])^(a[106] & b[190])^(a[105] & b[191])^(a[104] & b[192])^(a[103] & b[193])^(a[102] & b[194])^(a[101] & b[195])^(a[100] & b[196])^(a[99] & b[197])^(a[98] & b[198])^(a[97] & b[199])^(a[96] & b[200])^(a[95] & b[201])^(a[94] & b[202])^(a[93] & b[203])^(a[92] & b[204])^(a[91] & b[205])^(a[90] & b[206])^(a[89] & b[207])^(a[88] & b[208])^(a[87] & b[209])^(a[86] & b[210])^(a[85] & b[211])^(a[84] & b[212])^(a[83] & b[213])^(a[82] & b[214])^(a[81] & b[215])^(a[80] & b[216])^(a[79] & b[217])^(a[78] & b[218])^(a[77] & b[219])^(a[76] & b[220])^(a[75] & b[221])^(a[74] & b[222])^(a[73] & b[223])^(a[72] & b[224])^(a[71] & b[225])^(a[70] & b[226])^(a[69] & b[227])^(a[68] & b[228])^(a[67] & b[229])^(a[66] & b[230])^(a[65] & b[231])^(a[64] & b[232])^(a[63] & b[233])^(a[62] & b[234])^(a[61] & b[235])^(a[60] & b[236])^(a[59] & b[237])^(a[58] & b[238])^(a[57] & b[239])^(a[56] & b[240])^(a[55] & b[241])^(a[54] & b[242])^(a[53] & b[243])^(a[52] & b[244])^(a[51] & b[245])^(a[50] & b[246])^(a[49] & b[247])^(a[48] & b[248])^(a[47] & b[249])^(a[46] & b[250])^(a[45] & b[251])^(a[44] & b[252])^(a[43] & b[253])^(a[42] & b[254])^(a[41] & b[255])^(a[40] & b[256])^(a[39] & b[257])^(a[38] & b[258])^(a[37] & b[259])^(a[36] & b[260])^(a[35] & b[261])^(a[34] & b[262])^(a[33] & b[263])^(a[32] & b[264])^(a[31] & b[265])^(a[30] & b[266])^(a[29] & b[267])^(a[28] & b[268])^(a[27] & b[269])^(a[26] & b[270])^(a[25] & b[271])^(a[24] & b[272])^(a[23] & b[273])^(a[22] & b[274])^(a[21] & b[275])^(a[20] & b[276])^(a[19] & b[277])^(a[18] & b[278])^(a[17] & b[279])^(a[16] & b[280])^(a[15] & b[281])^(a[14] & b[282])^(a[13] & b[283])^(a[12] & b[284])^(a[11] & b[285])^(a[10] & b[286])^(a[9] & b[287])^(a[8] & b[288])^(a[7] & b[289])^(a[6] & b[290])^(a[5] & b[291])^(a[4] & b[292])^(a[3] & b[293])^(a[2] & b[294])^(a[1] & b[295])^(a[0] & b[296]);
assign y[297] = (a[297] & b[0])^(a[296] & b[1])^(a[295] & b[2])^(a[294] & b[3])^(a[293] & b[4])^(a[292] & b[5])^(a[291] & b[6])^(a[290] & b[7])^(a[289] & b[8])^(a[288] & b[9])^(a[287] & b[10])^(a[286] & b[11])^(a[285] & b[12])^(a[284] & b[13])^(a[283] & b[14])^(a[282] & b[15])^(a[281] & b[16])^(a[280] & b[17])^(a[279] & b[18])^(a[278] & b[19])^(a[277] & b[20])^(a[276] & b[21])^(a[275] & b[22])^(a[274] & b[23])^(a[273] & b[24])^(a[272] & b[25])^(a[271] & b[26])^(a[270] & b[27])^(a[269] & b[28])^(a[268] & b[29])^(a[267] & b[30])^(a[266] & b[31])^(a[265] & b[32])^(a[264] & b[33])^(a[263] & b[34])^(a[262] & b[35])^(a[261] & b[36])^(a[260] & b[37])^(a[259] & b[38])^(a[258] & b[39])^(a[257] & b[40])^(a[256] & b[41])^(a[255] & b[42])^(a[254] & b[43])^(a[253] & b[44])^(a[252] & b[45])^(a[251] & b[46])^(a[250] & b[47])^(a[249] & b[48])^(a[248] & b[49])^(a[247] & b[50])^(a[246] & b[51])^(a[245] & b[52])^(a[244] & b[53])^(a[243] & b[54])^(a[242] & b[55])^(a[241] & b[56])^(a[240] & b[57])^(a[239] & b[58])^(a[238] & b[59])^(a[237] & b[60])^(a[236] & b[61])^(a[235] & b[62])^(a[234] & b[63])^(a[233] & b[64])^(a[232] & b[65])^(a[231] & b[66])^(a[230] & b[67])^(a[229] & b[68])^(a[228] & b[69])^(a[227] & b[70])^(a[226] & b[71])^(a[225] & b[72])^(a[224] & b[73])^(a[223] & b[74])^(a[222] & b[75])^(a[221] & b[76])^(a[220] & b[77])^(a[219] & b[78])^(a[218] & b[79])^(a[217] & b[80])^(a[216] & b[81])^(a[215] & b[82])^(a[214] & b[83])^(a[213] & b[84])^(a[212] & b[85])^(a[211] & b[86])^(a[210] & b[87])^(a[209] & b[88])^(a[208] & b[89])^(a[207] & b[90])^(a[206] & b[91])^(a[205] & b[92])^(a[204] & b[93])^(a[203] & b[94])^(a[202] & b[95])^(a[201] & b[96])^(a[200] & b[97])^(a[199] & b[98])^(a[198] & b[99])^(a[197] & b[100])^(a[196] & b[101])^(a[195] & b[102])^(a[194] & b[103])^(a[193] & b[104])^(a[192] & b[105])^(a[191] & b[106])^(a[190] & b[107])^(a[189] & b[108])^(a[188] & b[109])^(a[187] & b[110])^(a[186] & b[111])^(a[185] & b[112])^(a[184] & b[113])^(a[183] & b[114])^(a[182] & b[115])^(a[181] & b[116])^(a[180] & b[117])^(a[179] & b[118])^(a[178] & b[119])^(a[177] & b[120])^(a[176] & b[121])^(a[175] & b[122])^(a[174] & b[123])^(a[173] & b[124])^(a[172] & b[125])^(a[171] & b[126])^(a[170] & b[127])^(a[169] & b[128])^(a[168] & b[129])^(a[167] & b[130])^(a[166] & b[131])^(a[165] & b[132])^(a[164] & b[133])^(a[163] & b[134])^(a[162] & b[135])^(a[161] & b[136])^(a[160] & b[137])^(a[159] & b[138])^(a[158] & b[139])^(a[157] & b[140])^(a[156] & b[141])^(a[155] & b[142])^(a[154] & b[143])^(a[153] & b[144])^(a[152] & b[145])^(a[151] & b[146])^(a[150] & b[147])^(a[149] & b[148])^(a[148] & b[149])^(a[147] & b[150])^(a[146] & b[151])^(a[145] & b[152])^(a[144] & b[153])^(a[143] & b[154])^(a[142] & b[155])^(a[141] & b[156])^(a[140] & b[157])^(a[139] & b[158])^(a[138] & b[159])^(a[137] & b[160])^(a[136] & b[161])^(a[135] & b[162])^(a[134] & b[163])^(a[133] & b[164])^(a[132] & b[165])^(a[131] & b[166])^(a[130] & b[167])^(a[129] & b[168])^(a[128] & b[169])^(a[127] & b[170])^(a[126] & b[171])^(a[125] & b[172])^(a[124] & b[173])^(a[123] & b[174])^(a[122] & b[175])^(a[121] & b[176])^(a[120] & b[177])^(a[119] & b[178])^(a[118] & b[179])^(a[117] & b[180])^(a[116] & b[181])^(a[115] & b[182])^(a[114] & b[183])^(a[113] & b[184])^(a[112] & b[185])^(a[111] & b[186])^(a[110] & b[187])^(a[109] & b[188])^(a[108] & b[189])^(a[107] & b[190])^(a[106] & b[191])^(a[105] & b[192])^(a[104] & b[193])^(a[103] & b[194])^(a[102] & b[195])^(a[101] & b[196])^(a[100] & b[197])^(a[99] & b[198])^(a[98] & b[199])^(a[97] & b[200])^(a[96] & b[201])^(a[95] & b[202])^(a[94] & b[203])^(a[93] & b[204])^(a[92] & b[205])^(a[91] & b[206])^(a[90] & b[207])^(a[89] & b[208])^(a[88] & b[209])^(a[87] & b[210])^(a[86] & b[211])^(a[85] & b[212])^(a[84] & b[213])^(a[83] & b[214])^(a[82] & b[215])^(a[81] & b[216])^(a[80] & b[217])^(a[79] & b[218])^(a[78] & b[219])^(a[77] & b[220])^(a[76] & b[221])^(a[75] & b[222])^(a[74] & b[223])^(a[73] & b[224])^(a[72] & b[225])^(a[71] & b[226])^(a[70] & b[227])^(a[69] & b[228])^(a[68] & b[229])^(a[67] & b[230])^(a[66] & b[231])^(a[65] & b[232])^(a[64] & b[233])^(a[63] & b[234])^(a[62] & b[235])^(a[61] & b[236])^(a[60] & b[237])^(a[59] & b[238])^(a[58] & b[239])^(a[57] & b[240])^(a[56] & b[241])^(a[55] & b[242])^(a[54] & b[243])^(a[53] & b[244])^(a[52] & b[245])^(a[51] & b[246])^(a[50] & b[247])^(a[49] & b[248])^(a[48] & b[249])^(a[47] & b[250])^(a[46] & b[251])^(a[45] & b[252])^(a[44] & b[253])^(a[43] & b[254])^(a[42] & b[255])^(a[41] & b[256])^(a[40] & b[257])^(a[39] & b[258])^(a[38] & b[259])^(a[37] & b[260])^(a[36] & b[261])^(a[35] & b[262])^(a[34] & b[263])^(a[33] & b[264])^(a[32] & b[265])^(a[31] & b[266])^(a[30] & b[267])^(a[29] & b[268])^(a[28] & b[269])^(a[27] & b[270])^(a[26] & b[271])^(a[25] & b[272])^(a[24] & b[273])^(a[23] & b[274])^(a[22] & b[275])^(a[21] & b[276])^(a[20] & b[277])^(a[19] & b[278])^(a[18] & b[279])^(a[17] & b[280])^(a[16] & b[281])^(a[15] & b[282])^(a[14] & b[283])^(a[13] & b[284])^(a[12] & b[285])^(a[11] & b[286])^(a[10] & b[287])^(a[9] & b[288])^(a[8] & b[289])^(a[7] & b[290])^(a[6] & b[291])^(a[5] & b[292])^(a[4] & b[293])^(a[3] & b[294])^(a[2] & b[295])^(a[1] & b[296])^(a[0] & b[297]);
assign y[298] = (a[298] & b[0])^(a[297] & b[1])^(a[296] & b[2])^(a[295] & b[3])^(a[294] & b[4])^(a[293] & b[5])^(a[292] & b[6])^(a[291] & b[7])^(a[290] & b[8])^(a[289] & b[9])^(a[288] & b[10])^(a[287] & b[11])^(a[286] & b[12])^(a[285] & b[13])^(a[284] & b[14])^(a[283] & b[15])^(a[282] & b[16])^(a[281] & b[17])^(a[280] & b[18])^(a[279] & b[19])^(a[278] & b[20])^(a[277] & b[21])^(a[276] & b[22])^(a[275] & b[23])^(a[274] & b[24])^(a[273] & b[25])^(a[272] & b[26])^(a[271] & b[27])^(a[270] & b[28])^(a[269] & b[29])^(a[268] & b[30])^(a[267] & b[31])^(a[266] & b[32])^(a[265] & b[33])^(a[264] & b[34])^(a[263] & b[35])^(a[262] & b[36])^(a[261] & b[37])^(a[260] & b[38])^(a[259] & b[39])^(a[258] & b[40])^(a[257] & b[41])^(a[256] & b[42])^(a[255] & b[43])^(a[254] & b[44])^(a[253] & b[45])^(a[252] & b[46])^(a[251] & b[47])^(a[250] & b[48])^(a[249] & b[49])^(a[248] & b[50])^(a[247] & b[51])^(a[246] & b[52])^(a[245] & b[53])^(a[244] & b[54])^(a[243] & b[55])^(a[242] & b[56])^(a[241] & b[57])^(a[240] & b[58])^(a[239] & b[59])^(a[238] & b[60])^(a[237] & b[61])^(a[236] & b[62])^(a[235] & b[63])^(a[234] & b[64])^(a[233] & b[65])^(a[232] & b[66])^(a[231] & b[67])^(a[230] & b[68])^(a[229] & b[69])^(a[228] & b[70])^(a[227] & b[71])^(a[226] & b[72])^(a[225] & b[73])^(a[224] & b[74])^(a[223] & b[75])^(a[222] & b[76])^(a[221] & b[77])^(a[220] & b[78])^(a[219] & b[79])^(a[218] & b[80])^(a[217] & b[81])^(a[216] & b[82])^(a[215] & b[83])^(a[214] & b[84])^(a[213] & b[85])^(a[212] & b[86])^(a[211] & b[87])^(a[210] & b[88])^(a[209] & b[89])^(a[208] & b[90])^(a[207] & b[91])^(a[206] & b[92])^(a[205] & b[93])^(a[204] & b[94])^(a[203] & b[95])^(a[202] & b[96])^(a[201] & b[97])^(a[200] & b[98])^(a[199] & b[99])^(a[198] & b[100])^(a[197] & b[101])^(a[196] & b[102])^(a[195] & b[103])^(a[194] & b[104])^(a[193] & b[105])^(a[192] & b[106])^(a[191] & b[107])^(a[190] & b[108])^(a[189] & b[109])^(a[188] & b[110])^(a[187] & b[111])^(a[186] & b[112])^(a[185] & b[113])^(a[184] & b[114])^(a[183] & b[115])^(a[182] & b[116])^(a[181] & b[117])^(a[180] & b[118])^(a[179] & b[119])^(a[178] & b[120])^(a[177] & b[121])^(a[176] & b[122])^(a[175] & b[123])^(a[174] & b[124])^(a[173] & b[125])^(a[172] & b[126])^(a[171] & b[127])^(a[170] & b[128])^(a[169] & b[129])^(a[168] & b[130])^(a[167] & b[131])^(a[166] & b[132])^(a[165] & b[133])^(a[164] & b[134])^(a[163] & b[135])^(a[162] & b[136])^(a[161] & b[137])^(a[160] & b[138])^(a[159] & b[139])^(a[158] & b[140])^(a[157] & b[141])^(a[156] & b[142])^(a[155] & b[143])^(a[154] & b[144])^(a[153] & b[145])^(a[152] & b[146])^(a[151] & b[147])^(a[150] & b[148])^(a[149] & b[149])^(a[148] & b[150])^(a[147] & b[151])^(a[146] & b[152])^(a[145] & b[153])^(a[144] & b[154])^(a[143] & b[155])^(a[142] & b[156])^(a[141] & b[157])^(a[140] & b[158])^(a[139] & b[159])^(a[138] & b[160])^(a[137] & b[161])^(a[136] & b[162])^(a[135] & b[163])^(a[134] & b[164])^(a[133] & b[165])^(a[132] & b[166])^(a[131] & b[167])^(a[130] & b[168])^(a[129] & b[169])^(a[128] & b[170])^(a[127] & b[171])^(a[126] & b[172])^(a[125] & b[173])^(a[124] & b[174])^(a[123] & b[175])^(a[122] & b[176])^(a[121] & b[177])^(a[120] & b[178])^(a[119] & b[179])^(a[118] & b[180])^(a[117] & b[181])^(a[116] & b[182])^(a[115] & b[183])^(a[114] & b[184])^(a[113] & b[185])^(a[112] & b[186])^(a[111] & b[187])^(a[110] & b[188])^(a[109] & b[189])^(a[108] & b[190])^(a[107] & b[191])^(a[106] & b[192])^(a[105] & b[193])^(a[104] & b[194])^(a[103] & b[195])^(a[102] & b[196])^(a[101] & b[197])^(a[100] & b[198])^(a[99] & b[199])^(a[98] & b[200])^(a[97] & b[201])^(a[96] & b[202])^(a[95] & b[203])^(a[94] & b[204])^(a[93] & b[205])^(a[92] & b[206])^(a[91] & b[207])^(a[90] & b[208])^(a[89] & b[209])^(a[88] & b[210])^(a[87] & b[211])^(a[86] & b[212])^(a[85] & b[213])^(a[84] & b[214])^(a[83] & b[215])^(a[82] & b[216])^(a[81] & b[217])^(a[80] & b[218])^(a[79] & b[219])^(a[78] & b[220])^(a[77] & b[221])^(a[76] & b[222])^(a[75] & b[223])^(a[74] & b[224])^(a[73] & b[225])^(a[72] & b[226])^(a[71] & b[227])^(a[70] & b[228])^(a[69] & b[229])^(a[68] & b[230])^(a[67] & b[231])^(a[66] & b[232])^(a[65] & b[233])^(a[64] & b[234])^(a[63] & b[235])^(a[62] & b[236])^(a[61] & b[237])^(a[60] & b[238])^(a[59] & b[239])^(a[58] & b[240])^(a[57] & b[241])^(a[56] & b[242])^(a[55] & b[243])^(a[54] & b[244])^(a[53] & b[245])^(a[52] & b[246])^(a[51] & b[247])^(a[50] & b[248])^(a[49] & b[249])^(a[48] & b[250])^(a[47] & b[251])^(a[46] & b[252])^(a[45] & b[253])^(a[44] & b[254])^(a[43] & b[255])^(a[42] & b[256])^(a[41] & b[257])^(a[40] & b[258])^(a[39] & b[259])^(a[38] & b[260])^(a[37] & b[261])^(a[36] & b[262])^(a[35] & b[263])^(a[34] & b[264])^(a[33] & b[265])^(a[32] & b[266])^(a[31] & b[267])^(a[30] & b[268])^(a[29] & b[269])^(a[28] & b[270])^(a[27] & b[271])^(a[26] & b[272])^(a[25] & b[273])^(a[24] & b[274])^(a[23] & b[275])^(a[22] & b[276])^(a[21] & b[277])^(a[20] & b[278])^(a[19] & b[279])^(a[18] & b[280])^(a[17] & b[281])^(a[16] & b[282])^(a[15] & b[283])^(a[14] & b[284])^(a[13] & b[285])^(a[12] & b[286])^(a[11] & b[287])^(a[10] & b[288])^(a[9] & b[289])^(a[8] & b[290])^(a[7] & b[291])^(a[6] & b[292])^(a[5] & b[293])^(a[4] & b[294])^(a[3] & b[295])^(a[2] & b[296])^(a[1] & b[297])^(a[0] & b[298]);
assign y[299] = (a[299] & b[0])^(a[298] & b[1])^(a[297] & b[2])^(a[296] & b[3])^(a[295] & b[4])^(a[294] & b[5])^(a[293] & b[6])^(a[292] & b[7])^(a[291] & b[8])^(a[290] & b[9])^(a[289] & b[10])^(a[288] & b[11])^(a[287] & b[12])^(a[286] & b[13])^(a[285] & b[14])^(a[284] & b[15])^(a[283] & b[16])^(a[282] & b[17])^(a[281] & b[18])^(a[280] & b[19])^(a[279] & b[20])^(a[278] & b[21])^(a[277] & b[22])^(a[276] & b[23])^(a[275] & b[24])^(a[274] & b[25])^(a[273] & b[26])^(a[272] & b[27])^(a[271] & b[28])^(a[270] & b[29])^(a[269] & b[30])^(a[268] & b[31])^(a[267] & b[32])^(a[266] & b[33])^(a[265] & b[34])^(a[264] & b[35])^(a[263] & b[36])^(a[262] & b[37])^(a[261] & b[38])^(a[260] & b[39])^(a[259] & b[40])^(a[258] & b[41])^(a[257] & b[42])^(a[256] & b[43])^(a[255] & b[44])^(a[254] & b[45])^(a[253] & b[46])^(a[252] & b[47])^(a[251] & b[48])^(a[250] & b[49])^(a[249] & b[50])^(a[248] & b[51])^(a[247] & b[52])^(a[246] & b[53])^(a[245] & b[54])^(a[244] & b[55])^(a[243] & b[56])^(a[242] & b[57])^(a[241] & b[58])^(a[240] & b[59])^(a[239] & b[60])^(a[238] & b[61])^(a[237] & b[62])^(a[236] & b[63])^(a[235] & b[64])^(a[234] & b[65])^(a[233] & b[66])^(a[232] & b[67])^(a[231] & b[68])^(a[230] & b[69])^(a[229] & b[70])^(a[228] & b[71])^(a[227] & b[72])^(a[226] & b[73])^(a[225] & b[74])^(a[224] & b[75])^(a[223] & b[76])^(a[222] & b[77])^(a[221] & b[78])^(a[220] & b[79])^(a[219] & b[80])^(a[218] & b[81])^(a[217] & b[82])^(a[216] & b[83])^(a[215] & b[84])^(a[214] & b[85])^(a[213] & b[86])^(a[212] & b[87])^(a[211] & b[88])^(a[210] & b[89])^(a[209] & b[90])^(a[208] & b[91])^(a[207] & b[92])^(a[206] & b[93])^(a[205] & b[94])^(a[204] & b[95])^(a[203] & b[96])^(a[202] & b[97])^(a[201] & b[98])^(a[200] & b[99])^(a[199] & b[100])^(a[198] & b[101])^(a[197] & b[102])^(a[196] & b[103])^(a[195] & b[104])^(a[194] & b[105])^(a[193] & b[106])^(a[192] & b[107])^(a[191] & b[108])^(a[190] & b[109])^(a[189] & b[110])^(a[188] & b[111])^(a[187] & b[112])^(a[186] & b[113])^(a[185] & b[114])^(a[184] & b[115])^(a[183] & b[116])^(a[182] & b[117])^(a[181] & b[118])^(a[180] & b[119])^(a[179] & b[120])^(a[178] & b[121])^(a[177] & b[122])^(a[176] & b[123])^(a[175] & b[124])^(a[174] & b[125])^(a[173] & b[126])^(a[172] & b[127])^(a[171] & b[128])^(a[170] & b[129])^(a[169] & b[130])^(a[168] & b[131])^(a[167] & b[132])^(a[166] & b[133])^(a[165] & b[134])^(a[164] & b[135])^(a[163] & b[136])^(a[162] & b[137])^(a[161] & b[138])^(a[160] & b[139])^(a[159] & b[140])^(a[158] & b[141])^(a[157] & b[142])^(a[156] & b[143])^(a[155] & b[144])^(a[154] & b[145])^(a[153] & b[146])^(a[152] & b[147])^(a[151] & b[148])^(a[150] & b[149])^(a[149] & b[150])^(a[148] & b[151])^(a[147] & b[152])^(a[146] & b[153])^(a[145] & b[154])^(a[144] & b[155])^(a[143] & b[156])^(a[142] & b[157])^(a[141] & b[158])^(a[140] & b[159])^(a[139] & b[160])^(a[138] & b[161])^(a[137] & b[162])^(a[136] & b[163])^(a[135] & b[164])^(a[134] & b[165])^(a[133] & b[166])^(a[132] & b[167])^(a[131] & b[168])^(a[130] & b[169])^(a[129] & b[170])^(a[128] & b[171])^(a[127] & b[172])^(a[126] & b[173])^(a[125] & b[174])^(a[124] & b[175])^(a[123] & b[176])^(a[122] & b[177])^(a[121] & b[178])^(a[120] & b[179])^(a[119] & b[180])^(a[118] & b[181])^(a[117] & b[182])^(a[116] & b[183])^(a[115] & b[184])^(a[114] & b[185])^(a[113] & b[186])^(a[112] & b[187])^(a[111] & b[188])^(a[110] & b[189])^(a[109] & b[190])^(a[108] & b[191])^(a[107] & b[192])^(a[106] & b[193])^(a[105] & b[194])^(a[104] & b[195])^(a[103] & b[196])^(a[102] & b[197])^(a[101] & b[198])^(a[100] & b[199])^(a[99] & b[200])^(a[98] & b[201])^(a[97] & b[202])^(a[96] & b[203])^(a[95] & b[204])^(a[94] & b[205])^(a[93] & b[206])^(a[92] & b[207])^(a[91] & b[208])^(a[90] & b[209])^(a[89] & b[210])^(a[88] & b[211])^(a[87] & b[212])^(a[86] & b[213])^(a[85] & b[214])^(a[84] & b[215])^(a[83] & b[216])^(a[82] & b[217])^(a[81] & b[218])^(a[80] & b[219])^(a[79] & b[220])^(a[78] & b[221])^(a[77] & b[222])^(a[76] & b[223])^(a[75] & b[224])^(a[74] & b[225])^(a[73] & b[226])^(a[72] & b[227])^(a[71] & b[228])^(a[70] & b[229])^(a[69] & b[230])^(a[68] & b[231])^(a[67] & b[232])^(a[66] & b[233])^(a[65] & b[234])^(a[64] & b[235])^(a[63] & b[236])^(a[62] & b[237])^(a[61] & b[238])^(a[60] & b[239])^(a[59] & b[240])^(a[58] & b[241])^(a[57] & b[242])^(a[56] & b[243])^(a[55] & b[244])^(a[54] & b[245])^(a[53] & b[246])^(a[52] & b[247])^(a[51] & b[248])^(a[50] & b[249])^(a[49] & b[250])^(a[48] & b[251])^(a[47] & b[252])^(a[46] & b[253])^(a[45] & b[254])^(a[44] & b[255])^(a[43] & b[256])^(a[42] & b[257])^(a[41] & b[258])^(a[40] & b[259])^(a[39] & b[260])^(a[38] & b[261])^(a[37] & b[262])^(a[36] & b[263])^(a[35] & b[264])^(a[34] & b[265])^(a[33] & b[266])^(a[32] & b[267])^(a[31] & b[268])^(a[30] & b[269])^(a[29] & b[270])^(a[28] & b[271])^(a[27] & b[272])^(a[26] & b[273])^(a[25] & b[274])^(a[24] & b[275])^(a[23] & b[276])^(a[22] & b[277])^(a[21] & b[278])^(a[20] & b[279])^(a[19] & b[280])^(a[18] & b[281])^(a[17] & b[282])^(a[16] & b[283])^(a[15] & b[284])^(a[14] & b[285])^(a[13] & b[286])^(a[12] & b[287])^(a[11] & b[288])^(a[10] & b[289])^(a[9] & b[290])^(a[8] & b[291])^(a[7] & b[292])^(a[6] & b[293])^(a[5] & b[294])^(a[4] & b[295])^(a[3] & b[296])^(a[2] & b[297])^(a[1] & b[298])^(a[0] & b[299]);
assign y[300] = (a[300] & b[0])^(a[299] & b[1])^(a[298] & b[2])^(a[297] & b[3])^(a[296] & b[4])^(a[295] & b[5])^(a[294] & b[6])^(a[293] & b[7])^(a[292] & b[8])^(a[291] & b[9])^(a[290] & b[10])^(a[289] & b[11])^(a[288] & b[12])^(a[287] & b[13])^(a[286] & b[14])^(a[285] & b[15])^(a[284] & b[16])^(a[283] & b[17])^(a[282] & b[18])^(a[281] & b[19])^(a[280] & b[20])^(a[279] & b[21])^(a[278] & b[22])^(a[277] & b[23])^(a[276] & b[24])^(a[275] & b[25])^(a[274] & b[26])^(a[273] & b[27])^(a[272] & b[28])^(a[271] & b[29])^(a[270] & b[30])^(a[269] & b[31])^(a[268] & b[32])^(a[267] & b[33])^(a[266] & b[34])^(a[265] & b[35])^(a[264] & b[36])^(a[263] & b[37])^(a[262] & b[38])^(a[261] & b[39])^(a[260] & b[40])^(a[259] & b[41])^(a[258] & b[42])^(a[257] & b[43])^(a[256] & b[44])^(a[255] & b[45])^(a[254] & b[46])^(a[253] & b[47])^(a[252] & b[48])^(a[251] & b[49])^(a[250] & b[50])^(a[249] & b[51])^(a[248] & b[52])^(a[247] & b[53])^(a[246] & b[54])^(a[245] & b[55])^(a[244] & b[56])^(a[243] & b[57])^(a[242] & b[58])^(a[241] & b[59])^(a[240] & b[60])^(a[239] & b[61])^(a[238] & b[62])^(a[237] & b[63])^(a[236] & b[64])^(a[235] & b[65])^(a[234] & b[66])^(a[233] & b[67])^(a[232] & b[68])^(a[231] & b[69])^(a[230] & b[70])^(a[229] & b[71])^(a[228] & b[72])^(a[227] & b[73])^(a[226] & b[74])^(a[225] & b[75])^(a[224] & b[76])^(a[223] & b[77])^(a[222] & b[78])^(a[221] & b[79])^(a[220] & b[80])^(a[219] & b[81])^(a[218] & b[82])^(a[217] & b[83])^(a[216] & b[84])^(a[215] & b[85])^(a[214] & b[86])^(a[213] & b[87])^(a[212] & b[88])^(a[211] & b[89])^(a[210] & b[90])^(a[209] & b[91])^(a[208] & b[92])^(a[207] & b[93])^(a[206] & b[94])^(a[205] & b[95])^(a[204] & b[96])^(a[203] & b[97])^(a[202] & b[98])^(a[201] & b[99])^(a[200] & b[100])^(a[199] & b[101])^(a[198] & b[102])^(a[197] & b[103])^(a[196] & b[104])^(a[195] & b[105])^(a[194] & b[106])^(a[193] & b[107])^(a[192] & b[108])^(a[191] & b[109])^(a[190] & b[110])^(a[189] & b[111])^(a[188] & b[112])^(a[187] & b[113])^(a[186] & b[114])^(a[185] & b[115])^(a[184] & b[116])^(a[183] & b[117])^(a[182] & b[118])^(a[181] & b[119])^(a[180] & b[120])^(a[179] & b[121])^(a[178] & b[122])^(a[177] & b[123])^(a[176] & b[124])^(a[175] & b[125])^(a[174] & b[126])^(a[173] & b[127])^(a[172] & b[128])^(a[171] & b[129])^(a[170] & b[130])^(a[169] & b[131])^(a[168] & b[132])^(a[167] & b[133])^(a[166] & b[134])^(a[165] & b[135])^(a[164] & b[136])^(a[163] & b[137])^(a[162] & b[138])^(a[161] & b[139])^(a[160] & b[140])^(a[159] & b[141])^(a[158] & b[142])^(a[157] & b[143])^(a[156] & b[144])^(a[155] & b[145])^(a[154] & b[146])^(a[153] & b[147])^(a[152] & b[148])^(a[151] & b[149])^(a[150] & b[150])^(a[149] & b[151])^(a[148] & b[152])^(a[147] & b[153])^(a[146] & b[154])^(a[145] & b[155])^(a[144] & b[156])^(a[143] & b[157])^(a[142] & b[158])^(a[141] & b[159])^(a[140] & b[160])^(a[139] & b[161])^(a[138] & b[162])^(a[137] & b[163])^(a[136] & b[164])^(a[135] & b[165])^(a[134] & b[166])^(a[133] & b[167])^(a[132] & b[168])^(a[131] & b[169])^(a[130] & b[170])^(a[129] & b[171])^(a[128] & b[172])^(a[127] & b[173])^(a[126] & b[174])^(a[125] & b[175])^(a[124] & b[176])^(a[123] & b[177])^(a[122] & b[178])^(a[121] & b[179])^(a[120] & b[180])^(a[119] & b[181])^(a[118] & b[182])^(a[117] & b[183])^(a[116] & b[184])^(a[115] & b[185])^(a[114] & b[186])^(a[113] & b[187])^(a[112] & b[188])^(a[111] & b[189])^(a[110] & b[190])^(a[109] & b[191])^(a[108] & b[192])^(a[107] & b[193])^(a[106] & b[194])^(a[105] & b[195])^(a[104] & b[196])^(a[103] & b[197])^(a[102] & b[198])^(a[101] & b[199])^(a[100] & b[200])^(a[99] & b[201])^(a[98] & b[202])^(a[97] & b[203])^(a[96] & b[204])^(a[95] & b[205])^(a[94] & b[206])^(a[93] & b[207])^(a[92] & b[208])^(a[91] & b[209])^(a[90] & b[210])^(a[89] & b[211])^(a[88] & b[212])^(a[87] & b[213])^(a[86] & b[214])^(a[85] & b[215])^(a[84] & b[216])^(a[83] & b[217])^(a[82] & b[218])^(a[81] & b[219])^(a[80] & b[220])^(a[79] & b[221])^(a[78] & b[222])^(a[77] & b[223])^(a[76] & b[224])^(a[75] & b[225])^(a[74] & b[226])^(a[73] & b[227])^(a[72] & b[228])^(a[71] & b[229])^(a[70] & b[230])^(a[69] & b[231])^(a[68] & b[232])^(a[67] & b[233])^(a[66] & b[234])^(a[65] & b[235])^(a[64] & b[236])^(a[63] & b[237])^(a[62] & b[238])^(a[61] & b[239])^(a[60] & b[240])^(a[59] & b[241])^(a[58] & b[242])^(a[57] & b[243])^(a[56] & b[244])^(a[55] & b[245])^(a[54] & b[246])^(a[53] & b[247])^(a[52] & b[248])^(a[51] & b[249])^(a[50] & b[250])^(a[49] & b[251])^(a[48] & b[252])^(a[47] & b[253])^(a[46] & b[254])^(a[45] & b[255])^(a[44] & b[256])^(a[43] & b[257])^(a[42] & b[258])^(a[41] & b[259])^(a[40] & b[260])^(a[39] & b[261])^(a[38] & b[262])^(a[37] & b[263])^(a[36] & b[264])^(a[35] & b[265])^(a[34] & b[266])^(a[33] & b[267])^(a[32] & b[268])^(a[31] & b[269])^(a[30] & b[270])^(a[29] & b[271])^(a[28] & b[272])^(a[27] & b[273])^(a[26] & b[274])^(a[25] & b[275])^(a[24] & b[276])^(a[23] & b[277])^(a[22] & b[278])^(a[21] & b[279])^(a[20] & b[280])^(a[19] & b[281])^(a[18] & b[282])^(a[17] & b[283])^(a[16] & b[284])^(a[15] & b[285])^(a[14] & b[286])^(a[13] & b[287])^(a[12] & b[288])^(a[11] & b[289])^(a[10] & b[290])^(a[9] & b[291])^(a[8] & b[292])^(a[7] & b[293])^(a[6] & b[294])^(a[5] & b[295])^(a[4] & b[296])^(a[3] & b[297])^(a[2] & b[298])^(a[1] & b[299])^(a[0] & b[300]);
assign y[301] = (a[301] & b[0])^(a[300] & b[1])^(a[299] & b[2])^(a[298] & b[3])^(a[297] & b[4])^(a[296] & b[5])^(a[295] & b[6])^(a[294] & b[7])^(a[293] & b[8])^(a[292] & b[9])^(a[291] & b[10])^(a[290] & b[11])^(a[289] & b[12])^(a[288] & b[13])^(a[287] & b[14])^(a[286] & b[15])^(a[285] & b[16])^(a[284] & b[17])^(a[283] & b[18])^(a[282] & b[19])^(a[281] & b[20])^(a[280] & b[21])^(a[279] & b[22])^(a[278] & b[23])^(a[277] & b[24])^(a[276] & b[25])^(a[275] & b[26])^(a[274] & b[27])^(a[273] & b[28])^(a[272] & b[29])^(a[271] & b[30])^(a[270] & b[31])^(a[269] & b[32])^(a[268] & b[33])^(a[267] & b[34])^(a[266] & b[35])^(a[265] & b[36])^(a[264] & b[37])^(a[263] & b[38])^(a[262] & b[39])^(a[261] & b[40])^(a[260] & b[41])^(a[259] & b[42])^(a[258] & b[43])^(a[257] & b[44])^(a[256] & b[45])^(a[255] & b[46])^(a[254] & b[47])^(a[253] & b[48])^(a[252] & b[49])^(a[251] & b[50])^(a[250] & b[51])^(a[249] & b[52])^(a[248] & b[53])^(a[247] & b[54])^(a[246] & b[55])^(a[245] & b[56])^(a[244] & b[57])^(a[243] & b[58])^(a[242] & b[59])^(a[241] & b[60])^(a[240] & b[61])^(a[239] & b[62])^(a[238] & b[63])^(a[237] & b[64])^(a[236] & b[65])^(a[235] & b[66])^(a[234] & b[67])^(a[233] & b[68])^(a[232] & b[69])^(a[231] & b[70])^(a[230] & b[71])^(a[229] & b[72])^(a[228] & b[73])^(a[227] & b[74])^(a[226] & b[75])^(a[225] & b[76])^(a[224] & b[77])^(a[223] & b[78])^(a[222] & b[79])^(a[221] & b[80])^(a[220] & b[81])^(a[219] & b[82])^(a[218] & b[83])^(a[217] & b[84])^(a[216] & b[85])^(a[215] & b[86])^(a[214] & b[87])^(a[213] & b[88])^(a[212] & b[89])^(a[211] & b[90])^(a[210] & b[91])^(a[209] & b[92])^(a[208] & b[93])^(a[207] & b[94])^(a[206] & b[95])^(a[205] & b[96])^(a[204] & b[97])^(a[203] & b[98])^(a[202] & b[99])^(a[201] & b[100])^(a[200] & b[101])^(a[199] & b[102])^(a[198] & b[103])^(a[197] & b[104])^(a[196] & b[105])^(a[195] & b[106])^(a[194] & b[107])^(a[193] & b[108])^(a[192] & b[109])^(a[191] & b[110])^(a[190] & b[111])^(a[189] & b[112])^(a[188] & b[113])^(a[187] & b[114])^(a[186] & b[115])^(a[185] & b[116])^(a[184] & b[117])^(a[183] & b[118])^(a[182] & b[119])^(a[181] & b[120])^(a[180] & b[121])^(a[179] & b[122])^(a[178] & b[123])^(a[177] & b[124])^(a[176] & b[125])^(a[175] & b[126])^(a[174] & b[127])^(a[173] & b[128])^(a[172] & b[129])^(a[171] & b[130])^(a[170] & b[131])^(a[169] & b[132])^(a[168] & b[133])^(a[167] & b[134])^(a[166] & b[135])^(a[165] & b[136])^(a[164] & b[137])^(a[163] & b[138])^(a[162] & b[139])^(a[161] & b[140])^(a[160] & b[141])^(a[159] & b[142])^(a[158] & b[143])^(a[157] & b[144])^(a[156] & b[145])^(a[155] & b[146])^(a[154] & b[147])^(a[153] & b[148])^(a[152] & b[149])^(a[151] & b[150])^(a[150] & b[151])^(a[149] & b[152])^(a[148] & b[153])^(a[147] & b[154])^(a[146] & b[155])^(a[145] & b[156])^(a[144] & b[157])^(a[143] & b[158])^(a[142] & b[159])^(a[141] & b[160])^(a[140] & b[161])^(a[139] & b[162])^(a[138] & b[163])^(a[137] & b[164])^(a[136] & b[165])^(a[135] & b[166])^(a[134] & b[167])^(a[133] & b[168])^(a[132] & b[169])^(a[131] & b[170])^(a[130] & b[171])^(a[129] & b[172])^(a[128] & b[173])^(a[127] & b[174])^(a[126] & b[175])^(a[125] & b[176])^(a[124] & b[177])^(a[123] & b[178])^(a[122] & b[179])^(a[121] & b[180])^(a[120] & b[181])^(a[119] & b[182])^(a[118] & b[183])^(a[117] & b[184])^(a[116] & b[185])^(a[115] & b[186])^(a[114] & b[187])^(a[113] & b[188])^(a[112] & b[189])^(a[111] & b[190])^(a[110] & b[191])^(a[109] & b[192])^(a[108] & b[193])^(a[107] & b[194])^(a[106] & b[195])^(a[105] & b[196])^(a[104] & b[197])^(a[103] & b[198])^(a[102] & b[199])^(a[101] & b[200])^(a[100] & b[201])^(a[99] & b[202])^(a[98] & b[203])^(a[97] & b[204])^(a[96] & b[205])^(a[95] & b[206])^(a[94] & b[207])^(a[93] & b[208])^(a[92] & b[209])^(a[91] & b[210])^(a[90] & b[211])^(a[89] & b[212])^(a[88] & b[213])^(a[87] & b[214])^(a[86] & b[215])^(a[85] & b[216])^(a[84] & b[217])^(a[83] & b[218])^(a[82] & b[219])^(a[81] & b[220])^(a[80] & b[221])^(a[79] & b[222])^(a[78] & b[223])^(a[77] & b[224])^(a[76] & b[225])^(a[75] & b[226])^(a[74] & b[227])^(a[73] & b[228])^(a[72] & b[229])^(a[71] & b[230])^(a[70] & b[231])^(a[69] & b[232])^(a[68] & b[233])^(a[67] & b[234])^(a[66] & b[235])^(a[65] & b[236])^(a[64] & b[237])^(a[63] & b[238])^(a[62] & b[239])^(a[61] & b[240])^(a[60] & b[241])^(a[59] & b[242])^(a[58] & b[243])^(a[57] & b[244])^(a[56] & b[245])^(a[55] & b[246])^(a[54] & b[247])^(a[53] & b[248])^(a[52] & b[249])^(a[51] & b[250])^(a[50] & b[251])^(a[49] & b[252])^(a[48] & b[253])^(a[47] & b[254])^(a[46] & b[255])^(a[45] & b[256])^(a[44] & b[257])^(a[43] & b[258])^(a[42] & b[259])^(a[41] & b[260])^(a[40] & b[261])^(a[39] & b[262])^(a[38] & b[263])^(a[37] & b[264])^(a[36] & b[265])^(a[35] & b[266])^(a[34] & b[267])^(a[33] & b[268])^(a[32] & b[269])^(a[31] & b[270])^(a[30] & b[271])^(a[29] & b[272])^(a[28] & b[273])^(a[27] & b[274])^(a[26] & b[275])^(a[25] & b[276])^(a[24] & b[277])^(a[23] & b[278])^(a[22] & b[279])^(a[21] & b[280])^(a[20] & b[281])^(a[19] & b[282])^(a[18] & b[283])^(a[17] & b[284])^(a[16] & b[285])^(a[15] & b[286])^(a[14] & b[287])^(a[13] & b[288])^(a[12] & b[289])^(a[11] & b[290])^(a[10] & b[291])^(a[9] & b[292])^(a[8] & b[293])^(a[7] & b[294])^(a[6] & b[295])^(a[5] & b[296])^(a[4] & b[297])^(a[3] & b[298])^(a[2] & b[299])^(a[1] & b[300])^(a[0] & b[301]);
assign y[302] = (a[302] & b[0])^(a[301] & b[1])^(a[300] & b[2])^(a[299] & b[3])^(a[298] & b[4])^(a[297] & b[5])^(a[296] & b[6])^(a[295] & b[7])^(a[294] & b[8])^(a[293] & b[9])^(a[292] & b[10])^(a[291] & b[11])^(a[290] & b[12])^(a[289] & b[13])^(a[288] & b[14])^(a[287] & b[15])^(a[286] & b[16])^(a[285] & b[17])^(a[284] & b[18])^(a[283] & b[19])^(a[282] & b[20])^(a[281] & b[21])^(a[280] & b[22])^(a[279] & b[23])^(a[278] & b[24])^(a[277] & b[25])^(a[276] & b[26])^(a[275] & b[27])^(a[274] & b[28])^(a[273] & b[29])^(a[272] & b[30])^(a[271] & b[31])^(a[270] & b[32])^(a[269] & b[33])^(a[268] & b[34])^(a[267] & b[35])^(a[266] & b[36])^(a[265] & b[37])^(a[264] & b[38])^(a[263] & b[39])^(a[262] & b[40])^(a[261] & b[41])^(a[260] & b[42])^(a[259] & b[43])^(a[258] & b[44])^(a[257] & b[45])^(a[256] & b[46])^(a[255] & b[47])^(a[254] & b[48])^(a[253] & b[49])^(a[252] & b[50])^(a[251] & b[51])^(a[250] & b[52])^(a[249] & b[53])^(a[248] & b[54])^(a[247] & b[55])^(a[246] & b[56])^(a[245] & b[57])^(a[244] & b[58])^(a[243] & b[59])^(a[242] & b[60])^(a[241] & b[61])^(a[240] & b[62])^(a[239] & b[63])^(a[238] & b[64])^(a[237] & b[65])^(a[236] & b[66])^(a[235] & b[67])^(a[234] & b[68])^(a[233] & b[69])^(a[232] & b[70])^(a[231] & b[71])^(a[230] & b[72])^(a[229] & b[73])^(a[228] & b[74])^(a[227] & b[75])^(a[226] & b[76])^(a[225] & b[77])^(a[224] & b[78])^(a[223] & b[79])^(a[222] & b[80])^(a[221] & b[81])^(a[220] & b[82])^(a[219] & b[83])^(a[218] & b[84])^(a[217] & b[85])^(a[216] & b[86])^(a[215] & b[87])^(a[214] & b[88])^(a[213] & b[89])^(a[212] & b[90])^(a[211] & b[91])^(a[210] & b[92])^(a[209] & b[93])^(a[208] & b[94])^(a[207] & b[95])^(a[206] & b[96])^(a[205] & b[97])^(a[204] & b[98])^(a[203] & b[99])^(a[202] & b[100])^(a[201] & b[101])^(a[200] & b[102])^(a[199] & b[103])^(a[198] & b[104])^(a[197] & b[105])^(a[196] & b[106])^(a[195] & b[107])^(a[194] & b[108])^(a[193] & b[109])^(a[192] & b[110])^(a[191] & b[111])^(a[190] & b[112])^(a[189] & b[113])^(a[188] & b[114])^(a[187] & b[115])^(a[186] & b[116])^(a[185] & b[117])^(a[184] & b[118])^(a[183] & b[119])^(a[182] & b[120])^(a[181] & b[121])^(a[180] & b[122])^(a[179] & b[123])^(a[178] & b[124])^(a[177] & b[125])^(a[176] & b[126])^(a[175] & b[127])^(a[174] & b[128])^(a[173] & b[129])^(a[172] & b[130])^(a[171] & b[131])^(a[170] & b[132])^(a[169] & b[133])^(a[168] & b[134])^(a[167] & b[135])^(a[166] & b[136])^(a[165] & b[137])^(a[164] & b[138])^(a[163] & b[139])^(a[162] & b[140])^(a[161] & b[141])^(a[160] & b[142])^(a[159] & b[143])^(a[158] & b[144])^(a[157] & b[145])^(a[156] & b[146])^(a[155] & b[147])^(a[154] & b[148])^(a[153] & b[149])^(a[152] & b[150])^(a[151] & b[151])^(a[150] & b[152])^(a[149] & b[153])^(a[148] & b[154])^(a[147] & b[155])^(a[146] & b[156])^(a[145] & b[157])^(a[144] & b[158])^(a[143] & b[159])^(a[142] & b[160])^(a[141] & b[161])^(a[140] & b[162])^(a[139] & b[163])^(a[138] & b[164])^(a[137] & b[165])^(a[136] & b[166])^(a[135] & b[167])^(a[134] & b[168])^(a[133] & b[169])^(a[132] & b[170])^(a[131] & b[171])^(a[130] & b[172])^(a[129] & b[173])^(a[128] & b[174])^(a[127] & b[175])^(a[126] & b[176])^(a[125] & b[177])^(a[124] & b[178])^(a[123] & b[179])^(a[122] & b[180])^(a[121] & b[181])^(a[120] & b[182])^(a[119] & b[183])^(a[118] & b[184])^(a[117] & b[185])^(a[116] & b[186])^(a[115] & b[187])^(a[114] & b[188])^(a[113] & b[189])^(a[112] & b[190])^(a[111] & b[191])^(a[110] & b[192])^(a[109] & b[193])^(a[108] & b[194])^(a[107] & b[195])^(a[106] & b[196])^(a[105] & b[197])^(a[104] & b[198])^(a[103] & b[199])^(a[102] & b[200])^(a[101] & b[201])^(a[100] & b[202])^(a[99] & b[203])^(a[98] & b[204])^(a[97] & b[205])^(a[96] & b[206])^(a[95] & b[207])^(a[94] & b[208])^(a[93] & b[209])^(a[92] & b[210])^(a[91] & b[211])^(a[90] & b[212])^(a[89] & b[213])^(a[88] & b[214])^(a[87] & b[215])^(a[86] & b[216])^(a[85] & b[217])^(a[84] & b[218])^(a[83] & b[219])^(a[82] & b[220])^(a[81] & b[221])^(a[80] & b[222])^(a[79] & b[223])^(a[78] & b[224])^(a[77] & b[225])^(a[76] & b[226])^(a[75] & b[227])^(a[74] & b[228])^(a[73] & b[229])^(a[72] & b[230])^(a[71] & b[231])^(a[70] & b[232])^(a[69] & b[233])^(a[68] & b[234])^(a[67] & b[235])^(a[66] & b[236])^(a[65] & b[237])^(a[64] & b[238])^(a[63] & b[239])^(a[62] & b[240])^(a[61] & b[241])^(a[60] & b[242])^(a[59] & b[243])^(a[58] & b[244])^(a[57] & b[245])^(a[56] & b[246])^(a[55] & b[247])^(a[54] & b[248])^(a[53] & b[249])^(a[52] & b[250])^(a[51] & b[251])^(a[50] & b[252])^(a[49] & b[253])^(a[48] & b[254])^(a[47] & b[255])^(a[46] & b[256])^(a[45] & b[257])^(a[44] & b[258])^(a[43] & b[259])^(a[42] & b[260])^(a[41] & b[261])^(a[40] & b[262])^(a[39] & b[263])^(a[38] & b[264])^(a[37] & b[265])^(a[36] & b[266])^(a[35] & b[267])^(a[34] & b[268])^(a[33] & b[269])^(a[32] & b[270])^(a[31] & b[271])^(a[30] & b[272])^(a[29] & b[273])^(a[28] & b[274])^(a[27] & b[275])^(a[26] & b[276])^(a[25] & b[277])^(a[24] & b[278])^(a[23] & b[279])^(a[22] & b[280])^(a[21] & b[281])^(a[20] & b[282])^(a[19] & b[283])^(a[18] & b[284])^(a[17] & b[285])^(a[16] & b[286])^(a[15] & b[287])^(a[14] & b[288])^(a[13] & b[289])^(a[12] & b[290])^(a[11] & b[291])^(a[10] & b[292])^(a[9] & b[293])^(a[8] & b[294])^(a[7] & b[295])^(a[6] & b[296])^(a[5] & b[297])^(a[4] & b[298])^(a[3] & b[299])^(a[2] & b[300])^(a[1] & b[301])^(a[0] & b[302]);
assign y[303] = (a[303] & b[0])^(a[302] & b[1])^(a[301] & b[2])^(a[300] & b[3])^(a[299] & b[4])^(a[298] & b[5])^(a[297] & b[6])^(a[296] & b[7])^(a[295] & b[8])^(a[294] & b[9])^(a[293] & b[10])^(a[292] & b[11])^(a[291] & b[12])^(a[290] & b[13])^(a[289] & b[14])^(a[288] & b[15])^(a[287] & b[16])^(a[286] & b[17])^(a[285] & b[18])^(a[284] & b[19])^(a[283] & b[20])^(a[282] & b[21])^(a[281] & b[22])^(a[280] & b[23])^(a[279] & b[24])^(a[278] & b[25])^(a[277] & b[26])^(a[276] & b[27])^(a[275] & b[28])^(a[274] & b[29])^(a[273] & b[30])^(a[272] & b[31])^(a[271] & b[32])^(a[270] & b[33])^(a[269] & b[34])^(a[268] & b[35])^(a[267] & b[36])^(a[266] & b[37])^(a[265] & b[38])^(a[264] & b[39])^(a[263] & b[40])^(a[262] & b[41])^(a[261] & b[42])^(a[260] & b[43])^(a[259] & b[44])^(a[258] & b[45])^(a[257] & b[46])^(a[256] & b[47])^(a[255] & b[48])^(a[254] & b[49])^(a[253] & b[50])^(a[252] & b[51])^(a[251] & b[52])^(a[250] & b[53])^(a[249] & b[54])^(a[248] & b[55])^(a[247] & b[56])^(a[246] & b[57])^(a[245] & b[58])^(a[244] & b[59])^(a[243] & b[60])^(a[242] & b[61])^(a[241] & b[62])^(a[240] & b[63])^(a[239] & b[64])^(a[238] & b[65])^(a[237] & b[66])^(a[236] & b[67])^(a[235] & b[68])^(a[234] & b[69])^(a[233] & b[70])^(a[232] & b[71])^(a[231] & b[72])^(a[230] & b[73])^(a[229] & b[74])^(a[228] & b[75])^(a[227] & b[76])^(a[226] & b[77])^(a[225] & b[78])^(a[224] & b[79])^(a[223] & b[80])^(a[222] & b[81])^(a[221] & b[82])^(a[220] & b[83])^(a[219] & b[84])^(a[218] & b[85])^(a[217] & b[86])^(a[216] & b[87])^(a[215] & b[88])^(a[214] & b[89])^(a[213] & b[90])^(a[212] & b[91])^(a[211] & b[92])^(a[210] & b[93])^(a[209] & b[94])^(a[208] & b[95])^(a[207] & b[96])^(a[206] & b[97])^(a[205] & b[98])^(a[204] & b[99])^(a[203] & b[100])^(a[202] & b[101])^(a[201] & b[102])^(a[200] & b[103])^(a[199] & b[104])^(a[198] & b[105])^(a[197] & b[106])^(a[196] & b[107])^(a[195] & b[108])^(a[194] & b[109])^(a[193] & b[110])^(a[192] & b[111])^(a[191] & b[112])^(a[190] & b[113])^(a[189] & b[114])^(a[188] & b[115])^(a[187] & b[116])^(a[186] & b[117])^(a[185] & b[118])^(a[184] & b[119])^(a[183] & b[120])^(a[182] & b[121])^(a[181] & b[122])^(a[180] & b[123])^(a[179] & b[124])^(a[178] & b[125])^(a[177] & b[126])^(a[176] & b[127])^(a[175] & b[128])^(a[174] & b[129])^(a[173] & b[130])^(a[172] & b[131])^(a[171] & b[132])^(a[170] & b[133])^(a[169] & b[134])^(a[168] & b[135])^(a[167] & b[136])^(a[166] & b[137])^(a[165] & b[138])^(a[164] & b[139])^(a[163] & b[140])^(a[162] & b[141])^(a[161] & b[142])^(a[160] & b[143])^(a[159] & b[144])^(a[158] & b[145])^(a[157] & b[146])^(a[156] & b[147])^(a[155] & b[148])^(a[154] & b[149])^(a[153] & b[150])^(a[152] & b[151])^(a[151] & b[152])^(a[150] & b[153])^(a[149] & b[154])^(a[148] & b[155])^(a[147] & b[156])^(a[146] & b[157])^(a[145] & b[158])^(a[144] & b[159])^(a[143] & b[160])^(a[142] & b[161])^(a[141] & b[162])^(a[140] & b[163])^(a[139] & b[164])^(a[138] & b[165])^(a[137] & b[166])^(a[136] & b[167])^(a[135] & b[168])^(a[134] & b[169])^(a[133] & b[170])^(a[132] & b[171])^(a[131] & b[172])^(a[130] & b[173])^(a[129] & b[174])^(a[128] & b[175])^(a[127] & b[176])^(a[126] & b[177])^(a[125] & b[178])^(a[124] & b[179])^(a[123] & b[180])^(a[122] & b[181])^(a[121] & b[182])^(a[120] & b[183])^(a[119] & b[184])^(a[118] & b[185])^(a[117] & b[186])^(a[116] & b[187])^(a[115] & b[188])^(a[114] & b[189])^(a[113] & b[190])^(a[112] & b[191])^(a[111] & b[192])^(a[110] & b[193])^(a[109] & b[194])^(a[108] & b[195])^(a[107] & b[196])^(a[106] & b[197])^(a[105] & b[198])^(a[104] & b[199])^(a[103] & b[200])^(a[102] & b[201])^(a[101] & b[202])^(a[100] & b[203])^(a[99] & b[204])^(a[98] & b[205])^(a[97] & b[206])^(a[96] & b[207])^(a[95] & b[208])^(a[94] & b[209])^(a[93] & b[210])^(a[92] & b[211])^(a[91] & b[212])^(a[90] & b[213])^(a[89] & b[214])^(a[88] & b[215])^(a[87] & b[216])^(a[86] & b[217])^(a[85] & b[218])^(a[84] & b[219])^(a[83] & b[220])^(a[82] & b[221])^(a[81] & b[222])^(a[80] & b[223])^(a[79] & b[224])^(a[78] & b[225])^(a[77] & b[226])^(a[76] & b[227])^(a[75] & b[228])^(a[74] & b[229])^(a[73] & b[230])^(a[72] & b[231])^(a[71] & b[232])^(a[70] & b[233])^(a[69] & b[234])^(a[68] & b[235])^(a[67] & b[236])^(a[66] & b[237])^(a[65] & b[238])^(a[64] & b[239])^(a[63] & b[240])^(a[62] & b[241])^(a[61] & b[242])^(a[60] & b[243])^(a[59] & b[244])^(a[58] & b[245])^(a[57] & b[246])^(a[56] & b[247])^(a[55] & b[248])^(a[54] & b[249])^(a[53] & b[250])^(a[52] & b[251])^(a[51] & b[252])^(a[50] & b[253])^(a[49] & b[254])^(a[48] & b[255])^(a[47] & b[256])^(a[46] & b[257])^(a[45] & b[258])^(a[44] & b[259])^(a[43] & b[260])^(a[42] & b[261])^(a[41] & b[262])^(a[40] & b[263])^(a[39] & b[264])^(a[38] & b[265])^(a[37] & b[266])^(a[36] & b[267])^(a[35] & b[268])^(a[34] & b[269])^(a[33] & b[270])^(a[32] & b[271])^(a[31] & b[272])^(a[30] & b[273])^(a[29] & b[274])^(a[28] & b[275])^(a[27] & b[276])^(a[26] & b[277])^(a[25] & b[278])^(a[24] & b[279])^(a[23] & b[280])^(a[22] & b[281])^(a[21] & b[282])^(a[20] & b[283])^(a[19] & b[284])^(a[18] & b[285])^(a[17] & b[286])^(a[16] & b[287])^(a[15] & b[288])^(a[14] & b[289])^(a[13] & b[290])^(a[12] & b[291])^(a[11] & b[292])^(a[10] & b[293])^(a[9] & b[294])^(a[8] & b[295])^(a[7] & b[296])^(a[6] & b[297])^(a[5] & b[298])^(a[4] & b[299])^(a[3] & b[300])^(a[2] & b[301])^(a[1] & b[302])^(a[0] & b[303]);
assign y[304] = (a[304] & b[0])^(a[303] & b[1])^(a[302] & b[2])^(a[301] & b[3])^(a[300] & b[4])^(a[299] & b[5])^(a[298] & b[6])^(a[297] & b[7])^(a[296] & b[8])^(a[295] & b[9])^(a[294] & b[10])^(a[293] & b[11])^(a[292] & b[12])^(a[291] & b[13])^(a[290] & b[14])^(a[289] & b[15])^(a[288] & b[16])^(a[287] & b[17])^(a[286] & b[18])^(a[285] & b[19])^(a[284] & b[20])^(a[283] & b[21])^(a[282] & b[22])^(a[281] & b[23])^(a[280] & b[24])^(a[279] & b[25])^(a[278] & b[26])^(a[277] & b[27])^(a[276] & b[28])^(a[275] & b[29])^(a[274] & b[30])^(a[273] & b[31])^(a[272] & b[32])^(a[271] & b[33])^(a[270] & b[34])^(a[269] & b[35])^(a[268] & b[36])^(a[267] & b[37])^(a[266] & b[38])^(a[265] & b[39])^(a[264] & b[40])^(a[263] & b[41])^(a[262] & b[42])^(a[261] & b[43])^(a[260] & b[44])^(a[259] & b[45])^(a[258] & b[46])^(a[257] & b[47])^(a[256] & b[48])^(a[255] & b[49])^(a[254] & b[50])^(a[253] & b[51])^(a[252] & b[52])^(a[251] & b[53])^(a[250] & b[54])^(a[249] & b[55])^(a[248] & b[56])^(a[247] & b[57])^(a[246] & b[58])^(a[245] & b[59])^(a[244] & b[60])^(a[243] & b[61])^(a[242] & b[62])^(a[241] & b[63])^(a[240] & b[64])^(a[239] & b[65])^(a[238] & b[66])^(a[237] & b[67])^(a[236] & b[68])^(a[235] & b[69])^(a[234] & b[70])^(a[233] & b[71])^(a[232] & b[72])^(a[231] & b[73])^(a[230] & b[74])^(a[229] & b[75])^(a[228] & b[76])^(a[227] & b[77])^(a[226] & b[78])^(a[225] & b[79])^(a[224] & b[80])^(a[223] & b[81])^(a[222] & b[82])^(a[221] & b[83])^(a[220] & b[84])^(a[219] & b[85])^(a[218] & b[86])^(a[217] & b[87])^(a[216] & b[88])^(a[215] & b[89])^(a[214] & b[90])^(a[213] & b[91])^(a[212] & b[92])^(a[211] & b[93])^(a[210] & b[94])^(a[209] & b[95])^(a[208] & b[96])^(a[207] & b[97])^(a[206] & b[98])^(a[205] & b[99])^(a[204] & b[100])^(a[203] & b[101])^(a[202] & b[102])^(a[201] & b[103])^(a[200] & b[104])^(a[199] & b[105])^(a[198] & b[106])^(a[197] & b[107])^(a[196] & b[108])^(a[195] & b[109])^(a[194] & b[110])^(a[193] & b[111])^(a[192] & b[112])^(a[191] & b[113])^(a[190] & b[114])^(a[189] & b[115])^(a[188] & b[116])^(a[187] & b[117])^(a[186] & b[118])^(a[185] & b[119])^(a[184] & b[120])^(a[183] & b[121])^(a[182] & b[122])^(a[181] & b[123])^(a[180] & b[124])^(a[179] & b[125])^(a[178] & b[126])^(a[177] & b[127])^(a[176] & b[128])^(a[175] & b[129])^(a[174] & b[130])^(a[173] & b[131])^(a[172] & b[132])^(a[171] & b[133])^(a[170] & b[134])^(a[169] & b[135])^(a[168] & b[136])^(a[167] & b[137])^(a[166] & b[138])^(a[165] & b[139])^(a[164] & b[140])^(a[163] & b[141])^(a[162] & b[142])^(a[161] & b[143])^(a[160] & b[144])^(a[159] & b[145])^(a[158] & b[146])^(a[157] & b[147])^(a[156] & b[148])^(a[155] & b[149])^(a[154] & b[150])^(a[153] & b[151])^(a[152] & b[152])^(a[151] & b[153])^(a[150] & b[154])^(a[149] & b[155])^(a[148] & b[156])^(a[147] & b[157])^(a[146] & b[158])^(a[145] & b[159])^(a[144] & b[160])^(a[143] & b[161])^(a[142] & b[162])^(a[141] & b[163])^(a[140] & b[164])^(a[139] & b[165])^(a[138] & b[166])^(a[137] & b[167])^(a[136] & b[168])^(a[135] & b[169])^(a[134] & b[170])^(a[133] & b[171])^(a[132] & b[172])^(a[131] & b[173])^(a[130] & b[174])^(a[129] & b[175])^(a[128] & b[176])^(a[127] & b[177])^(a[126] & b[178])^(a[125] & b[179])^(a[124] & b[180])^(a[123] & b[181])^(a[122] & b[182])^(a[121] & b[183])^(a[120] & b[184])^(a[119] & b[185])^(a[118] & b[186])^(a[117] & b[187])^(a[116] & b[188])^(a[115] & b[189])^(a[114] & b[190])^(a[113] & b[191])^(a[112] & b[192])^(a[111] & b[193])^(a[110] & b[194])^(a[109] & b[195])^(a[108] & b[196])^(a[107] & b[197])^(a[106] & b[198])^(a[105] & b[199])^(a[104] & b[200])^(a[103] & b[201])^(a[102] & b[202])^(a[101] & b[203])^(a[100] & b[204])^(a[99] & b[205])^(a[98] & b[206])^(a[97] & b[207])^(a[96] & b[208])^(a[95] & b[209])^(a[94] & b[210])^(a[93] & b[211])^(a[92] & b[212])^(a[91] & b[213])^(a[90] & b[214])^(a[89] & b[215])^(a[88] & b[216])^(a[87] & b[217])^(a[86] & b[218])^(a[85] & b[219])^(a[84] & b[220])^(a[83] & b[221])^(a[82] & b[222])^(a[81] & b[223])^(a[80] & b[224])^(a[79] & b[225])^(a[78] & b[226])^(a[77] & b[227])^(a[76] & b[228])^(a[75] & b[229])^(a[74] & b[230])^(a[73] & b[231])^(a[72] & b[232])^(a[71] & b[233])^(a[70] & b[234])^(a[69] & b[235])^(a[68] & b[236])^(a[67] & b[237])^(a[66] & b[238])^(a[65] & b[239])^(a[64] & b[240])^(a[63] & b[241])^(a[62] & b[242])^(a[61] & b[243])^(a[60] & b[244])^(a[59] & b[245])^(a[58] & b[246])^(a[57] & b[247])^(a[56] & b[248])^(a[55] & b[249])^(a[54] & b[250])^(a[53] & b[251])^(a[52] & b[252])^(a[51] & b[253])^(a[50] & b[254])^(a[49] & b[255])^(a[48] & b[256])^(a[47] & b[257])^(a[46] & b[258])^(a[45] & b[259])^(a[44] & b[260])^(a[43] & b[261])^(a[42] & b[262])^(a[41] & b[263])^(a[40] & b[264])^(a[39] & b[265])^(a[38] & b[266])^(a[37] & b[267])^(a[36] & b[268])^(a[35] & b[269])^(a[34] & b[270])^(a[33] & b[271])^(a[32] & b[272])^(a[31] & b[273])^(a[30] & b[274])^(a[29] & b[275])^(a[28] & b[276])^(a[27] & b[277])^(a[26] & b[278])^(a[25] & b[279])^(a[24] & b[280])^(a[23] & b[281])^(a[22] & b[282])^(a[21] & b[283])^(a[20] & b[284])^(a[19] & b[285])^(a[18] & b[286])^(a[17] & b[287])^(a[16] & b[288])^(a[15] & b[289])^(a[14] & b[290])^(a[13] & b[291])^(a[12] & b[292])^(a[11] & b[293])^(a[10] & b[294])^(a[9] & b[295])^(a[8] & b[296])^(a[7] & b[297])^(a[6] & b[298])^(a[5] & b[299])^(a[4] & b[300])^(a[3] & b[301])^(a[2] & b[302])^(a[1] & b[303])^(a[0] & b[304]);
assign y[305] = (a[305] & b[0])^(a[304] & b[1])^(a[303] & b[2])^(a[302] & b[3])^(a[301] & b[4])^(a[300] & b[5])^(a[299] & b[6])^(a[298] & b[7])^(a[297] & b[8])^(a[296] & b[9])^(a[295] & b[10])^(a[294] & b[11])^(a[293] & b[12])^(a[292] & b[13])^(a[291] & b[14])^(a[290] & b[15])^(a[289] & b[16])^(a[288] & b[17])^(a[287] & b[18])^(a[286] & b[19])^(a[285] & b[20])^(a[284] & b[21])^(a[283] & b[22])^(a[282] & b[23])^(a[281] & b[24])^(a[280] & b[25])^(a[279] & b[26])^(a[278] & b[27])^(a[277] & b[28])^(a[276] & b[29])^(a[275] & b[30])^(a[274] & b[31])^(a[273] & b[32])^(a[272] & b[33])^(a[271] & b[34])^(a[270] & b[35])^(a[269] & b[36])^(a[268] & b[37])^(a[267] & b[38])^(a[266] & b[39])^(a[265] & b[40])^(a[264] & b[41])^(a[263] & b[42])^(a[262] & b[43])^(a[261] & b[44])^(a[260] & b[45])^(a[259] & b[46])^(a[258] & b[47])^(a[257] & b[48])^(a[256] & b[49])^(a[255] & b[50])^(a[254] & b[51])^(a[253] & b[52])^(a[252] & b[53])^(a[251] & b[54])^(a[250] & b[55])^(a[249] & b[56])^(a[248] & b[57])^(a[247] & b[58])^(a[246] & b[59])^(a[245] & b[60])^(a[244] & b[61])^(a[243] & b[62])^(a[242] & b[63])^(a[241] & b[64])^(a[240] & b[65])^(a[239] & b[66])^(a[238] & b[67])^(a[237] & b[68])^(a[236] & b[69])^(a[235] & b[70])^(a[234] & b[71])^(a[233] & b[72])^(a[232] & b[73])^(a[231] & b[74])^(a[230] & b[75])^(a[229] & b[76])^(a[228] & b[77])^(a[227] & b[78])^(a[226] & b[79])^(a[225] & b[80])^(a[224] & b[81])^(a[223] & b[82])^(a[222] & b[83])^(a[221] & b[84])^(a[220] & b[85])^(a[219] & b[86])^(a[218] & b[87])^(a[217] & b[88])^(a[216] & b[89])^(a[215] & b[90])^(a[214] & b[91])^(a[213] & b[92])^(a[212] & b[93])^(a[211] & b[94])^(a[210] & b[95])^(a[209] & b[96])^(a[208] & b[97])^(a[207] & b[98])^(a[206] & b[99])^(a[205] & b[100])^(a[204] & b[101])^(a[203] & b[102])^(a[202] & b[103])^(a[201] & b[104])^(a[200] & b[105])^(a[199] & b[106])^(a[198] & b[107])^(a[197] & b[108])^(a[196] & b[109])^(a[195] & b[110])^(a[194] & b[111])^(a[193] & b[112])^(a[192] & b[113])^(a[191] & b[114])^(a[190] & b[115])^(a[189] & b[116])^(a[188] & b[117])^(a[187] & b[118])^(a[186] & b[119])^(a[185] & b[120])^(a[184] & b[121])^(a[183] & b[122])^(a[182] & b[123])^(a[181] & b[124])^(a[180] & b[125])^(a[179] & b[126])^(a[178] & b[127])^(a[177] & b[128])^(a[176] & b[129])^(a[175] & b[130])^(a[174] & b[131])^(a[173] & b[132])^(a[172] & b[133])^(a[171] & b[134])^(a[170] & b[135])^(a[169] & b[136])^(a[168] & b[137])^(a[167] & b[138])^(a[166] & b[139])^(a[165] & b[140])^(a[164] & b[141])^(a[163] & b[142])^(a[162] & b[143])^(a[161] & b[144])^(a[160] & b[145])^(a[159] & b[146])^(a[158] & b[147])^(a[157] & b[148])^(a[156] & b[149])^(a[155] & b[150])^(a[154] & b[151])^(a[153] & b[152])^(a[152] & b[153])^(a[151] & b[154])^(a[150] & b[155])^(a[149] & b[156])^(a[148] & b[157])^(a[147] & b[158])^(a[146] & b[159])^(a[145] & b[160])^(a[144] & b[161])^(a[143] & b[162])^(a[142] & b[163])^(a[141] & b[164])^(a[140] & b[165])^(a[139] & b[166])^(a[138] & b[167])^(a[137] & b[168])^(a[136] & b[169])^(a[135] & b[170])^(a[134] & b[171])^(a[133] & b[172])^(a[132] & b[173])^(a[131] & b[174])^(a[130] & b[175])^(a[129] & b[176])^(a[128] & b[177])^(a[127] & b[178])^(a[126] & b[179])^(a[125] & b[180])^(a[124] & b[181])^(a[123] & b[182])^(a[122] & b[183])^(a[121] & b[184])^(a[120] & b[185])^(a[119] & b[186])^(a[118] & b[187])^(a[117] & b[188])^(a[116] & b[189])^(a[115] & b[190])^(a[114] & b[191])^(a[113] & b[192])^(a[112] & b[193])^(a[111] & b[194])^(a[110] & b[195])^(a[109] & b[196])^(a[108] & b[197])^(a[107] & b[198])^(a[106] & b[199])^(a[105] & b[200])^(a[104] & b[201])^(a[103] & b[202])^(a[102] & b[203])^(a[101] & b[204])^(a[100] & b[205])^(a[99] & b[206])^(a[98] & b[207])^(a[97] & b[208])^(a[96] & b[209])^(a[95] & b[210])^(a[94] & b[211])^(a[93] & b[212])^(a[92] & b[213])^(a[91] & b[214])^(a[90] & b[215])^(a[89] & b[216])^(a[88] & b[217])^(a[87] & b[218])^(a[86] & b[219])^(a[85] & b[220])^(a[84] & b[221])^(a[83] & b[222])^(a[82] & b[223])^(a[81] & b[224])^(a[80] & b[225])^(a[79] & b[226])^(a[78] & b[227])^(a[77] & b[228])^(a[76] & b[229])^(a[75] & b[230])^(a[74] & b[231])^(a[73] & b[232])^(a[72] & b[233])^(a[71] & b[234])^(a[70] & b[235])^(a[69] & b[236])^(a[68] & b[237])^(a[67] & b[238])^(a[66] & b[239])^(a[65] & b[240])^(a[64] & b[241])^(a[63] & b[242])^(a[62] & b[243])^(a[61] & b[244])^(a[60] & b[245])^(a[59] & b[246])^(a[58] & b[247])^(a[57] & b[248])^(a[56] & b[249])^(a[55] & b[250])^(a[54] & b[251])^(a[53] & b[252])^(a[52] & b[253])^(a[51] & b[254])^(a[50] & b[255])^(a[49] & b[256])^(a[48] & b[257])^(a[47] & b[258])^(a[46] & b[259])^(a[45] & b[260])^(a[44] & b[261])^(a[43] & b[262])^(a[42] & b[263])^(a[41] & b[264])^(a[40] & b[265])^(a[39] & b[266])^(a[38] & b[267])^(a[37] & b[268])^(a[36] & b[269])^(a[35] & b[270])^(a[34] & b[271])^(a[33] & b[272])^(a[32] & b[273])^(a[31] & b[274])^(a[30] & b[275])^(a[29] & b[276])^(a[28] & b[277])^(a[27] & b[278])^(a[26] & b[279])^(a[25] & b[280])^(a[24] & b[281])^(a[23] & b[282])^(a[22] & b[283])^(a[21] & b[284])^(a[20] & b[285])^(a[19] & b[286])^(a[18] & b[287])^(a[17] & b[288])^(a[16] & b[289])^(a[15] & b[290])^(a[14] & b[291])^(a[13] & b[292])^(a[12] & b[293])^(a[11] & b[294])^(a[10] & b[295])^(a[9] & b[296])^(a[8] & b[297])^(a[7] & b[298])^(a[6] & b[299])^(a[5] & b[300])^(a[4] & b[301])^(a[3] & b[302])^(a[2] & b[303])^(a[1] & b[304])^(a[0] & b[305]);
assign y[306] = (a[306] & b[0])^(a[305] & b[1])^(a[304] & b[2])^(a[303] & b[3])^(a[302] & b[4])^(a[301] & b[5])^(a[300] & b[6])^(a[299] & b[7])^(a[298] & b[8])^(a[297] & b[9])^(a[296] & b[10])^(a[295] & b[11])^(a[294] & b[12])^(a[293] & b[13])^(a[292] & b[14])^(a[291] & b[15])^(a[290] & b[16])^(a[289] & b[17])^(a[288] & b[18])^(a[287] & b[19])^(a[286] & b[20])^(a[285] & b[21])^(a[284] & b[22])^(a[283] & b[23])^(a[282] & b[24])^(a[281] & b[25])^(a[280] & b[26])^(a[279] & b[27])^(a[278] & b[28])^(a[277] & b[29])^(a[276] & b[30])^(a[275] & b[31])^(a[274] & b[32])^(a[273] & b[33])^(a[272] & b[34])^(a[271] & b[35])^(a[270] & b[36])^(a[269] & b[37])^(a[268] & b[38])^(a[267] & b[39])^(a[266] & b[40])^(a[265] & b[41])^(a[264] & b[42])^(a[263] & b[43])^(a[262] & b[44])^(a[261] & b[45])^(a[260] & b[46])^(a[259] & b[47])^(a[258] & b[48])^(a[257] & b[49])^(a[256] & b[50])^(a[255] & b[51])^(a[254] & b[52])^(a[253] & b[53])^(a[252] & b[54])^(a[251] & b[55])^(a[250] & b[56])^(a[249] & b[57])^(a[248] & b[58])^(a[247] & b[59])^(a[246] & b[60])^(a[245] & b[61])^(a[244] & b[62])^(a[243] & b[63])^(a[242] & b[64])^(a[241] & b[65])^(a[240] & b[66])^(a[239] & b[67])^(a[238] & b[68])^(a[237] & b[69])^(a[236] & b[70])^(a[235] & b[71])^(a[234] & b[72])^(a[233] & b[73])^(a[232] & b[74])^(a[231] & b[75])^(a[230] & b[76])^(a[229] & b[77])^(a[228] & b[78])^(a[227] & b[79])^(a[226] & b[80])^(a[225] & b[81])^(a[224] & b[82])^(a[223] & b[83])^(a[222] & b[84])^(a[221] & b[85])^(a[220] & b[86])^(a[219] & b[87])^(a[218] & b[88])^(a[217] & b[89])^(a[216] & b[90])^(a[215] & b[91])^(a[214] & b[92])^(a[213] & b[93])^(a[212] & b[94])^(a[211] & b[95])^(a[210] & b[96])^(a[209] & b[97])^(a[208] & b[98])^(a[207] & b[99])^(a[206] & b[100])^(a[205] & b[101])^(a[204] & b[102])^(a[203] & b[103])^(a[202] & b[104])^(a[201] & b[105])^(a[200] & b[106])^(a[199] & b[107])^(a[198] & b[108])^(a[197] & b[109])^(a[196] & b[110])^(a[195] & b[111])^(a[194] & b[112])^(a[193] & b[113])^(a[192] & b[114])^(a[191] & b[115])^(a[190] & b[116])^(a[189] & b[117])^(a[188] & b[118])^(a[187] & b[119])^(a[186] & b[120])^(a[185] & b[121])^(a[184] & b[122])^(a[183] & b[123])^(a[182] & b[124])^(a[181] & b[125])^(a[180] & b[126])^(a[179] & b[127])^(a[178] & b[128])^(a[177] & b[129])^(a[176] & b[130])^(a[175] & b[131])^(a[174] & b[132])^(a[173] & b[133])^(a[172] & b[134])^(a[171] & b[135])^(a[170] & b[136])^(a[169] & b[137])^(a[168] & b[138])^(a[167] & b[139])^(a[166] & b[140])^(a[165] & b[141])^(a[164] & b[142])^(a[163] & b[143])^(a[162] & b[144])^(a[161] & b[145])^(a[160] & b[146])^(a[159] & b[147])^(a[158] & b[148])^(a[157] & b[149])^(a[156] & b[150])^(a[155] & b[151])^(a[154] & b[152])^(a[153] & b[153])^(a[152] & b[154])^(a[151] & b[155])^(a[150] & b[156])^(a[149] & b[157])^(a[148] & b[158])^(a[147] & b[159])^(a[146] & b[160])^(a[145] & b[161])^(a[144] & b[162])^(a[143] & b[163])^(a[142] & b[164])^(a[141] & b[165])^(a[140] & b[166])^(a[139] & b[167])^(a[138] & b[168])^(a[137] & b[169])^(a[136] & b[170])^(a[135] & b[171])^(a[134] & b[172])^(a[133] & b[173])^(a[132] & b[174])^(a[131] & b[175])^(a[130] & b[176])^(a[129] & b[177])^(a[128] & b[178])^(a[127] & b[179])^(a[126] & b[180])^(a[125] & b[181])^(a[124] & b[182])^(a[123] & b[183])^(a[122] & b[184])^(a[121] & b[185])^(a[120] & b[186])^(a[119] & b[187])^(a[118] & b[188])^(a[117] & b[189])^(a[116] & b[190])^(a[115] & b[191])^(a[114] & b[192])^(a[113] & b[193])^(a[112] & b[194])^(a[111] & b[195])^(a[110] & b[196])^(a[109] & b[197])^(a[108] & b[198])^(a[107] & b[199])^(a[106] & b[200])^(a[105] & b[201])^(a[104] & b[202])^(a[103] & b[203])^(a[102] & b[204])^(a[101] & b[205])^(a[100] & b[206])^(a[99] & b[207])^(a[98] & b[208])^(a[97] & b[209])^(a[96] & b[210])^(a[95] & b[211])^(a[94] & b[212])^(a[93] & b[213])^(a[92] & b[214])^(a[91] & b[215])^(a[90] & b[216])^(a[89] & b[217])^(a[88] & b[218])^(a[87] & b[219])^(a[86] & b[220])^(a[85] & b[221])^(a[84] & b[222])^(a[83] & b[223])^(a[82] & b[224])^(a[81] & b[225])^(a[80] & b[226])^(a[79] & b[227])^(a[78] & b[228])^(a[77] & b[229])^(a[76] & b[230])^(a[75] & b[231])^(a[74] & b[232])^(a[73] & b[233])^(a[72] & b[234])^(a[71] & b[235])^(a[70] & b[236])^(a[69] & b[237])^(a[68] & b[238])^(a[67] & b[239])^(a[66] & b[240])^(a[65] & b[241])^(a[64] & b[242])^(a[63] & b[243])^(a[62] & b[244])^(a[61] & b[245])^(a[60] & b[246])^(a[59] & b[247])^(a[58] & b[248])^(a[57] & b[249])^(a[56] & b[250])^(a[55] & b[251])^(a[54] & b[252])^(a[53] & b[253])^(a[52] & b[254])^(a[51] & b[255])^(a[50] & b[256])^(a[49] & b[257])^(a[48] & b[258])^(a[47] & b[259])^(a[46] & b[260])^(a[45] & b[261])^(a[44] & b[262])^(a[43] & b[263])^(a[42] & b[264])^(a[41] & b[265])^(a[40] & b[266])^(a[39] & b[267])^(a[38] & b[268])^(a[37] & b[269])^(a[36] & b[270])^(a[35] & b[271])^(a[34] & b[272])^(a[33] & b[273])^(a[32] & b[274])^(a[31] & b[275])^(a[30] & b[276])^(a[29] & b[277])^(a[28] & b[278])^(a[27] & b[279])^(a[26] & b[280])^(a[25] & b[281])^(a[24] & b[282])^(a[23] & b[283])^(a[22] & b[284])^(a[21] & b[285])^(a[20] & b[286])^(a[19] & b[287])^(a[18] & b[288])^(a[17] & b[289])^(a[16] & b[290])^(a[15] & b[291])^(a[14] & b[292])^(a[13] & b[293])^(a[12] & b[294])^(a[11] & b[295])^(a[10] & b[296])^(a[9] & b[297])^(a[8] & b[298])^(a[7] & b[299])^(a[6] & b[300])^(a[5] & b[301])^(a[4] & b[302])^(a[3] & b[303])^(a[2] & b[304])^(a[1] & b[305])^(a[0] & b[306]);
assign y[307] = (a[307] & b[0])^(a[306] & b[1])^(a[305] & b[2])^(a[304] & b[3])^(a[303] & b[4])^(a[302] & b[5])^(a[301] & b[6])^(a[300] & b[7])^(a[299] & b[8])^(a[298] & b[9])^(a[297] & b[10])^(a[296] & b[11])^(a[295] & b[12])^(a[294] & b[13])^(a[293] & b[14])^(a[292] & b[15])^(a[291] & b[16])^(a[290] & b[17])^(a[289] & b[18])^(a[288] & b[19])^(a[287] & b[20])^(a[286] & b[21])^(a[285] & b[22])^(a[284] & b[23])^(a[283] & b[24])^(a[282] & b[25])^(a[281] & b[26])^(a[280] & b[27])^(a[279] & b[28])^(a[278] & b[29])^(a[277] & b[30])^(a[276] & b[31])^(a[275] & b[32])^(a[274] & b[33])^(a[273] & b[34])^(a[272] & b[35])^(a[271] & b[36])^(a[270] & b[37])^(a[269] & b[38])^(a[268] & b[39])^(a[267] & b[40])^(a[266] & b[41])^(a[265] & b[42])^(a[264] & b[43])^(a[263] & b[44])^(a[262] & b[45])^(a[261] & b[46])^(a[260] & b[47])^(a[259] & b[48])^(a[258] & b[49])^(a[257] & b[50])^(a[256] & b[51])^(a[255] & b[52])^(a[254] & b[53])^(a[253] & b[54])^(a[252] & b[55])^(a[251] & b[56])^(a[250] & b[57])^(a[249] & b[58])^(a[248] & b[59])^(a[247] & b[60])^(a[246] & b[61])^(a[245] & b[62])^(a[244] & b[63])^(a[243] & b[64])^(a[242] & b[65])^(a[241] & b[66])^(a[240] & b[67])^(a[239] & b[68])^(a[238] & b[69])^(a[237] & b[70])^(a[236] & b[71])^(a[235] & b[72])^(a[234] & b[73])^(a[233] & b[74])^(a[232] & b[75])^(a[231] & b[76])^(a[230] & b[77])^(a[229] & b[78])^(a[228] & b[79])^(a[227] & b[80])^(a[226] & b[81])^(a[225] & b[82])^(a[224] & b[83])^(a[223] & b[84])^(a[222] & b[85])^(a[221] & b[86])^(a[220] & b[87])^(a[219] & b[88])^(a[218] & b[89])^(a[217] & b[90])^(a[216] & b[91])^(a[215] & b[92])^(a[214] & b[93])^(a[213] & b[94])^(a[212] & b[95])^(a[211] & b[96])^(a[210] & b[97])^(a[209] & b[98])^(a[208] & b[99])^(a[207] & b[100])^(a[206] & b[101])^(a[205] & b[102])^(a[204] & b[103])^(a[203] & b[104])^(a[202] & b[105])^(a[201] & b[106])^(a[200] & b[107])^(a[199] & b[108])^(a[198] & b[109])^(a[197] & b[110])^(a[196] & b[111])^(a[195] & b[112])^(a[194] & b[113])^(a[193] & b[114])^(a[192] & b[115])^(a[191] & b[116])^(a[190] & b[117])^(a[189] & b[118])^(a[188] & b[119])^(a[187] & b[120])^(a[186] & b[121])^(a[185] & b[122])^(a[184] & b[123])^(a[183] & b[124])^(a[182] & b[125])^(a[181] & b[126])^(a[180] & b[127])^(a[179] & b[128])^(a[178] & b[129])^(a[177] & b[130])^(a[176] & b[131])^(a[175] & b[132])^(a[174] & b[133])^(a[173] & b[134])^(a[172] & b[135])^(a[171] & b[136])^(a[170] & b[137])^(a[169] & b[138])^(a[168] & b[139])^(a[167] & b[140])^(a[166] & b[141])^(a[165] & b[142])^(a[164] & b[143])^(a[163] & b[144])^(a[162] & b[145])^(a[161] & b[146])^(a[160] & b[147])^(a[159] & b[148])^(a[158] & b[149])^(a[157] & b[150])^(a[156] & b[151])^(a[155] & b[152])^(a[154] & b[153])^(a[153] & b[154])^(a[152] & b[155])^(a[151] & b[156])^(a[150] & b[157])^(a[149] & b[158])^(a[148] & b[159])^(a[147] & b[160])^(a[146] & b[161])^(a[145] & b[162])^(a[144] & b[163])^(a[143] & b[164])^(a[142] & b[165])^(a[141] & b[166])^(a[140] & b[167])^(a[139] & b[168])^(a[138] & b[169])^(a[137] & b[170])^(a[136] & b[171])^(a[135] & b[172])^(a[134] & b[173])^(a[133] & b[174])^(a[132] & b[175])^(a[131] & b[176])^(a[130] & b[177])^(a[129] & b[178])^(a[128] & b[179])^(a[127] & b[180])^(a[126] & b[181])^(a[125] & b[182])^(a[124] & b[183])^(a[123] & b[184])^(a[122] & b[185])^(a[121] & b[186])^(a[120] & b[187])^(a[119] & b[188])^(a[118] & b[189])^(a[117] & b[190])^(a[116] & b[191])^(a[115] & b[192])^(a[114] & b[193])^(a[113] & b[194])^(a[112] & b[195])^(a[111] & b[196])^(a[110] & b[197])^(a[109] & b[198])^(a[108] & b[199])^(a[107] & b[200])^(a[106] & b[201])^(a[105] & b[202])^(a[104] & b[203])^(a[103] & b[204])^(a[102] & b[205])^(a[101] & b[206])^(a[100] & b[207])^(a[99] & b[208])^(a[98] & b[209])^(a[97] & b[210])^(a[96] & b[211])^(a[95] & b[212])^(a[94] & b[213])^(a[93] & b[214])^(a[92] & b[215])^(a[91] & b[216])^(a[90] & b[217])^(a[89] & b[218])^(a[88] & b[219])^(a[87] & b[220])^(a[86] & b[221])^(a[85] & b[222])^(a[84] & b[223])^(a[83] & b[224])^(a[82] & b[225])^(a[81] & b[226])^(a[80] & b[227])^(a[79] & b[228])^(a[78] & b[229])^(a[77] & b[230])^(a[76] & b[231])^(a[75] & b[232])^(a[74] & b[233])^(a[73] & b[234])^(a[72] & b[235])^(a[71] & b[236])^(a[70] & b[237])^(a[69] & b[238])^(a[68] & b[239])^(a[67] & b[240])^(a[66] & b[241])^(a[65] & b[242])^(a[64] & b[243])^(a[63] & b[244])^(a[62] & b[245])^(a[61] & b[246])^(a[60] & b[247])^(a[59] & b[248])^(a[58] & b[249])^(a[57] & b[250])^(a[56] & b[251])^(a[55] & b[252])^(a[54] & b[253])^(a[53] & b[254])^(a[52] & b[255])^(a[51] & b[256])^(a[50] & b[257])^(a[49] & b[258])^(a[48] & b[259])^(a[47] & b[260])^(a[46] & b[261])^(a[45] & b[262])^(a[44] & b[263])^(a[43] & b[264])^(a[42] & b[265])^(a[41] & b[266])^(a[40] & b[267])^(a[39] & b[268])^(a[38] & b[269])^(a[37] & b[270])^(a[36] & b[271])^(a[35] & b[272])^(a[34] & b[273])^(a[33] & b[274])^(a[32] & b[275])^(a[31] & b[276])^(a[30] & b[277])^(a[29] & b[278])^(a[28] & b[279])^(a[27] & b[280])^(a[26] & b[281])^(a[25] & b[282])^(a[24] & b[283])^(a[23] & b[284])^(a[22] & b[285])^(a[21] & b[286])^(a[20] & b[287])^(a[19] & b[288])^(a[18] & b[289])^(a[17] & b[290])^(a[16] & b[291])^(a[15] & b[292])^(a[14] & b[293])^(a[13] & b[294])^(a[12] & b[295])^(a[11] & b[296])^(a[10] & b[297])^(a[9] & b[298])^(a[8] & b[299])^(a[7] & b[300])^(a[6] & b[301])^(a[5] & b[302])^(a[4] & b[303])^(a[3] & b[304])^(a[2] & b[305])^(a[1] & b[306])^(a[0] & b[307]);
assign y[308] = (a[308] & b[0])^(a[307] & b[1])^(a[306] & b[2])^(a[305] & b[3])^(a[304] & b[4])^(a[303] & b[5])^(a[302] & b[6])^(a[301] & b[7])^(a[300] & b[8])^(a[299] & b[9])^(a[298] & b[10])^(a[297] & b[11])^(a[296] & b[12])^(a[295] & b[13])^(a[294] & b[14])^(a[293] & b[15])^(a[292] & b[16])^(a[291] & b[17])^(a[290] & b[18])^(a[289] & b[19])^(a[288] & b[20])^(a[287] & b[21])^(a[286] & b[22])^(a[285] & b[23])^(a[284] & b[24])^(a[283] & b[25])^(a[282] & b[26])^(a[281] & b[27])^(a[280] & b[28])^(a[279] & b[29])^(a[278] & b[30])^(a[277] & b[31])^(a[276] & b[32])^(a[275] & b[33])^(a[274] & b[34])^(a[273] & b[35])^(a[272] & b[36])^(a[271] & b[37])^(a[270] & b[38])^(a[269] & b[39])^(a[268] & b[40])^(a[267] & b[41])^(a[266] & b[42])^(a[265] & b[43])^(a[264] & b[44])^(a[263] & b[45])^(a[262] & b[46])^(a[261] & b[47])^(a[260] & b[48])^(a[259] & b[49])^(a[258] & b[50])^(a[257] & b[51])^(a[256] & b[52])^(a[255] & b[53])^(a[254] & b[54])^(a[253] & b[55])^(a[252] & b[56])^(a[251] & b[57])^(a[250] & b[58])^(a[249] & b[59])^(a[248] & b[60])^(a[247] & b[61])^(a[246] & b[62])^(a[245] & b[63])^(a[244] & b[64])^(a[243] & b[65])^(a[242] & b[66])^(a[241] & b[67])^(a[240] & b[68])^(a[239] & b[69])^(a[238] & b[70])^(a[237] & b[71])^(a[236] & b[72])^(a[235] & b[73])^(a[234] & b[74])^(a[233] & b[75])^(a[232] & b[76])^(a[231] & b[77])^(a[230] & b[78])^(a[229] & b[79])^(a[228] & b[80])^(a[227] & b[81])^(a[226] & b[82])^(a[225] & b[83])^(a[224] & b[84])^(a[223] & b[85])^(a[222] & b[86])^(a[221] & b[87])^(a[220] & b[88])^(a[219] & b[89])^(a[218] & b[90])^(a[217] & b[91])^(a[216] & b[92])^(a[215] & b[93])^(a[214] & b[94])^(a[213] & b[95])^(a[212] & b[96])^(a[211] & b[97])^(a[210] & b[98])^(a[209] & b[99])^(a[208] & b[100])^(a[207] & b[101])^(a[206] & b[102])^(a[205] & b[103])^(a[204] & b[104])^(a[203] & b[105])^(a[202] & b[106])^(a[201] & b[107])^(a[200] & b[108])^(a[199] & b[109])^(a[198] & b[110])^(a[197] & b[111])^(a[196] & b[112])^(a[195] & b[113])^(a[194] & b[114])^(a[193] & b[115])^(a[192] & b[116])^(a[191] & b[117])^(a[190] & b[118])^(a[189] & b[119])^(a[188] & b[120])^(a[187] & b[121])^(a[186] & b[122])^(a[185] & b[123])^(a[184] & b[124])^(a[183] & b[125])^(a[182] & b[126])^(a[181] & b[127])^(a[180] & b[128])^(a[179] & b[129])^(a[178] & b[130])^(a[177] & b[131])^(a[176] & b[132])^(a[175] & b[133])^(a[174] & b[134])^(a[173] & b[135])^(a[172] & b[136])^(a[171] & b[137])^(a[170] & b[138])^(a[169] & b[139])^(a[168] & b[140])^(a[167] & b[141])^(a[166] & b[142])^(a[165] & b[143])^(a[164] & b[144])^(a[163] & b[145])^(a[162] & b[146])^(a[161] & b[147])^(a[160] & b[148])^(a[159] & b[149])^(a[158] & b[150])^(a[157] & b[151])^(a[156] & b[152])^(a[155] & b[153])^(a[154] & b[154])^(a[153] & b[155])^(a[152] & b[156])^(a[151] & b[157])^(a[150] & b[158])^(a[149] & b[159])^(a[148] & b[160])^(a[147] & b[161])^(a[146] & b[162])^(a[145] & b[163])^(a[144] & b[164])^(a[143] & b[165])^(a[142] & b[166])^(a[141] & b[167])^(a[140] & b[168])^(a[139] & b[169])^(a[138] & b[170])^(a[137] & b[171])^(a[136] & b[172])^(a[135] & b[173])^(a[134] & b[174])^(a[133] & b[175])^(a[132] & b[176])^(a[131] & b[177])^(a[130] & b[178])^(a[129] & b[179])^(a[128] & b[180])^(a[127] & b[181])^(a[126] & b[182])^(a[125] & b[183])^(a[124] & b[184])^(a[123] & b[185])^(a[122] & b[186])^(a[121] & b[187])^(a[120] & b[188])^(a[119] & b[189])^(a[118] & b[190])^(a[117] & b[191])^(a[116] & b[192])^(a[115] & b[193])^(a[114] & b[194])^(a[113] & b[195])^(a[112] & b[196])^(a[111] & b[197])^(a[110] & b[198])^(a[109] & b[199])^(a[108] & b[200])^(a[107] & b[201])^(a[106] & b[202])^(a[105] & b[203])^(a[104] & b[204])^(a[103] & b[205])^(a[102] & b[206])^(a[101] & b[207])^(a[100] & b[208])^(a[99] & b[209])^(a[98] & b[210])^(a[97] & b[211])^(a[96] & b[212])^(a[95] & b[213])^(a[94] & b[214])^(a[93] & b[215])^(a[92] & b[216])^(a[91] & b[217])^(a[90] & b[218])^(a[89] & b[219])^(a[88] & b[220])^(a[87] & b[221])^(a[86] & b[222])^(a[85] & b[223])^(a[84] & b[224])^(a[83] & b[225])^(a[82] & b[226])^(a[81] & b[227])^(a[80] & b[228])^(a[79] & b[229])^(a[78] & b[230])^(a[77] & b[231])^(a[76] & b[232])^(a[75] & b[233])^(a[74] & b[234])^(a[73] & b[235])^(a[72] & b[236])^(a[71] & b[237])^(a[70] & b[238])^(a[69] & b[239])^(a[68] & b[240])^(a[67] & b[241])^(a[66] & b[242])^(a[65] & b[243])^(a[64] & b[244])^(a[63] & b[245])^(a[62] & b[246])^(a[61] & b[247])^(a[60] & b[248])^(a[59] & b[249])^(a[58] & b[250])^(a[57] & b[251])^(a[56] & b[252])^(a[55] & b[253])^(a[54] & b[254])^(a[53] & b[255])^(a[52] & b[256])^(a[51] & b[257])^(a[50] & b[258])^(a[49] & b[259])^(a[48] & b[260])^(a[47] & b[261])^(a[46] & b[262])^(a[45] & b[263])^(a[44] & b[264])^(a[43] & b[265])^(a[42] & b[266])^(a[41] & b[267])^(a[40] & b[268])^(a[39] & b[269])^(a[38] & b[270])^(a[37] & b[271])^(a[36] & b[272])^(a[35] & b[273])^(a[34] & b[274])^(a[33] & b[275])^(a[32] & b[276])^(a[31] & b[277])^(a[30] & b[278])^(a[29] & b[279])^(a[28] & b[280])^(a[27] & b[281])^(a[26] & b[282])^(a[25] & b[283])^(a[24] & b[284])^(a[23] & b[285])^(a[22] & b[286])^(a[21] & b[287])^(a[20] & b[288])^(a[19] & b[289])^(a[18] & b[290])^(a[17] & b[291])^(a[16] & b[292])^(a[15] & b[293])^(a[14] & b[294])^(a[13] & b[295])^(a[12] & b[296])^(a[11] & b[297])^(a[10] & b[298])^(a[9] & b[299])^(a[8] & b[300])^(a[7] & b[301])^(a[6] & b[302])^(a[5] & b[303])^(a[4] & b[304])^(a[3] & b[305])^(a[2] & b[306])^(a[1] & b[307])^(a[0] & b[308]);
assign y[309] = (a[309] & b[0])^(a[308] & b[1])^(a[307] & b[2])^(a[306] & b[3])^(a[305] & b[4])^(a[304] & b[5])^(a[303] & b[6])^(a[302] & b[7])^(a[301] & b[8])^(a[300] & b[9])^(a[299] & b[10])^(a[298] & b[11])^(a[297] & b[12])^(a[296] & b[13])^(a[295] & b[14])^(a[294] & b[15])^(a[293] & b[16])^(a[292] & b[17])^(a[291] & b[18])^(a[290] & b[19])^(a[289] & b[20])^(a[288] & b[21])^(a[287] & b[22])^(a[286] & b[23])^(a[285] & b[24])^(a[284] & b[25])^(a[283] & b[26])^(a[282] & b[27])^(a[281] & b[28])^(a[280] & b[29])^(a[279] & b[30])^(a[278] & b[31])^(a[277] & b[32])^(a[276] & b[33])^(a[275] & b[34])^(a[274] & b[35])^(a[273] & b[36])^(a[272] & b[37])^(a[271] & b[38])^(a[270] & b[39])^(a[269] & b[40])^(a[268] & b[41])^(a[267] & b[42])^(a[266] & b[43])^(a[265] & b[44])^(a[264] & b[45])^(a[263] & b[46])^(a[262] & b[47])^(a[261] & b[48])^(a[260] & b[49])^(a[259] & b[50])^(a[258] & b[51])^(a[257] & b[52])^(a[256] & b[53])^(a[255] & b[54])^(a[254] & b[55])^(a[253] & b[56])^(a[252] & b[57])^(a[251] & b[58])^(a[250] & b[59])^(a[249] & b[60])^(a[248] & b[61])^(a[247] & b[62])^(a[246] & b[63])^(a[245] & b[64])^(a[244] & b[65])^(a[243] & b[66])^(a[242] & b[67])^(a[241] & b[68])^(a[240] & b[69])^(a[239] & b[70])^(a[238] & b[71])^(a[237] & b[72])^(a[236] & b[73])^(a[235] & b[74])^(a[234] & b[75])^(a[233] & b[76])^(a[232] & b[77])^(a[231] & b[78])^(a[230] & b[79])^(a[229] & b[80])^(a[228] & b[81])^(a[227] & b[82])^(a[226] & b[83])^(a[225] & b[84])^(a[224] & b[85])^(a[223] & b[86])^(a[222] & b[87])^(a[221] & b[88])^(a[220] & b[89])^(a[219] & b[90])^(a[218] & b[91])^(a[217] & b[92])^(a[216] & b[93])^(a[215] & b[94])^(a[214] & b[95])^(a[213] & b[96])^(a[212] & b[97])^(a[211] & b[98])^(a[210] & b[99])^(a[209] & b[100])^(a[208] & b[101])^(a[207] & b[102])^(a[206] & b[103])^(a[205] & b[104])^(a[204] & b[105])^(a[203] & b[106])^(a[202] & b[107])^(a[201] & b[108])^(a[200] & b[109])^(a[199] & b[110])^(a[198] & b[111])^(a[197] & b[112])^(a[196] & b[113])^(a[195] & b[114])^(a[194] & b[115])^(a[193] & b[116])^(a[192] & b[117])^(a[191] & b[118])^(a[190] & b[119])^(a[189] & b[120])^(a[188] & b[121])^(a[187] & b[122])^(a[186] & b[123])^(a[185] & b[124])^(a[184] & b[125])^(a[183] & b[126])^(a[182] & b[127])^(a[181] & b[128])^(a[180] & b[129])^(a[179] & b[130])^(a[178] & b[131])^(a[177] & b[132])^(a[176] & b[133])^(a[175] & b[134])^(a[174] & b[135])^(a[173] & b[136])^(a[172] & b[137])^(a[171] & b[138])^(a[170] & b[139])^(a[169] & b[140])^(a[168] & b[141])^(a[167] & b[142])^(a[166] & b[143])^(a[165] & b[144])^(a[164] & b[145])^(a[163] & b[146])^(a[162] & b[147])^(a[161] & b[148])^(a[160] & b[149])^(a[159] & b[150])^(a[158] & b[151])^(a[157] & b[152])^(a[156] & b[153])^(a[155] & b[154])^(a[154] & b[155])^(a[153] & b[156])^(a[152] & b[157])^(a[151] & b[158])^(a[150] & b[159])^(a[149] & b[160])^(a[148] & b[161])^(a[147] & b[162])^(a[146] & b[163])^(a[145] & b[164])^(a[144] & b[165])^(a[143] & b[166])^(a[142] & b[167])^(a[141] & b[168])^(a[140] & b[169])^(a[139] & b[170])^(a[138] & b[171])^(a[137] & b[172])^(a[136] & b[173])^(a[135] & b[174])^(a[134] & b[175])^(a[133] & b[176])^(a[132] & b[177])^(a[131] & b[178])^(a[130] & b[179])^(a[129] & b[180])^(a[128] & b[181])^(a[127] & b[182])^(a[126] & b[183])^(a[125] & b[184])^(a[124] & b[185])^(a[123] & b[186])^(a[122] & b[187])^(a[121] & b[188])^(a[120] & b[189])^(a[119] & b[190])^(a[118] & b[191])^(a[117] & b[192])^(a[116] & b[193])^(a[115] & b[194])^(a[114] & b[195])^(a[113] & b[196])^(a[112] & b[197])^(a[111] & b[198])^(a[110] & b[199])^(a[109] & b[200])^(a[108] & b[201])^(a[107] & b[202])^(a[106] & b[203])^(a[105] & b[204])^(a[104] & b[205])^(a[103] & b[206])^(a[102] & b[207])^(a[101] & b[208])^(a[100] & b[209])^(a[99] & b[210])^(a[98] & b[211])^(a[97] & b[212])^(a[96] & b[213])^(a[95] & b[214])^(a[94] & b[215])^(a[93] & b[216])^(a[92] & b[217])^(a[91] & b[218])^(a[90] & b[219])^(a[89] & b[220])^(a[88] & b[221])^(a[87] & b[222])^(a[86] & b[223])^(a[85] & b[224])^(a[84] & b[225])^(a[83] & b[226])^(a[82] & b[227])^(a[81] & b[228])^(a[80] & b[229])^(a[79] & b[230])^(a[78] & b[231])^(a[77] & b[232])^(a[76] & b[233])^(a[75] & b[234])^(a[74] & b[235])^(a[73] & b[236])^(a[72] & b[237])^(a[71] & b[238])^(a[70] & b[239])^(a[69] & b[240])^(a[68] & b[241])^(a[67] & b[242])^(a[66] & b[243])^(a[65] & b[244])^(a[64] & b[245])^(a[63] & b[246])^(a[62] & b[247])^(a[61] & b[248])^(a[60] & b[249])^(a[59] & b[250])^(a[58] & b[251])^(a[57] & b[252])^(a[56] & b[253])^(a[55] & b[254])^(a[54] & b[255])^(a[53] & b[256])^(a[52] & b[257])^(a[51] & b[258])^(a[50] & b[259])^(a[49] & b[260])^(a[48] & b[261])^(a[47] & b[262])^(a[46] & b[263])^(a[45] & b[264])^(a[44] & b[265])^(a[43] & b[266])^(a[42] & b[267])^(a[41] & b[268])^(a[40] & b[269])^(a[39] & b[270])^(a[38] & b[271])^(a[37] & b[272])^(a[36] & b[273])^(a[35] & b[274])^(a[34] & b[275])^(a[33] & b[276])^(a[32] & b[277])^(a[31] & b[278])^(a[30] & b[279])^(a[29] & b[280])^(a[28] & b[281])^(a[27] & b[282])^(a[26] & b[283])^(a[25] & b[284])^(a[24] & b[285])^(a[23] & b[286])^(a[22] & b[287])^(a[21] & b[288])^(a[20] & b[289])^(a[19] & b[290])^(a[18] & b[291])^(a[17] & b[292])^(a[16] & b[293])^(a[15] & b[294])^(a[14] & b[295])^(a[13] & b[296])^(a[12] & b[297])^(a[11] & b[298])^(a[10] & b[299])^(a[9] & b[300])^(a[8] & b[301])^(a[7] & b[302])^(a[6] & b[303])^(a[5] & b[304])^(a[4] & b[305])^(a[3] & b[306])^(a[2] & b[307])^(a[1] & b[308])^(a[0] & b[309]);
assign y[310] = (a[310] & b[0])^(a[309] & b[1])^(a[308] & b[2])^(a[307] & b[3])^(a[306] & b[4])^(a[305] & b[5])^(a[304] & b[6])^(a[303] & b[7])^(a[302] & b[8])^(a[301] & b[9])^(a[300] & b[10])^(a[299] & b[11])^(a[298] & b[12])^(a[297] & b[13])^(a[296] & b[14])^(a[295] & b[15])^(a[294] & b[16])^(a[293] & b[17])^(a[292] & b[18])^(a[291] & b[19])^(a[290] & b[20])^(a[289] & b[21])^(a[288] & b[22])^(a[287] & b[23])^(a[286] & b[24])^(a[285] & b[25])^(a[284] & b[26])^(a[283] & b[27])^(a[282] & b[28])^(a[281] & b[29])^(a[280] & b[30])^(a[279] & b[31])^(a[278] & b[32])^(a[277] & b[33])^(a[276] & b[34])^(a[275] & b[35])^(a[274] & b[36])^(a[273] & b[37])^(a[272] & b[38])^(a[271] & b[39])^(a[270] & b[40])^(a[269] & b[41])^(a[268] & b[42])^(a[267] & b[43])^(a[266] & b[44])^(a[265] & b[45])^(a[264] & b[46])^(a[263] & b[47])^(a[262] & b[48])^(a[261] & b[49])^(a[260] & b[50])^(a[259] & b[51])^(a[258] & b[52])^(a[257] & b[53])^(a[256] & b[54])^(a[255] & b[55])^(a[254] & b[56])^(a[253] & b[57])^(a[252] & b[58])^(a[251] & b[59])^(a[250] & b[60])^(a[249] & b[61])^(a[248] & b[62])^(a[247] & b[63])^(a[246] & b[64])^(a[245] & b[65])^(a[244] & b[66])^(a[243] & b[67])^(a[242] & b[68])^(a[241] & b[69])^(a[240] & b[70])^(a[239] & b[71])^(a[238] & b[72])^(a[237] & b[73])^(a[236] & b[74])^(a[235] & b[75])^(a[234] & b[76])^(a[233] & b[77])^(a[232] & b[78])^(a[231] & b[79])^(a[230] & b[80])^(a[229] & b[81])^(a[228] & b[82])^(a[227] & b[83])^(a[226] & b[84])^(a[225] & b[85])^(a[224] & b[86])^(a[223] & b[87])^(a[222] & b[88])^(a[221] & b[89])^(a[220] & b[90])^(a[219] & b[91])^(a[218] & b[92])^(a[217] & b[93])^(a[216] & b[94])^(a[215] & b[95])^(a[214] & b[96])^(a[213] & b[97])^(a[212] & b[98])^(a[211] & b[99])^(a[210] & b[100])^(a[209] & b[101])^(a[208] & b[102])^(a[207] & b[103])^(a[206] & b[104])^(a[205] & b[105])^(a[204] & b[106])^(a[203] & b[107])^(a[202] & b[108])^(a[201] & b[109])^(a[200] & b[110])^(a[199] & b[111])^(a[198] & b[112])^(a[197] & b[113])^(a[196] & b[114])^(a[195] & b[115])^(a[194] & b[116])^(a[193] & b[117])^(a[192] & b[118])^(a[191] & b[119])^(a[190] & b[120])^(a[189] & b[121])^(a[188] & b[122])^(a[187] & b[123])^(a[186] & b[124])^(a[185] & b[125])^(a[184] & b[126])^(a[183] & b[127])^(a[182] & b[128])^(a[181] & b[129])^(a[180] & b[130])^(a[179] & b[131])^(a[178] & b[132])^(a[177] & b[133])^(a[176] & b[134])^(a[175] & b[135])^(a[174] & b[136])^(a[173] & b[137])^(a[172] & b[138])^(a[171] & b[139])^(a[170] & b[140])^(a[169] & b[141])^(a[168] & b[142])^(a[167] & b[143])^(a[166] & b[144])^(a[165] & b[145])^(a[164] & b[146])^(a[163] & b[147])^(a[162] & b[148])^(a[161] & b[149])^(a[160] & b[150])^(a[159] & b[151])^(a[158] & b[152])^(a[157] & b[153])^(a[156] & b[154])^(a[155] & b[155])^(a[154] & b[156])^(a[153] & b[157])^(a[152] & b[158])^(a[151] & b[159])^(a[150] & b[160])^(a[149] & b[161])^(a[148] & b[162])^(a[147] & b[163])^(a[146] & b[164])^(a[145] & b[165])^(a[144] & b[166])^(a[143] & b[167])^(a[142] & b[168])^(a[141] & b[169])^(a[140] & b[170])^(a[139] & b[171])^(a[138] & b[172])^(a[137] & b[173])^(a[136] & b[174])^(a[135] & b[175])^(a[134] & b[176])^(a[133] & b[177])^(a[132] & b[178])^(a[131] & b[179])^(a[130] & b[180])^(a[129] & b[181])^(a[128] & b[182])^(a[127] & b[183])^(a[126] & b[184])^(a[125] & b[185])^(a[124] & b[186])^(a[123] & b[187])^(a[122] & b[188])^(a[121] & b[189])^(a[120] & b[190])^(a[119] & b[191])^(a[118] & b[192])^(a[117] & b[193])^(a[116] & b[194])^(a[115] & b[195])^(a[114] & b[196])^(a[113] & b[197])^(a[112] & b[198])^(a[111] & b[199])^(a[110] & b[200])^(a[109] & b[201])^(a[108] & b[202])^(a[107] & b[203])^(a[106] & b[204])^(a[105] & b[205])^(a[104] & b[206])^(a[103] & b[207])^(a[102] & b[208])^(a[101] & b[209])^(a[100] & b[210])^(a[99] & b[211])^(a[98] & b[212])^(a[97] & b[213])^(a[96] & b[214])^(a[95] & b[215])^(a[94] & b[216])^(a[93] & b[217])^(a[92] & b[218])^(a[91] & b[219])^(a[90] & b[220])^(a[89] & b[221])^(a[88] & b[222])^(a[87] & b[223])^(a[86] & b[224])^(a[85] & b[225])^(a[84] & b[226])^(a[83] & b[227])^(a[82] & b[228])^(a[81] & b[229])^(a[80] & b[230])^(a[79] & b[231])^(a[78] & b[232])^(a[77] & b[233])^(a[76] & b[234])^(a[75] & b[235])^(a[74] & b[236])^(a[73] & b[237])^(a[72] & b[238])^(a[71] & b[239])^(a[70] & b[240])^(a[69] & b[241])^(a[68] & b[242])^(a[67] & b[243])^(a[66] & b[244])^(a[65] & b[245])^(a[64] & b[246])^(a[63] & b[247])^(a[62] & b[248])^(a[61] & b[249])^(a[60] & b[250])^(a[59] & b[251])^(a[58] & b[252])^(a[57] & b[253])^(a[56] & b[254])^(a[55] & b[255])^(a[54] & b[256])^(a[53] & b[257])^(a[52] & b[258])^(a[51] & b[259])^(a[50] & b[260])^(a[49] & b[261])^(a[48] & b[262])^(a[47] & b[263])^(a[46] & b[264])^(a[45] & b[265])^(a[44] & b[266])^(a[43] & b[267])^(a[42] & b[268])^(a[41] & b[269])^(a[40] & b[270])^(a[39] & b[271])^(a[38] & b[272])^(a[37] & b[273])^(a[36] & b[274])^(a[35] & b[275])^(a[34] & b[276])^(a[33] & b[277])^(a[32] & b[278])^(a[31] & b[279])^(a[30] & b[280])^(a[29] & b[281])^(a[28] & b[282])^(a[27] & b[283])^(a[26] & b[284])^(a[25] & b[285])^(a[24] & b[286])^(a[23] & b[287])^(a[22] & b[288])^(a[21] & b[289])^(a[20] & b[290])^(a[19] & b[291])^(a[18] & b[292])^(a[17] & b[293])^(a[16] & b[294])^(a[15] & b[295])^(a[14] & b[296])^(a[13] & b[297])^(a[12] & b[298])^(a[11] & b[299])^(a[10] & b[300])^(a[9] & b[301])^(a[8] & b[302])^(a[7] & b[303])^(a[6] & b[304])^(a[5] & b[305])^(a[4] & b[306])^(a[3] & b[307])^(a[2] & b[308])^(a[1] & b[309])^(a[0] & b[310]);
assign y[311] = (a[311] & b[0])^(a[310] & b[1])^(a[309] & b[2])^(a[308] & b[3])^(a[307] & b[4])^(a[306] & b[5])^(a[305] & b[6])^(a[304] & b[7])^(a[303] & b[8])^(a[302] & b[9])^(a[301] & b[10])^(a[300] & b[11])^(a[299] & b[12])^(a[298] & b[13])^(a[297] & b[14])^(a[296] & b[15])^(a[295] & b[16])^(a[294] & b[17])^(a[293] & b[18])^(a[292] & b[19])^(a[291] & b[20])^(a[290] & b[21])^(a[289] & b[22])^(a[288] & b[23])^(a[287] & b[24])^(a[286] & b[25])^(a[285] & b[26])^(a[284] & b[27])^(a[283] & b[28])^(a[282] & b[29])^(a[281] & b[30])^(a[280] & b[31])^(a[279] & b[32])^(a[278] & b[33])^(a[277] & b[34])^(a[276] & b[35])^(a[275] & b[36])^(a[274] & b[37])^(a[273] & b[38])^(a[272] & b[39])^(a[271] & b[40])^(a[270] & b[41])^(a[269] & b[42])^(a[268] & b[43])^(a[267] & b[44])^(a[266] & b[45])^(a[265] & b[46])^(a[264] & b[47])^(a[263] & b[48])^(a[262] & b[49])^(a[261] & b[50])^(a[260] & b[51])^(a[259] & b[52])^(a[258] & b[53])^(a[257] & b[54])^(a[256] & b[55])^(a[255] & b[56])^(a[254] & b[57])^(a[253] & b[58])^(a[252] & b[59])^(a[251] & b[60])^(a[250] & b[61])^(a[249] & b[62])^(a[248] & b[63])^(a[247] & b[64])^(a[246] & b[65])^(a[245] & b[66])^(a[244] & b[67])^(a[243] & b[68])^(a[242] & b[69])^(a[241] & b[70])^(a[240] & b[71])^(a[239] & b[72])^(a[238] & b[73])^(a[237] & b[74])^(a[236] & b[75])^(a[235] & b[76])^(a[234] & b[77])^(a[233] & b[78])^(a[232] & b[79])^(a[231] & b[80])^(a[230] & b[81])^(a[229] & b[82])^(a[228] & b[83])^(a[227] & b[84])^(a[226] & b[85])^(a[225] & b[86])^(a[224] & b[87])^(a[223] & b[88])^(a[222] & b[89])^(a[221] & b[90])^(a[220] & b[91])^(a[219] & b[92])^(a[218] & b[93])^(a[217] & b[94])^(a[216] & b[95])^(a[215] & b[96])^(a[214] & b[97])^(a[213] & b[98])^(a[212] & b[99])^(a[211] & b[100])^(a[210] & b[101])^(a[209] & b[102])^(a[208] & b[103])^(a[207] & b[104])^(a[206] & b[105])^(a[205] & b[106])^(a[204] & b[107])^(a[203] & b[108])^(a[202] & b[109])^(a[201] & b[110])^(a[200] & b[111])^(a[199] & b[112])^(a[198] & b[113])^(a[197] & b[114])^(a[196] & b[115])^(a[195] & b[116])^(a[194] & b[117])^(a[193] & b[118])^(a[192] & b[119])^(a[191] & b[120])^(a[190] & b[121])^(a[189] & b[122])^(a[188] & b[123])^(a[187] & b[124])^(a[186] & b[125])^(a[185] & b[126])^(a[184] & b[127])^(a[183] & b[128])^(a[182] & b[129])^(a[181] & b[130])^(a[180] & b[131])^(a[179] & b[132])^(a[178] & b[133])^(a[177] & b[134])^(a[176] & b[135])^(a[175] & b[136])^(a[174] & b[137])^(a[173] & b[138])^(a[172] & b[139])^(a[171] & b[140])^(a[170] & b[141])^(a[169] & b[142])^(a[168] & b[143])^(a[167] & b[144])^(a[166] & b[145])^(a[165] & b[146])^(a[164] & b[147])^(a[163] & b[148])^(a[162] & b[149])^(a[161] & b[150])^(a[160] & b[151])^(a[159] & b[152])^(a[158] & b[153])^(a[157] & b[154])^(a[156] & b[155])^(a[155] & b[156])^(a[154] & b[157])^(a[153] & b[158])^(a[152] & b[159])^(a[151] & b[160])^(a[150] & b[161])^(a[149] & b[162])^(a[148] & b[163])^(a[147] & b[164])^(a[146] & b[165])^(a[145] & b[166])^(a[144] & b[167])^(a[143] & b[168])^(a[142] & b[169])^(a[141] & b[170])^(a[140] & b[171])^(a[139] & b[172])^(a[138] & b[173])^(a[137] & b[174])^(a[136] & b[175])^(a[135] & b[176])^(a[134] & b[177])^(a[133] & b[178])^(a[132] & b[179])^(a[131] & b[180])^(a[130] & b[181])^(a[129] & b[182])^(a[128] & b[183])^(a[127] & b[184])^(a[126] & b[185])^(a[125] & b[186])^(a[124] & b[187])^(a[123] & b[188])^(a[122] & b[189])^(a[121] & b[190])^(a[120] & b[191])^(a[119] & b[192])^(a[118] & b[193])^(a[117] & b[194])^(a[116] & b[195])^(a[115] & b[196])^(a[114] & b[197])^(a[113] & b[198])^(a[112] & b[199])^(a[111] & b[200])^(a[110] & b[201])^(a[109] & b[202])^(a[108] & b[203])^(a[107] & b[204])^(a[106] & b[205])^(a[105] & b[206])^(a[104] & b[207])^(a[103] & b[208])^(a[102] & b[209])^(a[101] & b[210])^(a[100] & b[211])^(a[99] & b[212])^(a[98] & b[213])^(a[97] & b[214])^(a[96] & b[215])^(a[95] & b[216])^(a[94] & b[217])^(a[93] & b[218])^(a[92] & b[219])^(a[91] & b[220])^(a[90] & b[221])^(a[89] & b[222])^(a[88] & b[223])^(a[87] & b[224])^(a[86] & b[225])^(a[85] & b[226])^(a[84] & b[227])^(a[83] & b[228])^(a[82] & b[229])^(a[81] & b[230])^(a[80] & b[231])^(a[79] & b[232])^(a[78] & b[233])^(a[77] & b[234])^(a[76] & b[235])^(a[75] & b[236])^(a[74] & b[237])^(a[73] & b[238])^(a[72] & b[239])^(a[71] & b[240])^(a[70] & b[241])^(a[69] & b[242])^(a[68] & b[243])^(a[67] & b[244])^(a[66] & b[245])^(a[65] & b[246])^(a[64] & b[247])^(a[63] & b[248])^(a[62] & b[249])^(a[61] & b[250])^(a[60] & b[251])^(a[59] & b[252])^(a[58] & b[253])^(a[57] & b[254])^(a[56] & b[255])^(a[55] & b[256])^(a[54] & b[257])^(a[53] & b[258])^(a[52] & b[259])^(a[51] & b[260])^(a[50] & b[261])^(a[49] & b[262])^(a[48] & b[263])^(a[47] & b[264])^(a[46] & b[265])^(a[45] & b[266])^(a[44] & b[267])^(a[43] & b[268])^(a[42] & b[269])^(a[41] & b[270])^(a[40] & b[271])^(a[39] & b[272])^(a[38] & b[273])^(a[37] & b[274])^(a[36] & b[275])^(a[35] & b[276])^(a[34] & b[277])^(a[33] & b[278])^(a[32] & b[279])^(a[31] & b[280])^(a[30] & b[281])^(a[29] & b[282])^(a[28] & b[283])^(a[27] & b[284])^(a[26] & b[285])^(a[25] & b[286])^(a[24] & b[287])^(a[23] & b[288])^(a[22] & b[289])^(a[21] & b[290])^(a[20] & b[291])^(a[19] & b[292])^(a[18] & b[293])^(a[17] & b[294])^(a[16] & b[295])^(a[15] & b[296])^(a[14] & b[297])^(a[13] & b[298])^(a[12] & b[299])^(a[11] & b[300])^(a[10] & b[301])^(a[9] & b[302])^(a[8] & b[303])^(a[7] & b[304])^(a[6] & b[305])^(a[5] & b[306])^(a[4] & b[307])^(a[3] & b[308])^(a[2] & b[309])^(a[1] & b[310])^(a[0] & b[311]);
assign y[312] = (a[312] & b[0])^(a[311] & b[1])^(a[310] & b[2])^(a[309] & b[3])^(a[308] & b[4])^(a[307] & b[5])^(a[306] & b[6])^(a[305] & b[7])^(a[304] & b[8])^(a[303] & b[9])^(a[302] & b[10])^(a[301] & b[11])^(a[300] & b[12])^(a[299] & b[13])^(a[298] & b[14])^(a[297] & b[15])^(a[296] & b[16])^(a[295] & b[17])^(a[294] & b[18])^(a[293] & b[19])^(a[292] & b[20])^(a[291] & b[21])^(a[290] & b[22])^(a[289] & b[23])^(a[288] & b[24])^(a[287] & b[25])^(a[286] & b[26])^(a[285] & b[27])^(a[284] & b[28])^(a[283] & b[29])^(a[282] & b[30])^(a[281] & b[31])^(a[280] & b[32])^(a[279] & b[33])^(a[278] & b[34])^(a[277] & b[35])^(a[276] & b[36])^(a[275] & b[37])^(a[274] & b[38])^(a[273] & b[39])^(a[272] & b[40])^(a[271] & b[41])^(a[270] & b[42])^(a[269] & b[43])^(a[268] & b[44])^(a[267] & b[45])^(a[266] & b[46])^(a[265] & b[47])^(a[264] & b[48])^(a[263] & b[49])^(a[262] & b[50])^(a[261] & b[51])^(a[260] & b[52])^(a[259] & b[53])^(a[258] & b[54])^(a[257] & b[55])^(a[256] & b[56])^(a[255] & b[57])^(a[254] & b[58])^(a[253] & b[59])^(a[252] & b[60])^(a[251] & b[61])^(a[250] & b[62])^(a[249] & b[63])^(a[248] & b[64])^(a[247] & b[65])^(a[246] & b[66])^(a[245] & b[67])^(a[244] & b[68])^(a[243] & b[69])^(a[242] & b[70])^(a[241] & b[71])^(a[240] & b[72])^(a[239] & b[73])^(a[238] & b[74])^(a[237] & b[75])^(a[236] & b[76])^(a[235] & b[77])^(a[234] & b[78])^(a[233] & b[79])^(a[232] & b[80])^(a[231] & b[81])^(a[230] & b[82])^(a[229] & b[83])^(a[228] & b[84])^(a[227] & b[85])^(a[226] & b[86])^(a[225] & b[87])^(a[224] & b[88])^(a[223] & b[89])^(a[222] & b[90])^(a[221] & b[91])^(a[220] & b[92])^(a[219] & b[93])^(a[218] & b[94])^(a[217] & b[95])^(a[216] & b[96])^(a[215] & b[97])^(a[214] & b[98])^(a[213] & b[99])^(a[212] & b[100])^(a[211] & b[101])^(a[210] & b[102])^(a[209] & b[103])^(a[208] & b[104])^(a[207] & b[105])^(a[206] & b[106])^(a[205] & b[107])^(a[204] & b[108])^(a[203] & b[109])^(a[202] & b[110])^(a[201] & b[111])^(a[200] & b[112])^(a[199] & b[113])^(a[198] & b[114])^(a[197] & b[115])^(a[196] & b[116])^(a[195] & b[117])^(a[194] & b[118])^(a[193] & b[119])^(a[192] & b[120])^(a[191] & b[121])^(a[190] & b[122])^(a[189] & b[123])^(a[188] & b[124])^(a[187] & b[125])^(a[186] & b[126])^(a[185] & b[127])^(a[184] & b[128])^(a[183] & b[129])^(a[182] & b[130])^(a[181] & b[131])^(a[180] & b[132])^(a[179] & b[133])^(a[178] & b[134])^(a[177] & b[135])^(a[176] & b[136])^(a[175] & b[137])^(a[174] & b[138])^(a[173] & b[139])^(a[172] & b[140])^(a[171] & b[141])^(a[170] & b[142])^(a[169] & b[143])^(a[168] & b[144])^(a[167] & b[145])^(a[166] & b[146])^(a[165] & b[147])^(a[164] & b[148])^(a[163] & b[149])^(a[162] & b[150])^(a[161] & b[151])^(a[160] & b[152])^(a[159] & b[153])^(a[158] & b[154])^(a[157] & b[155])^(a[156] & b[156])^(a[155] & b[157])^(a[154] & b[158])^(a[153] & b[159])^(a[152] & b[160])^(a[151] & b[161])^(a[150] & b[162])^(a[149] & b[163])^(a[148] & b[164])^(a[147] & b[165])^(a[146] & b[166])^(a[145] & b[167])^(a[144] & b[168])^(a[143] & b[169])^(a[142] & b[170])^(a[141] & b[171])^(a[140] & b[172])^(a[139] & b[173])^(a[138] & b[174])^(a[137] & b[175])^(a[136] & b[176])^(a[135] & b[177])^(a[134] & b[178])^(a[133] & b[179])^(a[132] & b[180])^(a[131] & b[181])^(a[130] & b[182])^(a[129] & b[183])^(a[128] & b[184])^(a[127] & b[185])^(a[126] & b[186])^(a[125] & b[187])^(a[124] & b[188])^(a[123] & b[189])^(a[122] & b[190])^(a[121] & b[191])^(a[120] & b[192])^(a[119] & b[193])^(a[118] & b[194])^(a[117] & b[195])^(a[116] & b[196])^(a[115] & b[197])^(a[114] & b[198])^(a[113] & b[199])^(a[112] & b[200])^(a[111] & b[201])^(a[110] & b[202])^(a[109] & b[203])^(a[108] & b[204])^(a[107] & b[205])^(a[106] & b[206])^(a[105] & b[207])^(a[104] & b[208])^(a[103] & b[209])^(a[102] & b[210])^(a[101] & b[211])^(a[100] & b[212])^(a[99] & b[213])^(a[98] & b[214])^(a[97] & b[215])^(a[96] & b[216])^(a[95] & b[217])^(a[94] & b[218])^(a[93] & b[219])^(a[92] & b[220])^(a[91] & b[221])^(a[90] & b[222])^(a[89] & b[223])^(a[88] & b[224])^(a[87] & b[225])^(a[86] & b[226])^(a[85] & b[227])^(a[84] & b[228])^(a[83] & b[229])^(a[82] & b[230])^(a[81] & b[231])^(a[80] & b[232])^(a[79] & b[233])^(a[78] & b[234])^(a[77] & b[235])^(a[76] & b[236])^(a[75] & b[237])^(a[74] & b[238])^(a[73] & b[239])^(a[72] & b[240])^(a[71] & b[241])^(a[70] & b[242])^(a[69] & b[243])^(a[68] & b[244])^(a[67] & b[245])^(a[66] & b[246])^(a[65] & b[247])^(a[64] & b[248])^(a[63] & b[249])^(a[62] & b[250])^(a[61] & b[251])^(a[60] & b[252])^(a[59] & b[253])^(a[58] & b[254])^(a[57] & b[255])^(a[56] & b[256])^(a[55] & b[257])^(a[54] & b[258])^(a[53] & b[259])^(a[52] & b[260])^(a[51] & b[261])^(a[50] & b[262])^(a[49] & b[263])^(a[48] & b[264])^(a[47] & b[265])^(a[46] & b[266])^(a[45] & b[267])^(a[44] & b[268])^(a[43] & b[269])^(a[42] & b[270])^(a[41] & b[271])^(a[40] & b[272])^(a[39] & b[273])^(a[38] & b[274])^(a[37] & b[275])^(a[36] & b[276])^(a[35] & b[277])^(a[34] & b[278])^(a[33] & b[279])^(a[32] & b[280])^(a[31] & b[281])^(a[30] & b[282])^(a[29] & b[283])^(a[28] & b[284])^(a[27] & b[285])^(a[26] & b[286])^(a[25] & b[287])^(a[24] & b[288])^(a[23] & b[289])^(a[22] & b[290])^(a[21] & b[291])^(a[20] & b[292])^(a[19] & b[293])^(a[18] & b[294])^(a[17] & b[295])^(a[16] & b[296])^(a[15] & b[297])^(a[14] & b[298])^(a[13] & b[299])^(a[12] & b[300])^(a[11] & b[301])^(a[10] & b[302])^(a[9] & b[303])^(a[8] & b[304])^(a[7] & b[305])^(a[6] & b[306])^(a[5] & b[307])^(a[4] & b[308])^(a[3] & b[309])^(a[2] & b[310])^(a[1] & b[311])^(a[0] & b[312]);
assign y[313] = (a[313] & b[0])^(a[312] & b[1])^(a[311] & b[2])^(a[310] & b[3])^(a[309] & b[4])^(a[308] & b[5])^(a[307] & b[6])^(a[306] & b[7])^(a[305] & b[8])^(a[304] & b[9])^(a[303] & b[10])^(a[302] & b[11])^(a[301] & b[12])^(a[300] & b[13])^(a[299] & b[14])^(a[298] & b[15])^(a[297] & b[16])^(a[296] & b[17])^(a[295] & b[18])^(a[294] & b[19])^(a[293] & b[20])^(a[292] & b[21])^(a[291] & b[22])^(a[290] & b[23])^(a[289] & b[24])^(a[288] & b[25])^(a[287] & b[26])^(a[286] & b[27])^(a[285] & b[28])^(a[284] & b[29])^(a[283] & b[30])^(a[282] & b[31])^(a[281] & b[32])^(a[280] & b[33])^(a[279] & b[34])^(a[278] & b[35])^(a[277] & b[36])^(a[276] & b[37])^(a[275] & b[38])^(a[274] & b[39])^(a[273] & b[40])^(a[272] & b[41])^(a[271] & b[42])^(a[270] & b[43])^(a[269] & b[44])^(a[268] & b[45])^(a[267] & b[46])^(a[266] & b[47])^(a[265] & b[48])^(a[264] & b[49])^(a[263] & b[50])^(a[262] & b[51])^(a[261] & b[52])^(a[260] & b[53])^(a[259] & b[54])^(a[258] & b[55])^(a[257] & b[56])^(a[256] & b[57])^(a[255] & b[58])^(a[254] & b[59])^(a[253] & b[60])^(a[252] & b[61])^(a[251] & b[62])^(a[250] & b[63])^(a[249] & b[64])^(a[248] & b[65])^(a[247] & b[66])^(a[246] & b[67])^(a[245] & b[68])^(a[244] & b[69])^(a[243] & b[70])^(a[242] & b[71])^(a[241] & b[72])^(a[240] & b[73])^(a[239] & b[74])^(a[238] & b[75])^(a[237] & b[76])^(a[236] & b[77])^(a[235] & b[78])^(a[234] & b[79])^(a[233] & b[80])^(a[232] & b[81])^(a[231] & b[82])^(a[230] & b[83])^(a[229] & b[84])^(a[228] & b[85])^(a[227] & b[86])^(a[226] & b[87])^(a[225] & b[88])^(a[224] & b[89])^(a[223] & b[90])^(a[222] & b[91])^(a[221] & b[92])^(a[220] & b[93])^(a[219] & b[94])^(a[218] & b[95])^(a[217] & b[96])^(a[216] & b[97])^(a[215] & b[98])^(a[214] & b[99])^(a[213] & b[100])^(a[212] & b[101])^(a[211] & b[102])^(a[210] & b[103])^(a[209] & b[104])^(a[208] & b[105])^(a[207] & b[106])^(a[206] & b[107])^(a[205] & b[108])^(a[204] & b[109])^(a[203] & b[110])^(a[202] & b[111])^(a[201] & b[112])^(a[200] & b[113])^(a[199] & b[114])^(a[198] & b[115])^(a[197] & b[116])^(a[196] & b[117])^(a[195] & b[118])^(a[194] & b[119])^(a[193] & b[120])^(a[192] & b[121])^(a[191] & b[122])^(a[190] & b[123])^(a[189] & b[124])^(a[188] & b[125])^(a[187] & b[126])^(a[186] & b[127])^(a[185] & b[128])^(a[184] & b[129])^(a[183] & b[130])^(a[182] & b[131])^(a[181] & b[132])^(a[180] & b[133])^(a[179] & b[134])^(a[178] & b[135])^(a[177] & b[136])^(a[176] & b[137])^(a[175] & b[138])^(a[174] & b[139])^(a[173] & b[140])^(a[172] & b[141])^(a[171] & b[142])^(a[170] & b[143])^(a[169] & b[144])^(a[168] & b[145])^(a[167] & b[146])^(a[166] & b[147])^(a[165] & b[148])^(a[164] & b[149])^(a[163] & b[150])^(a[162] & b[151])^(a[161] & b[152])^(a[160] & b[153])^(a[159] & b[154])^(a[158] & b[155])^(a[157] & b[156])^(a[156] & b[157])^(a[155] & b[158])^(a[154] & b[159])^(a[153] & b[160])^(a[152] & b[161])^(a[151] & b[162])^(a[150] & b[163])^(a[149] & b[164])^(a[148] & b[165])^(a[147] & b[166])^(a[146] & b[167])^(a[145] & b[168])^(a[144] & b[169])^(a[143] & b[170])^(a[142] & b[171])^(a[141] & b[172])^(a[140] & b[173])^(a[139] & b[174])^(a[138] & b[175])^(a[137] & b[176])^(a[136] & b[177])^(a[135] & b[178])^(a[134] & b[179])^(a[133] & b[180])^(a[132] & b[181])^(a[131] & b[182])^(a[130] & b[183])^(a[129] & b[184])^(a[128] & b[185])^(a[127] & b[186])^(a[126] & b[187])^(a[125] & b[188])^(a[124] & b[189])^(a[123] & b[190])^(a[122] & b[191])^(a[121] & b[192])^(a[120] & b[193])^(a[119] & b[194])^(a[118] & b[195])^(a[117] & b[196])^(a[116] & b[197])^(a[115] & b[198])^(a[114] & b[199])^(a[113] & b[200])^(a[112] & b[201])^(a[111] & b[202])^(a[110] & b[203])^(a[109] & b[204])^(a[108] & b[205])^(a[107] & b[206])^(a[106] & b[207])^(a[105] & b[208])^(a[104] & b[209])^(a[103] & b[210])^(a[102] & b[211])^(a[101] & b[212])^(a[100] & b[213])^(a[99] & b[214])^(a[98] & b[215])^(a[97] & b[216])^(a[96] & b[217])^(a[95] & b[218])^(a[94] & b[219])^(a[93] & b[220])^(a[92] & b[221])^(a[91] & b[222])^(a[90] & b[223])^(a[89] & b[224])^(a[88] & b[225])^(a[87] & b[226])^(a[86] & b[227])^(a[85] & b[228])^(a[84] & b[229])^(a[83] & b[230])^(a[82] & b[231])^(a[81] & b[232])^(a[80] & b[233])^(a[79] & b[234])^(a[78] & b[235])^(a[77] & b[236])^(a[76] & b[237])^(a[75] & b[238])^(a[74] & b[239])^(a[73] & b[240])^(a[72] & b[241])^(a[71] & b[242])^(a[70] & b[243])^(a[69] & b[244])^(a[68] & b[245])^(a[67] & b[246])^(a[66] & b[247])^(a[65] & b[248])^(a[64] & b[249])^(a[63] & b[250])^(a[62] & b[251])^(a[61] & b[252])^(a[60] & b[253])^(a[59] & b[254])^(a[58] & b[255])^(a[57] & b[256])^(a[56] & b[257])^(a[55] & b[258])^(a[54] & b[259])^(a[53] & b[260])^(a[52] & b[261])^(a[51] & b[262])^(a[50] & b[263])^(a[49] & b[264])^(a[48] & b[265])^(a[47] & b[266])^(a[46] & b[267])^(a[45] & b[268])^(a[44] & b[269])^(a[43] & b[270])^(a[42] & b[271])^(a[41] & b[272])^(a[40] & b[273])^(a[39] & b[274])^(a[38] & b[275])^(a[37] & b[276])^(a[36] & b[277])^(a[35] & b[278])^(a[34] & b[279])^(a[33] & b[280])^(a[32] & b[281])^(a[31] & b[282])^(a[30] & b[283])^(a[29] & b[284])^(a[28] & b[285])^(a[27] & b[286])^(a[26] & b[287])^(a[25] & b[288])^(a[24] & b[289])^(a[23] & b[290])^(a[22] & b[291])^(a[21] & b[292])^(a[20] & b[293])^(a[19] & b[294])^(a[18] & b[295])^(a[17] & b[296])^(a[16] & b[297])^(a[15] & b[298])^(a[14] & b[299])^(a[13] & b[300])^(a[12] & b[301])^(a[11] & b[302])^(a[10] & b[303])^(a[9] & b[304])^(a[8] & b[305])^(a[7] & b[306])^(a[6] & b[307])^(a[5] & b[308])^(a[4] & b[309])^(a[3] & b[310])^(a[2] & b[311])^(a[1] & b[312])^(a[0] & b[313]);
assign y[314] = (a[314] & b[0])^(a[313] & b[1])^(a[312] & b[2])^(a[311] & b[3])^(a[310] & b[4])^(a[309] & b[5])^(a[308] & b[6])^(a[307] & b[7])^(a[306] & b[8])^(a[305] & b[9])^(a[304] & b[10])^(a[303] & b[11])^(a[302] & b[12])^(a[301] & b[13])^(a[300] & b[14])^(a[299] & b[15])^(a[298] & b[16])^(a[297] & b[17])^(a[296] & b[18])^(a[295] & b[19])^(a[294] & b[20])^(a[293] & b[21])^(a[292] & b[22])^(a[291] & b[23])^(a[290] & b[24])^(a[289] & b[25])^(a[288] & b[26])^(a[287] & b[27])^(a[286] & b[28])^(a[285] & b[29])^(a[284] & b[30])^(a[283] & b[31])^(a[282] & b[32])^(a[281] & b[33])^(a[280] & b[34])^(a[279] & b[35])^(a[278] & b[36])^(a[277] & b[37])^(a[276] & b[38])^(a[275] & b[39])^(a[274] & b[40])^(a[273] & b[41])^(a[272] & b[42])^(a[271] & b[43])^(a[270] & b[44])^(a[269] & b[45])^(a[268] & b[46])^(a[267] & b[47])^(a[266] & b[48])^(a[265] & b[49])^(a[264] & b[50])^(a[263] & b[51])^(a[262] & b[52])^(a[261] & b[53])^(a[260] & b[54])^(a[259] & b[55])^(a[258] & b[56])^(a[257] & b[57])^(a[256] & b[58])^(a[255] & b[59])^(a[254] & b[60])^(a[253] & b[61])^(a[252] & b[62])^(a[251] & b[63])^(a[250] & b[64])^(a[249] & b[65])^(a[248] & b[66])^(a[247] & b[67])^(a[246] & b[68])^(a[245] & b[69])^(a[244] & b[70])^(a[243] & b[71])^(a[242] & b[72])^(a[241] & b[73])^(a[240] & b[74])^(a[239] & b[75])^(a[238] & b[76])^(a[237] & b[77])^(a[236] & b[78])^(a[235] & b[79])^(a[234] & b[80])^(a[233] & b[81])^(a[232] & b[82])^(a[231] & b[83])^(a[230] & b[84])^(a[229] & b[85])^(a[228] & b[86])^(a[227] & b[87])^(a[226] & b[88])^(a[225] & b[89])^(a[224] & b[90])^(a[223] & b[91])^(a[222] & b[92])^(a[221] & b[93])^(a[220] & b[94])^(a[219] & b[95])^(a[218] & b[96])^(a[217] & b[97])^(a[216] & b[98])^(a[215] & b[99])^(a[214] & b[100])^(a[213] & b[101])^(a[212] & b[102])^(a[211] & b[103])^(a[210] & b[104])^(a[209] & b[105])^(a[208] & b[106])^(a[207] & b[107])^(a[206] & b[108])^(a[205] & b[109])^(a[204] & b[110])^(a[203] & b[111])^(a[202] & b[112])^(a[201] & b[113])^(a[200] & b[114])^(a[199] & b[115])^(a[198] & b[116])^(a[197] & b[117])^(a[196] & b[118])^(a[195] & b[119])^(a[194] & b[120])^(a[193] & b[121])^(a[192] & b[122])^(a[191] & b[123])^(a[190] & b[124])^(a[189] & b[125])^(a[188] & b[126])^(a[187] & b[127])^(a[186] & b[128])^(a[185] & b[129])^(a[184] & b[130])^(a[183] & b[131])^(a[182] & b[132])^(a[181] & b[133])^(a[180] & b[134])^(a[179] & b[135])^(a[178] & b[136])^(a[177] & b[137])^(a[176] & b[138])^(a[175] & b[139])^(a[174] & b[140])^(a[173] & b[141])^(a[172] & b[142])^(a[171] & b[143])^(a[170] & b[144])^(a[169] & b[145])^(a[168] & b[146])^(a[167] & b[147])^(a[166] & b[148])^(a[165] & b[149])^(a[164] & b[150])^(a[163] & b[151])^(a[162] & b[152])^(a[161] & b[153])^(a[160] & b[154])^(a[159] & b[155])^(a[158] & b[156])^(a[157] & b[157])^(a[156] & b[158])^(a[155] & b[159])^(a[154] & b[160])^(a[153] & b[161])^(a[152] & b[162])^(a[151] & b[163])^(a[150] & b[164])^(a[149] & b[165])^(a[148] & b[166])^(a[147] & b[167])^(a[146] & b[168])^(a[145] & b[169])^(a[144] & b[170])^(a[143] & b[171])^(a[142] & b[172])^(a[141] & b[173])^(a[140] & b[174])^(a[139] & b[175])^(a[138] & b[176])^(a[137] & b[177])^(a[136] & b[178])^(a[135] & b[179])^(a[134] & b[180])^(a[133] & b[181])^(a[132] & b[182])^(a[131] & b[183])^(a[130] & b[184])^(a[129] & b[185])^(a[128] & b[186])^(a[127] & b[187])^(a[126] & b[188])^(a[125] & b[189])^(a[124] & b[190])^(a[123] & b[191])^(a[122] & b[192])^(a[121] & b[193])^(a[120] & b[194])^(a[119] & b[195])^(a[118] & b[196])^(a[117] & b[197])^(a[116] & b[198])^(a[115] & b[199])^(a[114] & b[200])^(a[113] & b[201])^(a[112] & b[202])^(a[111] & b[203])^(a[110] & b[204])^(a[109] & b[205])^(a[108] & b[206])^(a[107] & b[207])^(a[106] & b[208])^(a[105] & b[209])^(a[104] & b[210])^(a[103] & b[211])^(a[102] & b[212])^(a[101] & b[213])^(a[100] & b[214])^(a[99] & b[215])^(a[98] & b[216])^(a[97] & b[217])^(a[96] & b[218])^(a[95] & b[219])^(a[94] & b[220])^(a[93] & b[221])^(a[92] & b[222])^(a[91] & b[223])^(a[90] & b[224])^(a[89] & b[225])^(a[88] & b[226])^(a[87] & b[227])^(a[86] & b[228])^(a[85] & b[229])^(a[84] & b[230])^(a[83] & b[231])^(a[82] & b[232])^(a[81] & b[233])^(a[80] & b[234])^(a[79] & b[235])^(a[78] & b[236])^(a[77] & b[237])^(a[76] & b[238])^(a[75] & b[239])^(a[74] & b[240])^(a[73] & b[241])^(a[72] & b[242])^(a[71] & b[243])^(a[70] & b[244])^(a[69] & b[245])^(a[68] & b[246])^(a[67] & b[247])^(a[66] & b[248])^(a[65] & b[249])^(a[64] & b[250])^(a[63] & b[251])^(a[62] & b[252])^(a[61] & b[253])^(a[60] & b[254])^(a[59] & b[255])^(a[58] & b[256])^(a[57] & b[257])^(a[56] & b[258])^(a[55] & b[259])^(a[54] & b[260])^(a[53] & b[261])^(a[52] & b[262])^(a[51] & b[263])^(a[50] & b[264])^(a[49] & b[265])^(a[48] & b[266])^(a[47] & b[267])^(a[46] & b[268])^(a[45] & b[269])^(a[44] & b[270])^(a[43] & b[271])^(a[42] & b[272])^(a[41] & b[273])^(a[40] & b[274])^(a[39] & b[275])^(a[38] & b[276])^(a[37] & b[277])^(a[36] & b[278])^(a[35] & b[279])^(a[34] & b[280])^(a[33] & b[281])^(a[32] & b[282])^(a[31] & b[283])^(a[30] & b[284])^(a[29] & b[285])^(a[28] & b[286])^(a[27] & b[287])^(a[26] & b[288])^(a[25] & b[289])^(a[24] & b[290])^(a[23] & b[291])^(a[22] & b[292])^(a[21] & b[293])^(a[20] & b[294])^(a[19] & b[295])^(a[18] & b[296])^(a[17] & b[297])^(a[16] & b[298])^(a[15] & b[299])^(a[14] & b[300])^(a[13] & b[301])^(a[12] & b[302])^(a[11] & b[303])^(a[10] & b[304])^(a[9] & b[305])^(a[8] & b[306])^(a[7] & b[307])^(a[6] & b[308])^(a[5] & b[309])^(a[4] & b[310])^(a[3] & b[311])^(a[2] & b[312])^(a[1] & b[313])^(a[0] & b[314]);
assign y[315] = (a[315] & b[0])^(a[314] & b[1])^(a[313] & b[2])^(a[312] & b[3])^(a[311] & b[4])^(a[310] & b[5])^(a[309] & b[6])^(a[308] & b[7])^(a[307] & b[8])^(a[306] & b[9])^(a[305] & b[10])^(a[304] & b[11])^(a[303] & b[12])^(a[302] & b[13])^(a[301] & b[14])^(a[300] & b[15])^(a[299] & b[16])^(a[298] & b[17])^(a[297] & b[18])^(a[296] & b[19])^(a[295] & b[20])^(a[294] & b[21])^(a[293] & b[22])^(a[292] & b[23])^(a[291] & b[24])^(a[290] & b[25])^(a[289] & b[26])^(a[288] & b[27])^(a[287] & b[28])^(a[286] & b[29])^(a[285] & b[30])^(a[284] & b[31])^(a[283] & b[32])^(a[282] & b[33])^(a[281] & b[34])^(a[280] & b[35])^(a[279] & b[36])^(a[278] & b[37])^(a[277] & b[38])^(a[276] & b[39])^(a[275] & b[40])^(a[274] & b[41])^(a[273] & b[42])^(a[272] & b[43])^(a[271] & b[44])^(a[270] & b[45])^(a[269] & b[46])^(a[268] & b[47])^(a[267] & b[48])^(a[266] & b[49])^(a[265] & b[50])^(a[264] & b[51])^(a[263] & b[52])^(a[262] & b[53])^(a[261] & b[54])^(a[260] & b[55])^(a[259] & b[56])^(a[258] & b[57])^(a[257] & b[58])^(a[256] & b[59])^(a[255] & b[60])^(a[254] & b[61])^(a[253] & b[62])^(a[252] & b[63])^(a[251] & b[64])^(a[250] & b[65])^(a[249] & b[66])^(a[248] & b[67])^(a[247] & b[68])^(a[246] & b[69])^(a[245] & b[70])^(a[244] & b[71])^(a[243] & b[72])^(a[242] & b[73])^(a[241] & b[74])^(a[240] & b[75])^(a[239] & b[76])^(a[238] & b[77])^(a[237] & b[78])^(a[236] & b[79])^(a[235] & b[80])^(a[234] & b[81])^(a[233] & b[82])^(a[232] & b[83])^(a[231] & b[84])^(a[230] & b[85])^(a[229] & b[86])^(a[228] & b[87])^(a[227] & b[88])^(a[226] & b[89])^(a[225] & b[90])^(a[224] & b[91])^(a[223] & b[92])^(a[222] & b[93])^(a[221] & b[94])^(a[220] & b[95])^(a[219] & b[96])^(a[218] & b[97])^(a[217] & b[98])^(a[216] & b[99])^(a[215] & b[100])^(a[214] & b[101])^(a[213] & b[102])^(a[212] & b[103])^(a[211] & b[104])^(a[210] & b[105])^(a[209] & b[106])^(a[208] & b[107])^(a[207] & b[108])^(a[206] & b[109])^(a[205] & b[110])^(a[204] & b[111])^(a[203] & b[112])^(a[202] & b[113])^(a[201] & b[114])^(a[200] & b[115])^(a[199] & b[116])^(a[198] & b[117])^(a[197] & b[118])^(a[196] & b[119])^(a[195] & b[120])^(a[194] & b[121])^(a[193] & b[122])^(a[192] & b[123])^(a[191] & b[124])^(a[190] & b[125])^(a[189] & b[126])^(a[188] & b[127])^(a[187] & b[128])^(a[186] & b[129])^(a[185] & b[130])^(a[184] & b[131])^(a[183] & b[132])^(a[182] & b[133])^(a[181] & b[134])^(a[180] & b[135])^(a[179] & b[136])^(a[178] & b[137])^(a[177] & b[138])^(a[176] & b[139])^(a[175] & b[140])^(a[174] & b[141])^(a[173] & b[142])^(a[172] & b[143])^(a[171] & b[144])^(a[170] & b[145])^(a[169] & b[146])^(a[168] & b[147])^(a[167] & b[148])^(a[166] & b[149])^(a[165] & b[150])^(a[164] & b[151])^(a[163] & b[152])^(a[162] & b[153])^(a[161] & b[154])^(a[160] & b[155])^(a[159] & b[156])^(a[158] & b[157])^(a[157] & b[158])^(a[156] & b[159])^(a[155] & b[160])^(a[154] & b[161])^(a[153] & b[162])^(a[152] & b[163])^(a[151] & b[164])^(a[150] & b[165])^(a[149] & b[166])^(a[148] & b[167])^(a[147] & b[168])^(a[146] & b[169])^(a[145] & b[170])^(a[144] & b[171])^(a[143] & b[172])^(a[142] & b[173])^(a[141] & b[174])^(a[140] & b[175])^(a[139] & b[176])^(a[138] & b[177])^(a[137] & b[178])^(a[136] & b[179])^(a[135] & b[180])^(a[134] & b[181])^(a[133] & b[182])^(a[132] & b[183])^(a[131] & b[184])^(a[130] & b[185])^(a[129] & b[186])^(a[128] & b[187])^(a[127] & b[188])^(a[126] & b[189])^(a[125] & b[190])^(a[124] & b[191])^(a[123] & b[192])^(a[122] & b[193])^(a[121] & b[194])^(a[120] & b[195])^(a[119] & b[196])^(a[118] & b[197])^(a[117] & b[198])^(a[116] & b[199])^(a[115] & b[200])^(a[114] & b[201])^(a[113] & b[202])^(a[112] & b[203])^(a[111] & b[204])^(a[110] & b[205])^(a[109] & b[206])^(a[108] & b[207])^(a[107] & b[208])^(a[106] & b[209])^(a[105] & b[210])^(a[104] & b[211])^(a[103] & b[212])^(a[102] & b[213])^(a[101] & b[214])^(a[100] & b[215])^(a[99] & b[216])^(a[98] & b[217])^(a[97] & b[218])^(a[96] & b[219])^(a[95] & b[220])^(a[94] & b[221])^(a[93] & b[222])^(a[92] & b[223])^(a[91] & b[224])^(a[90] & b[225])^(a[89] & b[226])^(a[88] & b[227])^(a[87] & b[228])^(a[86] & b[229])^(a[85] & b[230])^(a[84] & b[231])^(a[83] & b[232])^(a[82] & b[233])^(a[81] & b[234])^(a[80] & b[235])^(a[79] & b[236])^(a[78] & b[237])^(a[77] & b[238])^(a[76] & b[239])^(a[75] & b[240])^(a[74] & b[241])^(a[73] & b[242])^(a[72] & b[243])^(a[71] & b[244])^(a[70] & b[245])^(a[69] & b[246])^(a[68] & b[247])^(a[67] & b[248])^(a[66] & b[249])^(a[65] & b[250])^(a[64] & b[251])^(a[63] & b[252])^(a[62] & b[253])^(a[61] & b[254])^(a[60] & b[255])^(a[59] & b[256])^(a[58] & b[257])^(a[57] & b[258])^(a[56] & b[259])^(a[55] & b[260])^(a[54] & b[261])^(a[53] & b[262])^(a[52] & b[263])^(a[51] & b[264])^(a[50] & b[265])^(a[49] & b[266])^(a[48] & b[267])^(a[47] & b[268])^(a[46] & b[269])^(a[45] & b[270])^(a[44] & b[271])^(a[43] & b[272])^(a[42] & b[273])^(a[41] & b[274])^(a[40] & b[275])^(a[39] & b[276])^(a[38] & b[277])^(a[37] & b[278])^(a[36] & b[279])^(a[35] & b[280])^(a[34] & b[281])^(a[33] & b[282])^(a[32] & b[283])^(a[31] & b[284])^(a[30] & b[285])^(a[29] & b[286])^(a[28] & b[287])^(a[27] & b[288])^(a[26] & b[289])^(a[25] & b[290])^(a[24] & b[291])^(a[23] & b[292])^(a[22] & b[293])^(a[21] & b[294])^(a[20] & b[295])^(a[19] & b[296])^(a[18] & b[297])^(a[17] & b[298])^(a[16] & b[299])^(a[15] & b[300])^(a[14] & b[301])^(a[13] & b[302])^(a[12] & b[303])^(a[11] & b[304])^(a[10] & b[305])^(a[9] & b[306])^(a[8] & b[307])^(a[7] & b[308])^(a[6] & b[309])^(a[5] & b[310])^(a[4] & b[311])^(a[3] & b[312])^(a[2] & b[313])^(a[1] & b[314])^(a[0] & b[315]);
assign y[316] = (a[316] & b[0])^(a[315] & b[1])^(a[314] & b[2])^(a[313] & b[3])^(a[312] & b[4])^(a[311] & b[5])^(a[310] & b[6])^(a[309] & b[7])^(a[308] & b[8])^(a[307] & b[9])^(a[306] & b[10])^(a[305] & b[11])^(a[304] & b[12])^(a[303] & b[13])^(a[302] & b[14])^(a[301] & b[15])^(a[300] & b[16])^(a[299] & b[17])^(a[298] & b[18])^(a[297] & b[19])^(a[296] & b[20])^(a[295] & b[21])^(a[294] & b[22])^(a[293] & b[23])^(a[292] & b[24])^(a[291] & b[25])^(a[290] & b[26])^(a[289] & b[27])^(a[288] & b[28])^(a[287] & b[29])^(a[286] & b[30])^(a[285] & b[31])^(a[284] & b[32])^(a[283] & b[33])^(a[282] & b[34])^(a[281] & b[35])^(a[280] & b[36])^(a[279] & b[37])^(a[278] & b[38])^(a[277] & b[39])^(a[276] & b[40])^(a[275] & b[41])^(a[274] & b[42])^(a[273] & b[43])^(a[272] & b[44])^(a[271] & b[45])^(a[270] & b[46])^(a[269] & b[47])^(a[268] & b[48])^(a[267] & b[49])^(a[266] & b[50])^(a[265] & b[51])^(a[264] & b[52])^(a[263] & b[53])^(a[262] & b[54])^(a[261] & b[55])^(a[260] & b[56])^(a[259] & b[57])^(a[258] & b[58])^(a[257] & b[59])^(a[256] & b[60])^(a[255] & b[61])^(a[254] & b[62])^(a[253] & b[63])^(a[252] & b[64])^(a[251] & b[65])^(a[250] & b[66])^(a[249] & b[67])^(a[248] & b[68])^(a[247] & b[69])^(a[246] & b[70])^(a[245] & b[71])^(a[244] & b[72])^(a[243] & b[73])^(a[242] & b[74])^(a[241] & b[75])^(a[240] & b[76])^(a[239] & b[77])^(a[238] & b[78])^(a[237] & b[79])^(a[236] & b[80])^(a[235] & b[81])^(a[234] & b[82])^(a[233] & b[83])^(a[232] & b[84])^(a[231] & b[85])^(a[230] & b[86])^(a[229] & b[87])^(a[228] & b[88])^(a[227] & b[89])^(a[226] & b[90])^(a[225] & b[91])^(a[224] & b[92])^(a[223] & b[93])^(a[222] & b[94])^(a[221] & b[95])^(a[220] & b[96])^(a[219] & b[97])^(a[218] & b[98])^(a[217] & b[99])^(a[216] & b[100])^(a[215] & b[101])^(a[214] & b[102])^(a[213] & b[103])^(a[212] & b[104])^(a[211] & b[105])^(a[210] & b[106])^(a[209] & b[107])^(a[208] & b[108])^(a[207] & b[109])^(a[206] & b[110])^(a[205] & b[111])^(a[204] & b[112])^(a[203] & b[113])^(a[202] & b[114])^(a[201] & b[115])^(a[200] & b[116])^(a[199] & b[117])^(a[198] & b[118])^(a[197] & b[119])^(a[196] & b[120])^(a[195] & b[121])^(a[194] & b[122])^(a[193] & b[123])^(a[192] & b[124])^(a[191] & b[125])^(a[190] & b[126])^(a[189] & b[127])^(a[188] & b[128])^(a[187] & b[129])^(a[186] & b[130])^(a[185] & b[131])^(a[184] & b[132])^(a[183] & b[133])^(a[182] & b[134])^(a[181] & b[135])^(a[180] & b[136])^(a[179] & b[137])^(a[178] & b[138])^(a[177] & b[139])^(a[176] & b[140])^(a[175] & b[141])^(a[174] & b[142])^(a[173] & b[143])^(a[172] & b[144])^(a[171] & b[145])^(a[170] & b[146])^(a[169] & b[147])^(a[168] & b[148])^(a[167] & b[149])^(a[166] & b[150])^(a[165] & b[151])^(a[164] & b[152])^(a[163] & b[153])^(a[162] & b[154])^(a[161] & b[155])^(a[160] & b[156])^(a[159] & b[157])^(a[158] & b[158])^(a[157] & b[159])^(a[156] & b[160])^(a[155] & b[161])^(a[154] & b[162])^(a[153] & b[163])^(a[152] & b[164])^(a[151] & b[165])^(a[150] & b[166])^(a[149] & b[167])^(a[148] & b[168])^(a[147] & b[169])^(a[146] & b[170])^(a[145] & b[171])^(a[144] & b[172])^(a[143] & b[173])^(a[142] & b[174])^(a[141] & b[175])^(a[140] & b[176])^(a[139] & b[177])^(a[138] & b[178])^(a[137] & b[179])^(a[136] & b[180])^(a[135] & b[181])^(a[134] & b[182])^(a[133] & b[183])^(a[132] & b[184])^(a[131] & b[185])^(a[130] & b[186])^(a[129] & b[187])^(a[128] & b[188])^(a[127] & b[189])^(a[126] & b[190])^(a[125] & b[191])^(a[124] & b[192])^(a[123] & b[193])^(a[122] & b[194])^(a[121] & b[195])^(a[120] & b[196])^(a[119] & b[197])^(a[118] & b[198])^(a[117] & b[199])^(a[116] & b[200])^(a[115] & b[201])^(a[114] & b[202])^(a[113] & b[203])^(a[112] & b[204])^(a[111] & b[205])^(a[110] & b[206])^(a[109] & b[207])^(a[108] & b[208])^(a[107] & b[209])^(a[106] & b[210])^(a[105] & b[211])^(a[104] & b[212])^(a[103] & b[213])^(a[102] & b[214])^(a[101] & b[215])^(a[100] & b[216])^(a[99] & b[217])^(a[98] & b[218])^(a[97] & b[219])^(a[96] & b[220])^(a[95] & b[221])^(a[94] & b[222])^(a[93] & b[223])^(a[92] & b[224])^(a[91] & b[225])^(a[90] & b[226])^(a[89] & b[227])^(a[88] & b[228])^(a[87] & b[229])^(a[86] & b[230])^(a[85] & b[231])^(a[84] & b[232])^(a[83] & b[233])^(a[82] & b[234])^(a[81] & b[235])^(a[80] & b[236])^(a[79] & b[237])^(a[78] & b[238])^(a[77] & b[239])^(a[76] & b[240])^(a[75] & b[241])^(a[74] & b[242])^(a[73] & b[243])^(a[72] & b[244])^(a[71] & b[245])^(a[70] & b[246])^(a[69] & b[247])^(a[68] & b[248])^(a[67] & b[249])^(a[66] & b[250])^(a[65] & b[251])^(a[64] & b[252])^(a[63] & b[253])^(a[62] & b[254])^(a[61] & b[255])^(a[60] & b[256])^(a[59] & b[257])^(a[58] & b[258])^(a[57] & b[259])^(a[56] & b[260])^(a[55] & b[261])^(a[54] & b[262])^(a[53] & b[263])^(a[52] & b[264])^(a[51] & b[265])^(a[50] & b[266])^(a[49] & b[267])^(a[48] & b[268])^(a[47] & b[269])^(a[46] & b[270])^(a[45] & b[271])^(a[44] & b[272])^(a[43] & b[273])^(a[42] & b[274])^(a[41] & b[275])^(a[40] & b[276])^(a[39] & b[277])^(a[38] & b[278])^(a[37] & b[279])^(a[36] & b[280])^(a[35] & b[281])^(a[34] & b[282])^(a[33] & b[283])^(a[32] & b[284])^(a[31] & b[285])^(a[30] & b[286])^(a[29] & b[287])^(a[28] & b[288])^(a[27] & b[289])^(a[26] & b[290])^(a[25] & b[291])^(a[24] & b[292])^(a[23] & b[293])^(a[22] & b[294])^(a[21] & b[295])^(a[20] & b[296])^(a[19] & b[297])^(a[18] & b[298])^(a[17] & b[299])^(a[16] & b[300])^(a[15] & b[301])^(a[14] & b[302])^(a[13] & b[303])^(a[12] & b[304])^(a[11] & b[305])^(a[10] & b[306])^(a[9] & b[307])^(a[8] & b[308])^(a[7] & b[309])^(a[6] & b[310])^(a[5] & b[311])^(a[4] & b[312])^(a[3] & b[313])^(a[2] & b[314])^(a[1] & b[315])^(a[0] & b[316]);
assign y[317] = (a[317] & b[0])^(a[316] & b[1])^(a[315] & b[2])^(a[314] & b[3])^(a[313] & b[4])^(a[312] & b[5])^(a[311] & b[6])^(a[310] & b[7])^(a[309] & b[8])^(a[308] & b[9])^(a[307] & b[10])^(a[306] & b[11])^(a[305] & b[12])^(a[304] & b[13])^(a[303] & b[14])^(a[302] & b[15])^(a[301] & b[16])^(a[300] & b[17])^(a[299] & b[18])^(a[298] & b[19])^(a[297] & b[20])^(a[296] & b[21])^(a[295] & b[22])^(a[294] & b[23])^(a[293] & b[24])^(a[292] & b[25])^(a[291] & b[26])^(a[290] & b[27])^(a[289] & b[28])^(a[288] & b[29])^(a[287] & b[30])^(a[286] & b[31])^(a[285] & b[32])^(a[284] & b[33])^(a[283] & b[34])^(a[282] & b[35])^(a[281] & b[36])^(a[280] & b[37])^(a[279] & b[38])^(a[278] & b[39])^(a[277] & b[40])^(a[276] & b[41])^(a[275] & b[42])^(a[274] & b[43])^(a[273] & b[44])^(a[272] & b[45])^(a[271] & b[46])^(a[270] & b[47])^(a[269] & b[48])^(a[268] & b[49])^(a[267] & b[50])^(a[266] & b[51])^(a[265] & b[52])^(a[264] & b[53])^(a[263] & b[54])^(a[262] & b[55])^(a[261] & b[56])^(a[260] & b[57])^(a[259] & b[58])^(a[258] & b[59])^(a[257] & b[60])^(a[256] & b[61])^(a[255] & b[62])^(a[254] & b[63])^(a[253] & b[64])^(a[252] & b[65])^(a[251] & b[66])^(a[250] & b[67])^(a[249] & b[68])^(a[248] & b[69])^(a[247] & b[70])^(a[246] & b[71])^(a[245] & b[72])^(a[244] & b[73])^(a[243] & b[74])^(a[242] & b[75])^(a[241] & b[76])^(a[240] & b[77])^(a[239] & b[78])^(a[238] & b[79])^(a[237] & b[80])^(a[236] & b[81])^(a[235] & b[82])^(a[234] & b[83])^(a[233] & b[84])^(a[232] & b[85])^(a[231] & b[86])^(a[230] & b[87])^(a[229] & b[88])^(a[228] & b[89])^(a[227] & b[90])^(a[226] & b[91])^(a[225] & b[92])^(a[224] & b[93])^(a[223] & b[94])^(a[222] & b[95])^(a[221] & b[96])^(a[220] & b[97])^(a[219] & b[98])^(a[218] & b[99])^(a[217] & b[100])^(a[216] & b[101])^(a[215] & b[102])^(a[214] & b[103])^(a[213] & b[104])^(a[212] & b[105])^(a[211] & b[106])^(a[210] & b[107])^(a[209] & b[108])^(a[208] & b[109])^(a[207] & b[110])^(a[206] & b[111])^(a[205] & b[112])^(a[204] & b[113])^(a[203] & b[114])^(a[202] & b[115])^(a[201] & b[116])^(a[200] & b[117])^(a[199] & b[118])^(a[198] & b[119])^(a[197] & b[120])^(a[196] & b[121])^(a[195] & b[122])^(a[194] & b[123])^(a[193] & b[124])^(a[192] & b[125])^(a[191] & b[126])^(a[190] & b[127])^(a[189] & b[128])^(a[188] & b[129])^(a[187] & b[130])^(a[186] & b[131])^(a[185] & b[132])^(a[184] & b[133])^(a[183] & b[134])^(a[182] & b[135])^(a[181] & b[136])^(a[180] & b[137])^(a[179] & b[138])^(a[178] & b[139])^(a[177] & b[140])^(a[176] & b[141])^(a[175] & b[142])^(a[174] & b[143])^(a[173] & b[144])^(a[172] & b[145])^(a[171] & b[146])^(a[170] & b[147])^(a[169] & b[148])^(a[168] & b[149])^(a[167] & b[150])^(a[166] & b[151])^(a[165] & b[152])^(a[164] & b[153])^(a[163] & b[154])^(a[162] & b[155])^(a[161] & b[156])^(a[160] & b[157])^(a[159] & b[158])^(a[158] & b[159])^(a[157] & b[160])^(a[156] & b[161])^(a[155] & b[162])^(a[154] & b[163])^(a[153] & b[164])^(a[152] & b[165])^(a[151] & b[166])^(a[150] & b[167])^(a[149] & b[168])^(a[148] & b[169])^(a[147] & b[170])^(a[146] & b[171])^(a[145] & b[172])^(a[144] & b[173])^(a[143] & b[174])^(a[142] & b[175])^(a[141] & b[176])^(a[140] & b[177])^(a[139] & b[178])^(a[138] & b[179])^(a[137] & b[180])^(a[136] & b[181])^(a[135] & b[182])^(a[134] & b[183])^(a[133] & b[184])^(a[132] & b[185])^(a[131] & b[186])^(a[130] & b[187])^(a[129] & b[188])^(a[128] & b[189])^(a[127] & b[190])^(a[126] & b[191])^(a[125] & b[192])^(a[124] & b[193])^(a[123] & b[194])^(a[122] & b[195])^(a[121] & b[196])^(a[120] & b[197])^(a[119] & b[198])^(a[118] & b[199])^(a[117] & b[200])^(a[116] & b[201])^(a[115] & b[202])^(a[114] & b[203])^(a[113] & b[204])^(a[112] & b[205])^(a[111] & b[206])^(a[110] & b[207])^(a[109] & b[208])^(a[108] & b[209])^(a[107] & b[210])^(a[106] & b[211])^(a[105] & b[212])^(a[104] & b[213])^(a[103] & b[214])^(a[102] & b[215])^(a[101] & b[216])^(a[100] & b[217])^(a[99] & b[218])^(a[98] & b[219])^(a[97] & b[220])^(a[96] & b[221])^(a[95] & b[222])^(a[94] & b[223])^(a[93] & b[224])^(a[92] & b[225])^(a[91] & b[226])^(a[90] & b[227])^(a[89] & b[228])^(a[88] & b[229])^(a[87] & b[230])^(a[86] & b[231])^(a[85] & b[232])^(a[84] & b[233])^(a[83] & b[234])^(a[82] & b[235])^(a[81] & b[236])^(a[80] & b[237])^(a[79] & b[238])^(a[78] & b[239])^(a[77] & b[240])^(a[76] & b[241])^(a[75] & b[242])^(a[74] & b[243])^(a[73] & b[244])^(a[72] & b[245])^(a[71] & b[246])^(a[70] & b[247])^(a[69] & b[248])^(a[68] & b[249])^(a[67] & b[250])^(a[66] & b[251])^(a[65] & b[252])^(a[64] & b[253])^(a[63] & b[254])^(a[62] & b[255])^(a[61] & b[256])^(a[60] & b[257])^(a[59] & b[258])^(a[58] & b[259])^(a[57] & b[260])^(a[56] & b[261])^(a[55] & b[262])^(a[54] & b[263])^(a[53] & b[264])^(a[52] & b[265])^(a[51] & b[266])^(a[50] & b[267])^(a[49] & b[268])^(a[48] & b[269])^(a[47] & b[270])^(a[46] & b[271])^(a[45] & b[272])^(a[44] & b[273])^(a[43] & b[274])^(a[42] & b[275])^(a[41] & b[276])^(a[40] & b[277])^(a[39] & b[278])^(a[38] & b[279])^(a[37] & b[280])^(a[36] & b[281])^(a[35] & b[282])^(a[34] & b[283])^(a[33] & b[284])^(a[32] & b[285])^(a[31] & b[286])^(a[30] & b[287])^(a[29] & b[288])^(a[28] & b[289])^(a[27] & b[290])^(a[26] & b[291])^(a[25] & b[292])^(a[24] & b[293])^(a[23] & b[294])^(a[22] & b[295])^(a[21] & b[296])^(a[20] & b[297])^(a[19] & b[298])^(a[18] & b[299])^(a[17] & b[300])^(a[16] & b[301])^(a[15] & b[302])^(a[14] & b[303])^(a[13] & b[304])^(a[12] & b[305])^(a[11] & b[306])^(a[10] & b[307])^(a[9] & b[308])^(a[8] & b[309])^(a[7] & b[310])^(a[6] & b[311])^(a[5] & b[312])^(a[4] & b[313])^(a[3] & b[314])^(a[2] & b[315])^(a[1] & b[316])^(a[0] & b[317]);
assign y[318] = (a[318] & b[0])^(a[317] & b[1])^(a[316] & b[2])^(a[315] & b[3])^(a[314] & b[4])^(a[313] & b[5])^(a[312] & b[6])^(a[311] & b[7])^(a[310] & b[8])^(a[309] & b[9])^(a[308] & b[10])^(a[307] & b[11])^(a[306] & b[12])^(a[305] & b[13])^(a[304] & b[14])^(a[303] & b[15])^(a[302] & b[16])^(a[301] & b[17])^(a[300] & b[18])^(a[299] & b[19])^(a[298] & b[20])^(a[297] & b[21])^(a[296] & b[22])^(a[295] & b[23])^(a[294] & b[24])^(a[293] & b[25])^(a[292] & b[26])^(a[291] & b[27])^(a[290] & b[28])^(a[289] & b[29])^(a[288] & b[30])^(a[287] & b[31])^(a[286] & b[32])^(a[285] & b[33])^(a[284] & b[34])^(a[283] & b[35])^(a[282] & b[36])^(a[281] & b[37])^(a[280] & b[38])^(a[279] & b[39])^(a[278] & b[40])^(a[277] & b[41])^(a[276] & b[42])^(a[275] & b[43])^(a[274] & b[44])^(a[273] & b[45])^(a[272] & b[46])^(a[271] & b[47])^(a[270] & b[48])^(a[269] & b[49])^(a[268] & b[50])^(a[267] & b[51])^(a[266] & b[52])^(a[265] & b[53])^(a[264] & b[54])^(a[263] & b[55])^(a[262] & b[56])^(a[261] & b[57])^(a[260] & b[58])^(a[259] & b[59])^(a[258] & b[60])^(a[257] & b[61])^(a[256] & b[62])^(a[255] & b[63])^(a[254] & b[64])^(a[253] & b[65])^(a[252] & b[66])^(a[251] & b[67])^(a[250] & b[68])^(a[249] & b[69])^(a[248] & b[70])^(a[247] & b[71])^(a[246] & b[72])^(a[245] & b[73])^(a[244] & b[74])^(a[243] & b[75])^(a[242] & b[76])^(a[241] & b[77])^(a[240] & b[78])^(a[239] & b[79])^(a[238] & b[80])^(a[237] & b[81])^(a[236] & b[82])^(a[235] & b[83])^(a[234] & b[84])^(a[233] & b[85])^(a[232] & b[86])^(a[231] & b[87])^(a[230] & b[88])^(a[229] & b[89])^(a[228] & b[90])^(a[227] & b[91])^(a[226] & b[92])^(a[225] & b[93])^(a[224] & b[94])^(a[223] & b[95])^(a[222] & b[96])^(a[221] & b[97])^(a[220] & b[98])^(a[219] & b[99])^(a[218] & b[100])^(a[217] & b[101])^(a[216] & b[102])^(a[215] & b[103])^(a[214] & b[104])^(a[213] & b[105])^(a[212] & b[106])^(a[211] & b[107])^(a[210] & b[108])^(a[209] & b[109])^(a[208] & b[110])^(a[207] & b[111])^(a[206] & b[112])^(a[205] & b[113])^(a[204] & b[114])^(a[203] & b[115])^(a[202] & b[116])^(a[201] & b[117])^(a[200] & b[118])^(a[199] & b[119])^(a[198] & b[120])^(a[197] & b[121])^(a[196] & b[122])^(a[195] & b[123])^(a[194] & b[124])^(a[193] & b[125])^(a[192] & b[126])^(a[191] & b[127])^(a[190] & b[128])^(a[189] & b[129])^(a[188] & b[130])^(a[187] & b[131])^(a[186] & b[132])^(a[185] & b[133])^(a[184] & b[134])^(a[183] & b[135])^(a[182] & b[136])^(a[181] & b[137])^(a[180] & b[138])^(a[179] & b[139])^(a[178] & b[140])^(a[177] & b[141])^(a[176] & b[142])^(a[175] & b[143])^(a[174] & b[144])^(a[173] & b[145])^(a[172] & b[146])^(a[171] & b[147])^(a[170] & b[148])^(a[169] & b[149])^(a[168] & b[150])^(a[167] & b[151])^(a[166] & b[152])^(a[165] & b[153])^(a[164] & b[154])^(a[163] & b[155])^(a[162] & b[156])^(a[161] & b[157])^(a[160] & b[158])^(a[159] & b[159])^(a[158] & b[160])^(a[157] & b[161])^(a[156] & b[162])^(a[155] & b[163])^(a[154] & b[164])^(a[153] & b[165])^(a[152] & b[166])^(a[151] & b[167])^(a[150] & b[168])^(a[149] & b[169])^(a[148] & b[170])^(a[147] & b[171])^(a[146] & b[172])^(a[145] & b[173])^(a[144] & b[174])^(a[143] & b[175])^(a[142] & b[176])^(a[141] & b[177])^(a[140] & b[178])^(a[139] & b[179])^(a[138] & b[180])^(a[137] & b[181])^(a[136] & b[182])^(a[135] & b[183])^(a[134] & b[184])^(a[133] & b[185])^(a[132] & b[186])^(a[131] & b[187])^(a[130] & b[188])^(a[129] & b[189])^(a[128] & b[190])^(a[127] & b[191])^(a[126] & b[192])^(a[125] & b[193])^(a[124] & b[194])^(a[123] & b[195])^(a[122] & b[196])^(a[121] & b[197])^(a[120] & b[198])^(a[119] & b[199])^(a[118] & b[200])^(a[117] & b[201])^(a[116] & b[202])^(a[115] & b[203])^(a[114] & b[204])^(a[113] & b[205])^(a[112] & b[206])^(a[111] & b[207])^(a[110] & b[208])^(a[109] & b[209])^(a[108] & b[210])^(a[107] & b[211])^(a[106] & b[212])^(a[105] & b[213])^(a[104] & b[214])^(a[103] & b[215])^(a[102] & b[216])^(a[101] & b[217])^(a[100] & b[218])^(a[99] & b[219])^(a[98] & b[220])^(a[97] & b[221])^(a[96] & b[222])^(a[95] & b[223])^(a[94] & b[224])^(a[93] & b[225])^(a[92] & b[226])^(a[91] & b[227])^(a[90] & b[228])^(a[89] & b[229])^(a[88] & b[230])^(a[87] & b[231])^(a[86] & b[232])^(a[85] & b[233])^(a[84] & b[234])^(a[83] & b[235])^(a[82] & b[236])^(a[81] & b[237])^(a[80] & b[238])^(a[79] & b[239])^(a[78] & b[240])^(a[77] & b[241])^(a[76] & b[242])^(a[75] & b[243])^(a[74] & b[244])^(a[73] & b[245])^(a[72] & b[246])^(a[71] & b[247])^(a[70] & b[248])^(a[69] & b[249])^(a[68] & b[250])^(a[67] & b[251])^(a[66] & b[252])^(a[65] & b[253])^(a[64] & b[254])^(a[63] & b[255])^(a[62] & b[256])^(a[61] & b[257])^(a[60] & b[258])^(a[59] & b[259])^(a[58] & b[260])^(a[57] & b[261])^(a[56] & b[262])^(a[55] & b[263])^(a[54] & b[264])^(a[53] & b[265])^(a[52] & b[266])^(a[51] & b[267])^(a[50] & b[268])^(a[49] & b[269])^(a[48] & b[270])^(a[47] & b[271])^(a[46] & b[272])^(a[45] & b[273])^(a[44] & b[274])^(a[43] & b[275])^(a[42] & b[276])^(a[41] & b[277])^(a[40] & b[278])^(a[39] & b[279])^(a[38] & b[280])^(a[37] & b[281])^(a[36] & b[282])^(a[35] & b[283])^(a[34] & b[284])^(a[33] & b[285])^(a[32] & b[286])^(a[31] & b[287])^(a[30] & b[288])^(a[29] & b[289])^(a[28] & b[290])^(a[27] & b[291])^(a[26] & b[292])^(a[25] & b[293])^(a[24] & b[294])^(a[23] & b[295])^(a[22] & b[296])^(a[21] & b[297])^(a[20] & b[298])^(a[19] & b[299])^(a[18] & b[300])^(a[17] & b[301])^(a[16] & b[302])^(a[15] & b[303])^(a[14] & b[304])^(a[13] & b[305])^(a[12] & b[306])^(a[11] & b[307])^(a[10] & b[308])^(a[9] & b[309])^(a[8] & b[310])^(a[7] & b[311])^(a[6] & b[312])^(a[5] & b[313])^(a[4] & b[314])^(a[3] & b[315])^(a[2] & b[316])^(a[1] & b[317])^(a[0] & b[318]);
assign y[319] = (a[319] & b[0])^(a[318] & b[1])^(a[317] & b[2])^(a[316] & b[3])^(a[315] & b[4])^(a[314] & b[5])^(a[313] & b[6])^(a[312] & b[7])^(a[311] & b[8])^(a[310] & b[9])^(a[309] & b[10])^(a[308] & b[11])^(a[307] & b[12])^(a[306] & b[13])^(a[305] & b[14])^(a[304] & b[15])^(a[303] & b[16])^(a[302] & b[17])^(a[301] & b[18])^(a[300] & b[19])^(a[299] & b[20])^(a[298] & b[21])^(a[297] & b[22])^(a[296] & b[23])^(a[295] & b[24])^(a[294] & b[25])^(a[293] & b[26])^(a[292] & b[27])^(a[291] & b[28])^(a[290] & b[29])^(a[289] & b[30])^(a[288] & b[31])^(a[287] & b[32])^(a[286] & b[33])^(a[285] & b[34])^(a[284] & b[35])^(a[283] & b[36])^(a[282] & b[37])^(a[281] & b[38])^(a[280] & b[39])^(a[279] & b[40])^(a[278] & b[41])^(a[277] & b[42])^(a[276] & b[43])^(a[275] & b[44])^(a[274] & b[45])^(a[273] & b[46])^(a[272] & b[47])^(a[271] & b[48])^(a[270] & b[49])^(a[269] & b[50])^(a[268] & b[51])^(a[267] & b[52])^(a[266] & b[53])^(a[265] & b[54])^(a[264] & b[55])^(a[263] & b[56])^(a[262] & b[57])^(a[261] & b[58])^(a[260] & b[59])^(a[259] & b[60])^(a[258] & b[61])^(a[257] & b[62])^(a[256] & b[63])^(a[255] & b[64])^(a[254] & b[65])^(a[253] & b[66])^(a[252] & b[67])^(a[251] & b[68])^(a[250] & b[69])^(a[249] & b[70])^(a[248] & b[71])^(a[247] & b[72])^(a[246] & b[73])^(a[245] & b[74])^(a[244] & b[75])^(a[243] & b[76])^(a[242] & b[77])^(a[241] & b[78])^(a[240] & b[79])^(a[239] & b[80])^(a[238] & b[81])^(a[237] & b[82])^(a[236] & b[83])^(a[235] & b[84])^(a[234] & b[85])^(a[233] & b[86])^(a[232] & b[87])^(a[231] & b[88])^(a[230] & b[89])^(a[229] & b[90])^(a[228] & b[91])^(a[227] & b[92])^(a[226] & b[93])^(a[225] & b[94])^(a[224] & b[95])^(a[223] & b[96])^(a[222] & b[97])^(a[221] & b[98])^(a[220] & b[99])^(a[219] & b[100])^(a[218] & b[101])^(a[217] & b[102])^(a[216] & b[103])^(a[215] & b[104])^(a[214] & b[105])^(a[213] & b[106])^(a[212] & b[107])^(a[211] & b[108])^(a[210] & b[109])^(a[209] & b[110])^(a[208] & b[111])^(a[207] & b[112])^(a[206] & b[113])^(a[205] & b[114])^(a[204] & b[115])^(a[203] & b[116])^(a[202] & b[117])^(a[201] & b[118])^(a[200] & b[119])^(a[199] & b[120])^(a[198] & b[121])^(a[197] & b[122])^(a[196] & b[123])^(a[195] & b[124])^(a[194] & b[125])^(a[193] & b[126])^(a[192] & b[127])^(a[191] & b[128])^(a[190] & b[129])^(a[189] & b[130])^(a[188] & b[131])^(a[187] & b[132])^(a[186] & b[133])^(a[185] & b[134])^(a[184] & b[135])^(a[183] & b[136])^(a[182] & b[137])^(a[181] & b[138])^(a[180] & b[139])^(a[179] & b[140])^(a[178] & b[141])^(a[177] & b[142])^(a[176] & b[143])^(a[175] & b[144])^(a[174] & b[145])^(a[173] & b[146])^(a[172] & b[147])^(a[171] & b[148])^(a[170] & b[149])^(a[169] & b[150])^(a[168] & b[151])^(a[167] & b[152])^(a[166] & b[153])^(a[165] & b[154])^(a[164] & b[155])^(a[163] & b[156])^(a[162] & b[157])^(a[161] & b[158])^(a[160] & b[159])^(a[159] & b[160])^(a[158] & b[161])^(a[157] & b[162])^(a[156] & b[163])^(a[155] & b[164])^(a[154] & b[165])^(a[153] & b[166])^(a[152] & b[167])^(a[151] & b[168])^(a[150] & b[169])^(a[149] & b[170])^(a[148] & b[171])^(a[147] & b[172])^(a[146] & b[173])^(a[145] & b[174])^(a[144] & b[175])^(a[143] & b[176])^(a[142] & b[177])^(a[141] & b[178])^(a[140] & b[179])^(a[139] & b[180])^(a[138] & b[181])^(a[137] & b[182])^(a[136] & b[183])^(a[135] & b[184])^(a[134] & b[185])^(a[133] & b[186])^(a[132] & b[187])^(a[131] & b[188])^(a[130] & b[189])^(a[129] & b[190])^(a[128] & b[191])^(a[127] & b[192])^(a[126] & b[193])^(a[125] & b[194])^(a[124] & b[195])^(a[123] & b[196])^(a[122] & b[197])^(a[121] & b[198])^(a[120] & b[199])^(a[119] & b[200])^(a[118] & b[201])^(a[117] & b[202])^(a[116] & b[203])^(a[115] & b[204])^(a[114] & b[205])^(a[113] & b[206])^(a[112] & b[207])^(a[111] & b[208])^(a[110] & b[209])^(a[109] & b[210])^(a[108] & b[211])^(a[107] & b[212])^(a[106] & b[213])^(a[105] & b[214])^(a[104] & b[215])^(a[103] & b[216])^(a[102] & b[217])^(a[101] & b[218])^(a[100] & b[219])^(a[99] & b[220])^(a[98] & b[221])^(a[97] & b[222])^(a[96] & b[223])^(a[95] & b[224])^(a[94] & b[225])^(a[93] & b[226])^(a[92] & b[227])^(a[91] & b[228])^(a[90] & b[229])^(a[89] & b[230])^(a[88] & b[231])^(a[87] & b[232])^(a[86] & b[233])^(a[85] & b[234])^(a[84] & b[235])^(a[83] & b[236])^(a[82] & b[237])^(a[81] & b[238])^(a[80] & b[239])^(a[79] & b[240])^(a[78] & b[241])^(a[77] & b[242])^(a[76] & b[243])^(a[75] & b[244])^(a[74] & b[245])^(a[73] & b[246])^(a[72] & b[247])^(a[71] & b[248])^(a[70] & b[249])^(a[69] & b[250])^(a[68] & b[251])^(a[67] & b[252])^(a[66] & b[253])^(a[65] & b[254])^(a[64] & b[255])^(a[63] & b[256])^(a[62] & b[257])^(a[61] & b[258])^(a[60] & b[259])^(a[59] & b[260])^(a[58] & b[261])^(a[57] & b[262])^(a[56] & b[263])^(a[55] & b[264])^(a[54] & b[265])^(a[53] & b[266])^(a[52] & b[267])^(a[51] & b[268])^(a[50] & b[269])^(a[49] & b[270])^(a[48] & b[271])^(a[47] & b[272])^(a[46] & b[273])^(a[45] & b[274])^(a[44] & b[275])^(a[43] & b[276])^(a[42] & b[277])^(a[41] & b[278])^(a[40] & b[279])^(a[39] & b[280])^(a[38] & b[281])^(a[37] & b[282])^(a[36] & b[283])^(a[35] & b[284])^(a[34] & b[285])^(a[33] & b[286])^(a[32] & b[287])^(a[31] & b[288])^(a[30] & b[289])^(a[29] & b[290])^(a[28] & b[291])^(a[27] & b[292])^(a[26] & b[293])^(a[25] & b[294])^(a[24] & b[295])^(a[23] & b[296])^(a[22] & b[297])^(a[21] & b[298])^(a[20] & b[299])^(a[19] & b[300])^(a[18] & b[301])^(a[17] & b[302])^(a[16] & b[303])^(a[15] & b[304])^(a[14] & b[305])^(a[13] & b[306])^(a[12] & b[307])^(a[11] & b[308])^(a[10] & b[309])^(a[9] & b[310])^(a[8] & b[311])^(a[7] & b[312])^(a[6] & b[313])^(a[5] & b[314])^(a[4] & b[315])^(a[3] & b[316])^(a[2] & b[317])^(a[1] & b[318])^(a[0] & b[319]);
assign y[320] = (a[320] & b[0])^(a[319] & b[1])^(a[318] & b[2])^(a[317] & b[3])^(a[316] & b[4])^(a[315] & b[5])^(a[314] & b[6])^(a[313] & b[7])^(a[312] & b[8])^(a[311] & b[9])^(a[310] & b[10])^(a[309] & b[11])^(a[308] & b[12])^(a[307] & b[13])^(a[306] & b[14])^(a[305] & b[15])^(a[304] & b[16])^(a[303] & b[17])^(a[302] & b[18])^(a[301] & b[19])^(a[300] & b[20])^(a[299] & b[21])^(a[298] & b[22])^(a[297] & b[23])^(a[296] & b[24])^(a[295] & b[25])^(a[294] & b[26])^(a[293] & b[27])^(a[292] & b[28])^(a[291] & b[29])^(a[290] & b[30])^(a[289] & b[31])^(a[288] & b[32])^(a[287] & b[33])^(a[286] & b[34])^(a[285] & b[35])^(a[284] & b[36])^(a[283] & b[37])^(a[282] & b[38])^(a[281] & b[39])^(a[280] & b[40])^(a[279] & b[41])^(a[278] & b[42])^(a[277] & b[43])^(a[276] & b[44])^(a[275] & b[45])^(a[274] & b[46])^(a[273] & b[47])^(a[272] & b[48])^(a[271] & b[49])^(a[270] & b[50])^(a[269] & b[51])^(a[268] & b[52])^(a[267] & b[53])^(a[266] & b[54])^(a[265] & b[55])^(a[264] & b[56])^(a[263] & b[57])^(a[262] & b[58])^(a[261] & b[59])^(a[260] & b[60])^(a[259] & b[61])^(a[258] & b[62])^(a[257] & b[63])^(a[256] & b[64])^(a[255] & b[65])^(a[254] & b[66])^(a[253] & b[67])^(a[252] & b[68])^(a[251] & b[69])^(a[250] & b[70])^(a[249] & b[71])^(a[248] & b[72])^(a[247] & b[73])^(a[246] & b[74])^(a[245] & b[75])^(a[244] & b[76])^(a[243] & b[77])^(a[242] & b[78])^(a[241] & b[79])^(a[240] & b[80])^(a[239] & b[81])^(a[238] & b[82])^(a[237] & b[83])^(a[236] & b[84])^(a[235] & b[85])^(a[234] & b[86])^(a[233] & b[87])^(a[232] & b[88])^(a[231] & b[89])^(a[230] & b[90])^(a[229] & b[91])^(a[228] & b[92])^(a[227] & b[93])^(a[226] & b[94])^(a[225] & b[95])^(a[224] & b[96])^(a[223] & b[97])^(a[222] & b[98])^(a[221] & b[99])^(a[220] & b[100])^(a[219] & b[101])^(a[218] & b[102])^(a[217] & b[103])^(a[216] & b[104])^(a[215] & b[105])^(a[214] & b[106])^(a[213] & b[107])^(a[212] & b[108])^(a[211] & b[109])^(a[210] & b[110])^(a[209] & b[111])^(a[208] & b[112])^(a[207] & b[113])^(a[206] & b[114])^(a[205] & b[115])^(a[204] & b[116])^(a[203] & b[117])^(a[202] & b[118])^(a[201] & b[119])^(a[200] & b[120])^(a[199] & b[121])^(a[198] & b[122])^(a[197] & b[123])^(a[196] & b[124])^(a[195] & b[125])^(a[194] & b[126])^(a[193] & b[127])^(a[192] & b[128])^(a[191] & b[129])^(a[190] & b[130])^(a[189] & b[131])^(a[188] & b[132])^(a[187] & b[133])^(a[186] & b[134])^(a[185] & b[135])^(a[184] & b[136])^(a[183] & b[137])^(a[182] & b[138])^(a[181] & b[139])^(a[180] & b[140])^(a[179] & b[141])^(a[178] & b[142])^(a[177] & b[143])^(a[176] & b[144])^(a[175] & b[145])^(a[174] & b[146])^(a[173] & b[147])^(a[172] & b[148])^(a[171] & b[149])^(a[170] & b[150])^(a[169] & b[151])^(a[168] & b[152])^(a[167] & b[153])^(a[166] & b[154])^(a[165] & b[155])^(a[164] & b[156])^(a[163] & b[157])^(a[162] & b[158])^(a[161] & b[159])^(a[160] & b[160])^(a[159] & b[161])^(a[158] & b[162])^(a[157] & b[163])^(a[156] & b[164])^(a[155] & b[165])^(a[154] & b[166])^(a[153] & b[167])^(a[152] & b[168])^(a[151] & b[169])^(a[150] & b[170])^(a[149] & b[171])^(a[148] & b[172])^(a[147] & b[173])^(a[146] & b[174])^(a[145] & b[175])^(a[144] & b[176])^(a[143] & b[177])^(a[142] & b[178])^(a[141] & b[179])^(a[140] & b[180])^(a[139] & b[181])^(a[138] & b[182])^(a[137] & b[183])^(a[136] & b[184])^(a[135] & b[185])^(a[134] & b[186])^(a[133] & b[187])^(a[132] & b[188])^(a[131] & b[189])^(a[130] & b[190])^(a[129] & b[191])^(a[128] & b[192])^(a[127] & b[193])^(a[126] & b[194])^(a[125] & b[195])^(a[124] & b[196])^(a[123] & b[197])^(a[122] & b[198])^(a[121] & b[199])^(a[120] & b[200])^(a[119] & b[201])^(a[118] & b[202])^(a[117] & b[203])^(a[116] & b[204])^(a[115] & b[205])^(a[114] & b[206])^(a[113] & b[207])^(a[112] & b[208])^(a[111] & b[209])^(a[110] & b[210])^(a[109] & b[211])^(a[108] & b[212])^(a[107] & b[213])^(a[106] & b[214])^(a[105] & b[215])^(a[104] & b[216])^(a[103] & b[217])^(a[102] & b[218])^(a[101] & b[219])^(a[100] & b[220])^(a[99] & b[221])^(a[98] & b[222])^(a[97] & b[223])^(a[96] & b[224])^(a[95] & b[225])^(a[94] & b[226])^(a[93] & b[227])^(a[92] & b[228])^(a[91] & b[229])^(a[90] & b[230])^(a[89] & b[231])^(a[88] & b[232])^(a[87] & b[233])^(a[86] & b[234])^(a[85] & b[235])^(a[84] & b[236])^(a[83] & b[237])^(a[82] & b[238])^(a[81] & b[239])^(a[80] & b[240])^(a[79] & b[241])^(a[78] & b[242])^(a[77] & b[243])^(a[76] & b[244])^(a[75] & b[245])^(a[74] & b[246])^(a[73] & b[247])^(a[72] & b[248])^(a[71] & b[249])^(a[70] & b[250])^(a[69] & b[251])^(a[68] & b[252])^(a[67] & b[253])^(a[66] & b[254])^(a[65] & b[255])^(a[64] & b[256])^(a[63] & b[257])^(a[62] & b[258])^(a[61] & b[259])^(a[60] & b[260])^(a[59] & b[261])^(a[58] & b[262])^(a[57] & b[263])^(a[56] & b[264])^(a[55] & b[265])^(a[54] & b[266])^(a[53] & b[267])^(a[52] & b[268])^(a[51] & b[269])^(a[50] & b[270])^(a[49] & b[271])^(a[48] & b[272])^(a[47] & b[273])^(a[46] & b[274])^(a[45] & b[275])^(a[44] & b[276])^(a[43] & b[277])^(a[42] & b[278])^(a[41] & b[279])^(a[40] & b[280])^(a[39] & b[281])^(a[38] & b[282])^(a[37] & b[283])^(a[36] & b[284])^(a[35] & b[285])^(a[34] & b[286])^(a[33] & b[287])^(a[32] & b[288])^(a[31] & b[289])^(a[30] & b[290])^(a[29] & b[291])^(a[28] & b[292])^(a[27] & b[293])^(a[26] & b[294])^(a[25] & b[295])^(a[24] & b[296])^(a[23] & b[297])^(a[22] & b[298])^(a[21] & b[299])^(a[20] & b[300])^(a[19] & b[301])^(a[18] & b[302])^(a[17] & b[303])^(a[16] & b[304])^(a[15] & b[305])^(a[14] & b[306])^(a[13] & b[307])^(a[12] & b[308])^(a[11] & b[309])^(a[10] & b[310])^(a[9] & b[311])^(a[8] & b[312])^(a[7] & b[313])^(a[6] & b[314])^(a[5] & b[315])^(a[4] & b[316])^(a[3] & b[317])^(a[2] & b[318])^(a[1] & b[319])^(a[0] & b[320]);
assign y[321] = (a[321] & b[0])^(a[320] & b[1])^(a[319] & b[2])^(a[318] & b[3])^(a[317] & b[4])^(a[316] & b[5])^(a[315] & b[6])^(a[314] & b[7])^(a[313] & b[8])^(a[312] & b[9])^(a[311] & b[10])^(a[310] & b[11])^(a[309] & b[12])^(a[308] & b[13])^(a[307] & b[14])^(a[306] & b[15])^(a[305] & b[16])^(a[304] & b[17])^(a[303] & b[18])^(a[302] & b[19])^(a[301] & b[20])^(a[300] & b[21])^(a[299] & b[22])^(a[298] & b[23])^(a[297] & b[24])^(a[296] & b[25])^(a[295] & b[26])^(a[294] & b[27])^(a[293] & b[28])^(a[292] & b[29])^(a[291] & b[30])^(a[290] & b[31])^(a[289] & b[32])^(a[288] & b[33])^(a[287] & b[34])^(a[286] & b[35])^(a[285] & b[36])^(a[284] & b[37])^(a[283] & b[38])^(a[282] & b[39])^(a[281] & b[40])^(a[280] & b[41])^(a[279] & b[42])^(a[278] & b[43])^(a[277] & b[44])^(a[276] & b[45])^(a[275] & b[46])^(a[274] & b[47])^(a[273] & b[48])^(a[272] & b[49])^(a[271] & b[50])^(a[270] & b[51])^(a[269] & b[52])^(a[268] & b[53])^(a[267] & b[54])^(a[266] & b[55])^(a[265] & b[56])^(a[264] & b[57])^(a[263] & b[58])^(a[262] & b[59])^(a[261] & b[60])^(a[260] & b[61])^(a[259] & b[62])^(a[258] & b[63])^(a[257] & b[64])^(a[256] & b[65])^(a[255] & b[66])^(a[254] & b[67])^(a[253] & b[68])^(a[252] & b[69])^(a[251] & b[70])^(a[250] & b[71])^(a[249] & b[72])^(a[248] & b[73])^(a[247] & b[74])^(a[246] & b[75])^(a[245] & b[76])^(a[244] & b[77])^(a[243] & b[78])^(a[242] & b[79])^(a[241] & b[80])^(a[240] & b[81])^(a[239] & b[82])^(a[238] & b[83])^(a[237] & b[84])^(a[236] & b[85])^(a[235] & b[86])^(a[234] & b[87])^(a[233] & b[88])^(a[232] & b[89])^(a[231] & b[90])^(a[230] & b[91])^(a[229] & b[92])^(a[228] & b[93])^(a[227] & b[94])^(a[226] & b[95])^(a[225] & b[96])^(a[224] & b[97])^(a[223] & b[98])^(a[222] & b[99])^(a[221] & b[100])^(a[220] & b[101])^(a[219] & b[102])^(a[218] & b[103])^(a[217] & b[104])^(a[216] & b[105])^(a[215] & b[106])^(a[214] & b[107])^(a[213] & b[108])^(a[212] & b[109])^(a[211] & b[110])^(a[210] & b[111])^(a[209] & b[112])^(a[208] & b[113])^(a[207] & b[114])^(a[206] & b[115])^(a[205] & b[116])^(a[204] & b[117])^(a[203] & b[118])^(a[202] & b[119])^(a[201] & b[120])^(a[200] & b[121])^(a[199] & b[122])^(a[198] & b[123])^(a[197] & b[124])^(a[196] & b[125])^(a[195] & b[126])^(a[194] & b[127])^(a[193] & b[128])^(a[192] & b[129])^(a[191] & b[130])^(a[190] & b[131])^(a[189] & b[132])^(a[188] & b[133])^(a[187] & b[134])^(a[186] & b[135])^(a[185] & b[136])^(a[184] & b[137])^(a[183] & b[138])^(a[182] & b[139])^(a[181] & b[140])^(a[180] & b[141])^(a[179] & b[142])^(a[178] & b[143])^(a[177] & b[144])^(a[176] & b[145])^(a[175] & b[146])^(a[174] & b[147])^(a[173] & b[148])^(a[172] & b[149])^(a[171] & b[150])^(a[170] & b[151])^(a[169] & b[152])^(a[168] & b[153])^(a[167] & b[154])^(a[166] & b[155])^(a[165] & b[156])^(a[164] & b[157])^(a[163] & b[158])^(a[162] & b[159])^(a[161] & b[160])^(a[160] & b[161])^(a[159] & b[162])^(a[158] & b[163])^(a[157] & b[164])^(a[156] & b[165])^(a[155] & b[166])^(a[154] & b[167])^(a[153] & b[168])^(a[152] & b[169])^(a[151] & b[170])^(a[150] & b[171])^(a[149] & b[172])^(a[148] & b[173])^(a[147] & b[174])^(a[146] & b[175])^(a[145] & b[176])^(a[144] & b[177])^(a[143] & b[178])^(a[142] & b[179])^(a[141] & b[180])^(a[140] & b[181])^(a[139] & b[182])^(a[138] & b[183])^(a[137] & b[184])^(a[136] & b[185])^(a[135] & b[186])^(a[134] & b[187])^(a[133] & b[188])^(a[132] & b[189])^(a[131] & b[190])^(a[130] & b[191])^(a[129] & b[192])^(a[128] & b[193])^(a[127] & b[194])^(a[126] & b[195])^(a[125] & b[196])^(a[124] & b[197])^(a[123] & b[198])^(a[122] & b[199])^(a[121] & b[200])^(a[120] & b[201])^(a[119] & b[202])^(a[118] & b[203])^(a[117] & b[204])^(a[116] & b[205])^(a[115] & b[206])^(a[114] & b[207])^(a[113] & b[208])^(a[112] & b[209])^(a[111] & b[210])^(a[110] & b[211])^(a[109] & b[212])^(a[108] & b[213])^(a[107] & b[214])^(a[106] & b[215])^(a[105] & b[216])^(a[104] & b[217])^(a[103] & b[218])^(a[102] & b[219])^(a[101] & b[220])^(a[100] & b[221])^(a[99] & b[222])^(a[98] & b[223])^(a[97] & b[224])^(a[96] & b[225])^(a[95] & b[226])^(a[94] & b[227])^(a[93] & b[228])^(a[92] & b[229])^(a[91] & b[230])^(a[90] & b[231])^(a[89] & b[232])^(a[88] & b[233])^(a[87] & b[234])^(a[86] & b[235])^(a[85] & b[236])^(a[84] & b[237])^(a[83] & b[238])^(a[82] & b[239])^(a[81] & b[240])^(a[80] & b[241])^(a[79] & b[242])^(a[78] & b[243])^(a[77] & b[244])^(a[76] & b[245])^(a[75] & b[246])^(a[74] & b[247])^(a[73] & b[248])^(a[72] & b[249])^(a[71] & b[250])^(a[70] & b[251])^(a[69] & b[252])^(a[68] & b[253])^(a[67] & b[254])^(a[66] & b[255])^(a[65] & b[256])^(a[64] & b[257])^(a[63] & b[258])^(a[62] & b[259])^(a[61] & b[260])^(a[60] & b[261])^(a[59] & b[262])^(a[58] & b[263])^(a[57] & b[264])^(a[56] & b[265])^(a[55] & b[266])^(a[54] & b[267])^(a[53] & b[268])^(a[52] & b[269])^(a[51] & b[270])^(a[50] & b[271])^(a[49] & b[272])^(a[48] & b[273])^(a[47] & b[274])^(a[46] & b[275])^(a[45] & b[276])^(a[44] & b[277])^(a[43] & b[278])^(a[42] & b[279])^(a[41] & b[280])^(a[40] & b[281])^(a[39] & b[282])^(a[38] & b[283])^(a[37] & b[284])^(a[36] & b[285])^(a[35] & b[286])^(a[34] & b[287])^(a[33] & b[288])^(a[32] & b[289])^(a[31] & b[290])^(a[30] & b[291])^(a[29] & b[292])^(a[28] & b[293])^(a[27] & b[294])^(a[26] & b[295])^(a[25] & b[296])^(a[24] & b[297])^(a[23] & b[298])^(a[22] & b[299])^(a[21] & b[300])^(a[20] & b[301])^(a[19] & b[302])^(a[18] & b[303])^(a[17] & b[304])^(a[16] & b[305])^(a[15] & b[306])^(a[14] & b[307])^(a[13] & b[308])^(a[12] & b[309])^(a[11] & b[310])^(a[10] & b[311])^(a[9] & b[312])^(a[8] & b[313])^(a[7] & b[314])^(a[6] & b[315])^(a[5] & b[316])^(a[4] & b[317])^(a[3] & b[318])^(a[2] & b[319])^(a[1] & b[320])^(a[0] & b[321]);
assign y[322] = (a[322] & b[0])^(a[321] & b[1])^(a[320] & b[2])^(a[319] & b[3])^(a[318] & b[4])^(a[317] & b[5])^(a[316] & b[6])^(a[315] & b[7])^(a[314] & b[8])^(a[313] & b[9])^(a[312] & b[10])^(a[311] & b[11])^(a[310] & b[12])^(a[309] & b[13])^(a[308] & b[14])^(a[307] & b[15])^(a[306] & b[16])^(a[305] & b[17])^(a[304] & b[18])^(a[303] & b[19])^(a[302] & b[20])^(a[301] & b[21])^(a[300] & b[22])^(a[299] & b[23])^(a[298] & b[24])^(a[297] & b[25])^(a[296] & b[26])^(a[295] & b[27])^(a[294] & b[28])^(a[293] & b[29])^(a[292] & b[30])^(a[291] & b[31])^(a[290] & b[32])^(a[289] & b[33])^(a[288] & b[34])^(a[287] & b[35])^(a[286] & b[36])^(a[285] & b[37])^(a[284] & b[38])^(a[283] & b[39])^(a[282] & b[40])^(a[281] & b[41])^(a[280] & b[42])^(a[279] & b[43])^(a[278] & b[44])^(a[277] & b[45])^(a[276] & b[46])^(a[275] & b[47])^(a[274] & b[48])^(a[273] & b[49])^(a[272] & b[50])^(a[271] & b[51])^(a[270] & b[52])^(a[269] & b[53])^(a[268] & b[54])^(a[267] & b[55])^(a[266] & b[56])^(a[265] & b[57])^(a[264] & b[58])^(a[263] & b[59])^(a[262] & b[60])^(a[261] & b[61])^(a[260] & b[62])^(a[259] & b[63])^(a[258] & b[64])^(a[257] & b[65])^(a[256] & b[66])^(a[255] & b[67])^(a[254] & b[68])^(a[253] & b[69])^(a[252] & b[70])^(a[251] & b[71])^(a[250] & b[72])^(a[249] & b[73])^(a[248] & b[74])^(a[247] & b[75])^(a[246] & b[76])^(a[245] & b[77])^(a[244] & b[78])^(a[243] & b[79])^(a[242] & b[80])^(a[241] & b[81])^(a[240] & b[82])^(a[239] & b[83])^(a[238] & b[84])^(a[237] & b[85])^(a[236] & b[86])^(a[235] & b[87])^(a[234] & b[88])^(a[233] & b[89])^(a[232] & b[90])^(a[231] & b[91])^(a[230] & b[92])^(a[229] & b[93])^(a[228] & b[94])^(a[227] & b[95])^(a[226] & b[96])^(a[225] & b[97])^(a[224] & b[98])^(a[223] & b[99])^(a[222] & b[100])^(a[221] & b[101])^(a[220] & b[102])^(a[219] & b[103])^(a[218] & b[104])^(a[217] & b[105])^(a[216] & b[106])^(a[215] & b[107])^(a[214] & b[108])^(a[213] & b[109])^(a[212] & b[110])^(a[211] & b[111])^(a[210] & b[112])^(a[209] & b[113])^(a[208] & b[114])^(a[207] & b[115])^(a[206] & b[116])^(a[205] & b[117])^(a[204] & b[118])^(a[203] & b[119])^(a[202] & b[120])^(a[201] & b[121])^(a[200] & b[122])^(a[199] & b[123])^(a[198] & b[124])^(a[197] & b[125])^(a[196] & b[126])^(a[195] & b[127])^(a[194] & b[128])^(a[193] & b[129])^(a[192] & b[130])^(a[191] & b[131])^(a[190] & b[132])^(a[189] & b[133])^(a[188] & b[134])^(a[187] & b[135])^(a[186] & b[136])^(a[185] & b[137])^(a[184] & b[138])^(a[183] & b[139])^(a[182] & b[140])^(a[181] & b[141])^(a[180] & b[142])^(a[179] & b[143])^(a[178] & b[144])^(a[177] & b[145])^(a[176] & b[146])^(a[175] & b[147])^(a[174] & b[148])^(a[173] & b[149])^(a[172] & b[150])^(a[171] & b[151])^(a[170] & b[152])^(a[169] & b[153])^(a[168] & b[154])^(a[167] & b[155])^(a[166] & b[156])^(a[165] & b[157])^(a[164] & b[158])^(a[163] & b[159])^(a[162] & b[160])^(a[161] & b[161])^(a[160] & b[162])^(a[159] & b[163])^(a[158] & b[164])^(a[157] & b[165])^(a[156] & b[166])^(a[155] & b[167])^(a[154] & b[168])^(a[153] & b[169])^(a[152] & b[170])^(a[151] & b[171])^(a[150] & b[172])^(a[149] & b[173])^(a[148] & b[174])^(a[147] & b[175])^(a[146] & b[176])^(a[145] & b[177])^(a[144] & b[178])^(a[143] & b[179])^(a[142] & b[180])^(a[141] & b[181])^(a[140] & b[182])^(a[139] & b[183])^(a[138] & b[184])^(a[137] & b[185])^(a[136] & b[186])^(a[135] & b[187])^(a[134] & b[188])^(a[133] & b[189])^(a[132] & b[190])^(a[131] & b[191])^(a[130] & b[192])^(a[129] & b[193])^(a[128] & b[194])^(a[127] & b[195])^(a[126] & b[196])^(a[125] & b[197])^(a[124] & b[198])^(a[123] & b[199])^(a[122] & b[200])^(a[121] & b[201])^(a[120] & b[202])^(a[119] & b[203])^(a[118] & b[204])^(a[117] & b[205])^(a[116] & b[206])^(a[115] & b[207])^(a[114] & b[208])^(a[113] & b[209])^(a[112] & b[210])^(a[111] & b[211])^(a[110] & b[212])^(a[109] & b[213])^(a[108] & b[214])^(a[107] & b[215])^(a[106] & b[216])^(a[105] & b[217])^(a[104] & b[218])^(a[103] & b[219])^(a[102] & b[220])^(a[101] & b[221])^(a[100] & b[222])^(a[99] & b[223])^(a[98] & b[224])^(a[97] & b[225])^(a[96] & b[226])^(a[95] & b[227])^(a[94] & b[228])^(a[93] & b[229])^(a[92] & b[230])^(a[91] & b[231])^(a[90] & b[232])^(a[89] & b[233])^(a[88] & b[234])^(a[87] & b[235])^(a[86] & b[236])^(a[85] & b[237])^(a[84] & b[238])^(a[83] & b[239])^(a[82] & b[240])^(a[81] & b[241])^(a[80] & b[242])^(a[79] & b[243])^(a[78] & b[244])^(a[77] & b[245])^(a[76] & b[246])^(a[75] & b[247])^(a[74] & b[248])^(a[73] & b[249])^(a[72] & b[250])^(a[71] & b[251])^(a[70] & b[252])^(a[69] & b[253])^(a[68] & b[254])^(a[67] & b[255])^(a[66] & b[256])^(a[65] & b[257])^(a[64] & b[258])^(a[63] & b[259])^(a[62] & b[260])^(a[61] & b[261])^(a[60] & b[262])^(a[59] & b[263])^(a[58] & b[264])^(a[57] & b[265])^(a[56] & b[266])^(a[55] & b[267])^(a[54] & b[268])^(a[53] & b[269])^(a[52] & b[270])^(a[51] & b[271])^(a[50] & b[272])^(a[49] & b[273])^(a[48] & b[274])^(a[47] & b[275])^(a[46] & b[276])^(a[45] & b[277])^(a[44] & b[278])^(a[43] & b[279])^(a[42] & b[280])^(a[41] & b[281])^(a[40] & b[282])^(a[39] & b[283])^(a[38] & b[284])^(a[37] & b[285])^(a[36] & b[286])^(a[35] & b[287])^(a[34] & b[288])^(a[33] & b[289])^(a[32] & b[290])^(a[31] & b[291])^(a[30] & b[292])^(a[29] & b[293])^(a[28] & b[294])^(a[27] & b[295])^(a[26] & b[296])^(a[25] & b[297])^(a[24] & b[298])^(a[23] & b[299])^(a[22] & b[300])^(a[21] & b[301])^(a[20] & b[302])^(a[19] & b[303])^(a[18] & b[304])^(a[17] & b[305])^(a[16] & b[306])^(a[15] & b[307])^(a[14] & b[308])^(a[13] & b[309])^(a[12] & b[310])^(a[11] & b[311])^(a[10] & b[312])^(a[9] & b[313])^(a[8] & b[314])^(a[7] & b[315])^(a[6] & b[316])^(a[5] & b[317])^(a[4] & b[318])^(a[3] & b[319])^(a[2] & b[320])^(a[1] & b[321])^(a[0] & b[322]);
assign y[323] = (a[323] & b[0])^(a[322] & b[1])^(a[321] & b[2])^(a[320] & b[3])^(a[319] & b[4])^(a[318] & b[5])^(a[317] & b[6])^(a[316] & b[7])^(a[315] & b[8])^(a[314] & b[9])^(a[313] & b[10])^(a[312] & b[11])^(a[311] & b[12])^(a[310] & b[13])^(a[309] & b[14])^(a[308] & b[15])^(a[307] & b[16])^(a[306] & b[17])^(a[305] & b[18])^(a[304] & b[19])^(a[303] & b[20])^(a[302] & b[21])^(a[301] & b[22])^(a[300] & b[23])^(a[299] & b[24])^(a[298] & b[25])^(a[297] & b[26])^(a[296] & b[27])^(a[295] & b[28])^(a[294] & b[29])^(a[293] & b[30])^(a[292] & b[31])^(a[291] & b[32])^(a[290] & b[33])^(a[289] & b[34])^(a[288] & b[35])^(a[287] & b[36])^(a[286] & b[37])^(a[285] & b[38])^(a[284] & b[39])^(a[283] & b[40])^(a[282] & b[41])^(a[281] & b[42])^(a[280] & b[43])^(a[279] & b[44])^(a[278] & b[45])^(a[277] & b[46])^(a[276] & b[47])^(a[275] & b[48])^(a[274] & b[49])^(a[273] & b[50])^(a[272] & b[51])^(a[271] & b[52])^(a[270] & b[53])^(a[269] & b[54])^(a[268] & b[55])^(a[267] & b[56])^(a[266] & b[57])^(a[265] & b[58])^(a[264] & b[59])^(a[263] & b[60])^(a[262] & b[61])^(a[261] & b[62])^(a[260] & b[63])^(a[259] & b[64])^(a[258] & b[65])^(a[257] & b[66])^(a[256] & b[67])^(a[255] & b[68])^(a[254] & b[69])^(a[253] & b[70])^(a[252] & b[71])^(a[251] & b[72])^(a[250] & b[73])^(a[249] & b[74])^(a[248] & b[75])^(a[247] & b[76])^(a[246] & b[77])^(a[245] & b[78])^(a[244] & b[79])^(a[243] & b[80])^(a[242] & b[81])^(a[241] & b[82])^(a[240] & b[83])^(a[239] & b[84])^(a[238] & b[85])^(a[237] & b[86])^(a[236] & b[87])^(a[235] & b[88])^(a[234] & b[89])^(a[233] & b[90])^(a[232] & b[91])^(a[231] & b[92])^(a[230] & b[93])^(a[229] & b[94])^(a[228] & b[95])^(a[227] & b[96])^(a[226] & b[97])^(a[225] & b[98])^(a[224] & b[99])^(a[223] & b[100])^(a[222] & b[101])^(a[221] & b[102])^(a[220] & b[103])^(a[219] & b[104])^(a[218] & b[105])^(a[217] & b[106])^(a[216] & b[107])^(a[215] & b[108])^(a[214] & b[109])^(a[213] & b[110])^(a[212] & b[111])^(a[211] & b[112])^(a[210] & b[113])^(a[209] & b[114])^(a[208] & b[115])^(a[207] & b[116])^(a[206] & b[117])^(a[205] & b[118])^(a[204] & b[119])^(a[203] & b[120])^(a[202] & b[121])^(a[201] & b[122])^(a[200] & b[123])^(a[199] & b[124])^(a[198] & b[125])^(a[197] & b[126])^(a[196] & b[127])^(a[195] & b[128])^(a[194] & b[129])^(a[193] & b[130])^(a[192] & b[131])^(a[191] & b[132])^(a[190] & b[133])^(a[189] & b[134])^(a[188] & b[135])^(a[187] & b[136])^(a[186] & b[137])^(a[185] & b[138])^(a[184] & b[139])^(a[183] & b[140])^(a[182] & b[141])^(a[181] & b[142])^(a[180] & b[143])^(a[179] & b[144])^(a[178] & b[145])^(a[177] & b[146])^(a[176] & b[147])^(a[175] & b[148])^(a[174] & b[149])^(a[173] & b[150])^(a[172] & b[151])^(a[171] & b[152])^(a[170] & b[153])^(a[169] & b[154])^(a[168] & b[155])^(a[167] & b[156])^(a[166] & b[157])^(a[165] & b[158])^(a[164] & b[159])^(a[163] & b[160])^(a[162] & b[161])^(a[161] & b[162])^(a[160] & b[163])^(a[159] & b[164])^(a[158] & b[165])^(a[157] & b[166])^(a[156] & b[167])^(a[155] & b[168])^(a[154] & b[169])^(a[153] & b[170])^(a[152] & b[171])^(a[151] & b[172])^(a[150] & b[173])^(a[149] & b[174])^(a[148] & b[175])^(a[147] & b[176])^(a[146] & b[177])^(a[145] & b[178])^(a[144] & b[179])^(a[143] & b[180])^(a[142] & b[181])^(a[141] & b[182])^(a[140] & b[183])^(a[139] & b[184])^(a[138] & b[185])^(a[137] & b[186])^(a[136] & b[187])^(a[135] & b[188])^(a[134] & b[189])^(a[133] & b[190])^(a[132] & b[191])^(a[131] & b[192])^(a[130] & b[193])^(a[129] & b[194])^(a[128] & b[195])^(a[127] & b[196])^(a[126] & b[197])^(a[125] & b[198])^(a[124] & b[199])^(a[123] & b[200])^(a[122] & b[201])^(a[121] & b[202])^(a[120] & b[203])^(a[119] & b[204])^(a[118] & b[205])^(a[117] & b[206])^(a[116] & b[207])^(a[115] & b[208])^(a[114] & b[209])^(a[113] & b[210])^(a[112] & b[211])^(a[111] & b[212])^(a[110] & b[213])^(a[109] & b[214])^(a[108] & b[215])^(a[107] & b[216])^(a[106] & b[217])^(a[105] & b[218])^(a[104] & b[219])^(a[103] & b[220])^(a[102] & b[221])^(a[101] & b[222])^(a[100] & b[223])^(a[99] & b[224])^(a[98] & b[225])^(a[97] & b[226])^(a[96] & b[227])^(a[95] & b[228])^(a[94] & b[229])^(a[93] & b[230])^(a[92] & b[231])^(a[91] & b[232])^(a[90] & b[233])^(a[89] & b[234])^(a[88] & b[235])^(a[87] & b[236])^(a[86] & b[237])^(a[85] & b[238])^(a[84] & b[239])^(a[83] & b[240])^(a[82] & b[241])^(a[81] & b[242])^(a[80] & b[243])^(a[79] & b[244])^(a[78] & b[245])^(a[77] & b[246])^(a[76] & b[247])^(a[75] & b[248])^(a[74] & b[249])^(a[73] & b[250])^(a[72] & b[251])^(a[71] & b[252])^(a[70] & b[253])^(a[69] & b[254])^(a[68] & b[255])^(a[67] & b[256])^(a[66] & b[257])^(a[65] & b[258])^(a[64] & b[259])^(a[63] & b[260])^(a[62] & b[261])^(a[61] & b[262])^(a[60] & b[263])^(a[59] & b[264])^(a[58] & b[265])^(a[57] & b[266])^(a[56] & b[267])^(a[55] & b[268])^(a[54] & b[269])^(a[53] & b[270])^(a[52] & b[271])^(a[51] & b[272])^(a[50] & b[273])^(a[49] & b[274])^(a[48] & b[275])^(a[47] & b[276])^(a[46] & b[277])^(a[45] & b[278])^(a[44] & b[279])^(a[43] & b[280])^(a[42] & b[281])^(a[41] & b[282])^(a[40] & b[283])^(a[39] & b[284])^(a[38] & b[285])^(a[37] & b[286])^(a[36] & b[287])^(a[35] & b[288])^(a[34] & b[289])^(a[33] & b[290])^(a[32] & b[291])^(a[31] & b[292])^(a[30] & b[293])^(a[29] & b[294])^(a[28] & b[295])^(a[27] & b[296])^(a[26] & b[297])^(a[25] & b[298])^(a[24] & b[299])^(a[23] & b[300])^(a[22] & b[301])^(a[21] & b[302])^(a[20] & b[303])^(a[19] & b[304])^(a[18] & b[305])^(a[17] & b[306])^(a[16] & b[307])^(a[15] & b[308])^(a[14] & b[309])^(a[13] & b[310])^(a[12] & b[311])^(a[11] & b[312])^(a[10] & b[313])^(a[9] & b[314])^(a[8] & b[315])^(a[7] & b[316])^(a[6] & b[317])^(a[5] & b[318])^(a[4] & b[319])^(a[3] & b[320])^(a[2] & b[321])^(a[1] & b[322])^(a[0] & b[323]);
assign y[324] = (a[324] & b[0])^(a[323] & b[1])^(a[322] & b[2])^(a[321] & b[3])^(a[320] & b[4])^(a[319] & b[5])^(a[318] & b[6])^(a[317] & b[7])^(a[316] & b[8])^(a[315] & b[9])^(a[314] & b[10])^(a[313] & b[11])^(a[312] & b[12])^(a[311] & b[13])^(a[310] & b[14])^(a[309] & b[15])^(a[308] & b[16])^(a[307] & b[17])^(a[306] & b[18])^(a[305] & b[19])^(a[304] & b[20])^(a[303] & b[21])^(a[302] & b[22])^(a[301] & b[23])^(a[300] & b[24])^(a[299] & b[25])^(a[298] & b[26])^(a[297] & b[27])^(a[296] & b[28])^(a[295] & b[29])^(a[294] & b[30])^(a[293] & b[31])^(a[292] & b[32])^(a[291] & b[33])^(a[290] & b[34])^(a[289] & b[35])^(a[288] & b[36])^(a[287] & b[37])^(a[286] & b[38])^(a[285] & b[39])^(a[284] & b[40])^(a[283] & b[41])^(a[282] & b[42])^(a[281] & b[43])^(a[280] & b[44])^(a[279] & b[45])^(a[278] & b[46])^(a[277] & b[47])^(a[276] & b[48])^(a[275] & b[49])^(a[274] & b[50])^(a[273] & b[51])^(a[272] & b[52])^(a[271] & b[53])^(a[270] & b[54])^(a[269] & b[55])^(a[268] & b[56])^(a[267] & b[57])^(a[266] & b[58])^(a[265] & b[59])^(a[264] & b[60])^(a[263] & b[61])^(a[262] & b[62])^(a[261] & b[63])^(a[260] & b[64])^(a[259] & b[65])^(a[258] & b[66])^(a[257] & b[67])^(a[256] & b[68])^(a[255] & b[69])^(a[254] & b[70])^(a[253] & b[71])^(a[252] & b[72])^(a[251] & b[73])^(a[250] & b[74])^(a[249] & b[75])^(a[248] & b[76])^(a[247] & b[77])^(a[246] & b[78])^(a[245] & b[79])^(a[244] & b[80])^(a[243] & b[81])^(a[242] & b[82])^(a[241] & b[83])^(a[240] & b[84])^(a[239] & b[85])^(a[238] & b[86])^(a[237] & b[87])^(a[236] & b[88])^(a[235] & b[89])^(a[234] & b[90])^(a[233] & b[91])^(a[232] & b[92])^(a[231] & b[93])^(a[230] & b[94])^(a[229] & b[95])^(a[228] & b[96])^(a[227] & b[97])^(a[226] & b[98])^(a[225] & b[99])^(a[224] & b[100])^(a[223] & b[101])^(a[222] & b[102])^(a[221] & b[103])^(a[220] & b[104])^(a[219] & b[105])^(a[218] & b[106])^(a[217] & b[107])^(a[216] & b[108])^(a[215] & b[109])^(a[214] & b[110])^(a[213] & b[111])^(a[212] & b[112])^(a[211] & b[113])^(a[210] & b[114])^(a[209] & b[115])^(a[208] & b[116])^(a[207] & b[117])^(a[206] & b[118])^(a[205] & b[119])^(a[204] & b[120])^(a[203] & b[121])^(a[202] & b[122])^(a[201] & b[123])^(a[200] & b[124])^(a[199] & b[125])^(a[198] & b[126])^(a[197] & b[127])^(a[196] & b[128])^(a[195] & b[129])^(a[194] & b[130])^(a[193] & b[131])^(a[192] & b[132])^(a[191] & b[133])^(a[190] & b[134])^(a[189] & b[135])^(a[188] & b[136])^(a[187] & b[137])^(a[186] & b[138])^(a[185] & b[139])^(a[184] & b[140])^(a[183] & b[141])^(a[182] & b[142])^(a[181] & b[143])^(a[180] & b[144])^(a[179] & b[145])^(a[178] & b[146])^(a[177] & b[147])^(a[176] & b[148])^(a[175] & b[149])^(a[174] & b[150])^(a[173] & b[151])^(a[172] & b[152])^(a[171] & b[153])^(a[170] & b[154])^(a[169] & b[155])^(a[168] & b[156])^(a[167] & b[157])^(a[166] & b[158])^(a[165] & b[159])^(a[164] & b[160])^(a[163] & b[161])^(a[162] & b[162])^(a[161] & b[163])^(a[160] & b[164])^(a[159] & b[165])^(a[158] & b[166])^(a[157] & b[167])^(a[156] & b[168])^(a[155] & b[169])^(a[154] & b[170])^(a[153] & b[171])^(a[152] & b[172])^(a[151] & b[173])^(a[150] & b[174])^(a[149] & b[175])^(a[148] & b[176])^(a[147] & b[177])^(a[146] & b[178])^(a[145] & b[179])^(a[144] & b[180])^(a[143] & b[181])^(a[142] & b[182])^(a[141] & b[183])^(a[140] & b[184])^(a[139] & b[185])^(a[138] & b[186])^(a[137] & b[187])^(a[136] & b[188])^(a[135] & b[189])^(a[134] & b[190])^(a[133] & b[191])^(a[132] & b[192])^(a[131] & b[193])^(a[130] & b[194])^(a[129] & b[195])^(a[128] & b[196])^(a[127] & b[197])^(a[126] & b[198])^(a[125] & b[199])^(a[124] & b[200])^(a[123] & b[201])^(a[122] & b[202])^(a[121] & b[203])^(a[120] & b[204])^(a[119] & b[205])^(a[118] & b[206])^(a[117] & b[207])^(a[116] & b[208])^(a[115] & b[209])^(a[114] & b[210])^(a[113] & b[211])^(a[112] & b[212])^(a[111] & b[213])^(a[110] & b[214])^(a[109] & b[215])^(a[108] & b[216])^(a[107] & b[217])^(a[106] & b[218])^(a[105] & b[219])^(a[104] & b[220])^(a[103] & b[221])^(a[102] & b[222])^(a[101] & b[223])^(a[100] & b[224])^(a[99] & b[225])^(a[98] & b[226])^(a[97] & b[227])^(a[96] & b[228])^(a[95] & b[229])^(a[94] & b[230])^(a[93] & b[231])^(a[92] & b[232])^(a[91] & b[233])^(a[90] & b[234])^(a[89] & b[235])^(a[88] & b[236])^(a[87] & b[237])^(a[86] & b[238])^(a[85] & b[239])^(a[84] & b[240])^(a[83] & b[241])^(a[82] & b[242])^(a[81] & b[243])^(a[80] & b[244])^(a[79] & b[245])^(a[78] & b[246])^(a[77] & b[247])^(a[76] & b[248])^(a[75] & b[249])^(a[74] & b[250])^(a[73] & b[251])^(a[72] & b[252])^(a[71] & b[253])^(a[70] & b[254])^(a[69] & b[255])^(a[68] & b[256])^(a[67] & b[257])^(a[66] & b[258])^(a[65] & b[259])^(a[64] & b[260])^(a[63] & b[261])^(a[62] & b[262])^(a[61] & b[263])^(a[60] & b[264])^(a[59] & b[265])^(a[58] & b[266])^(a[57] & b[267])^(a[56] & b[268])^(a[55] & b[269])^(a[54] & b[270])^(a[53] & b[271])^(a[52] & b[272])^(a[51] & b[273])^(a[50] & b[274])^(a[49] & b[275])^(a[48] & b[276])^(a[47] & b[277])^(a[46] & b[278])^(a[45] & b[279])^(a[44] & b[280])^(a[43] & b[281])^(a[42] & b[282])^(a[41] & b[283])^(a[40] & b[284])^(a[39] & b[285])^(a[38] & b[286])^(a[37] & b[287])^(a[36] & b[288])^(a[35] & b[289])^(a[34] & b[290])^(a[33] & b[291])^(a[32] & b[292])^(a[31] & b[293])^(a[30] & b[294])^(a[29] & b[295])^(a[28] & b[296])^(a[27] & b[297])^(a[26] & b[298])^(a[25] & b[299])^(a[24] & b[300])^(a[23] & b[301])^(a[22] & b[302])^(a[21] & b[303])^(a[20] & b[304])^(a[19] & b[305])^(a[18] & b[306])^(a[17] & b[307])^(a[16] & b[308])^(a[15] & b[309])^(a[14] & b[310])^(a[13] & b[311])^(a[12] & b[312])^(a[11] & b[313])^(a[10] & b[314])^(a[9] & b[315])^(a[8] & b[316])^(a[7] & b[317])^(a[6] & b[318])^(a[5] & b[319])^(a[4] & b[320])^(a[3] & b[321])^(a[2] & b[322])^(a[1] & b[323])^(a[0] & b[324]);
assign y[325] = (a[325] & b[0])^(a[324] & b[1])^(a[323] & b[2])^(a[322] & b[3])^(a[321] & b[4])^(a[320] & b[5])^(a[319] & b[6])^(a[318] & b[7])^(a[317] & b[8])^(a[316] & b[9])^(a[315] & b[10])^(a[314] & b[11])^(a[313] & b[12])^(a[312] & b[13])^(a[311] & b[14])^(a[310] & b[15])^(a[309] & b[16])^(a[308] & b[17])^(a[307] & b[18])^(a[306] & b[19])^(a[305] & b[20])^(a[304] & b[21])^(a[303] & b[22])^(a[302] & b[23])^(a[301] & b[24])^(a[300] & b[25])^(a[299] & b[26])^(a[298] & b[27])^(a[297] & b[28])^(a[296] & b[29])^(a[295] & b[30])^(a[294] & b[31])^(a[293] & b[32])^(a[292] & b[33])^(a[291] & b[34])^(a[290] & b[35])^(a[289] & b[36])^(a[288] & b[37])^(a[287] & b[38])^(a[286] & b[39])^(a[285] & b[40])^(a[284] & b[41])^(a[283] & b[42])^(a[282] & b[43])^(a[281] & b[44])^(a[280] & b[45])^(a[279] & b[46])^(a[278] & b[47])^(a[277] & b[48])^(a[276] & b[49])^(a[275] & b[50])^(a[274] & b[51])^(a[273] & b[52])^(a[272] & b[53])^(a[271] & b[54])^(a[270] & b[55])^(a[269] & b[56])^(a[268] & b[57])^(a[267] & b[58])^(a[266] & b[59])^(a[265] & b[60])^(a[264] & b[61])^(a[263] & b[62])^(a[262] & b[63])^(a[261] & b[64])^(a[260] & b[65])^(a[259] & b[66])^(a[258] & b[67])^(a[257] & b[68])^(a[256] & b[69])^(a[255] & b[70])^(a[254] & b[71])^(a[253] & b[72])^(a[252] & b[73])^(a[251] & b[74])^(a[250] & b[75])^(a[249] & b[76])^(a[248] & b[77])^(a[247] & b[78])^(a[246] & b[79])^(a[245] & b[80])^(a[244] & b[81])^(a[243] & b[82])^(a[242] & b[83])^(a[241] & b[84])^(a[240] & b[85])^(a[239] & b[86])^(a[238] & b[87])^(a[237] & b[88])^(a[236] & b[89])^(a[235] & b[90])^(a[234] & b[91])^(a[233] & b[92])^(a[232] & b[93])^(a[231] & b[94])^(a[230] & b[95])^(a[229] & b[96])^(a[228] & b[97])^(a[227] & b[98])^(a[226] & b[99])^(a[225] & b[100])^(a[224] & b[101])^(a[223] & b[102])^(a[222] & b[103])^(a[221] & b[104])^(a[220] & b[105])^(a[219] & b[106])^(a[218] & b[107])^(a[217] & b[108])^(a[216] & b[109])^(a[215] & b[110])^(a[214] & b[111])^(a[213] & b[112])^(a[212] & b[113])^(a[211] & b[114])^(a[210] & b[115])^(a[209] & b[116])^(a[208] & b[117])^(a[207] & b[118])^(a[206] & b[119])^(a[205] & b[120])^(a[204] & b[121])^(a[203] & b[122])^(a[202] & b[123])^(a[201] & b[124])^(a[200] & b[125])^(a[199] & b[126])^(a[198] & b[127])^(a[197] & b[128])^(a[196] & b[129])^(a[195] & b[130])^(a[194] & b[131])^(a[193] & b[132])^(a[192] & b[133])^(a[191] & b[134])^(a[190] & b[135])^(a[189] & b[136])^(a[188] & b[137])^(a[187] & b[138])^(a[186] & b[139])^(a[185] & b[140])^(a[184] & b[141])^(a[183] & b[142])^(a[182] & b[143])^(a[181] & b[144])^(a[180] & b[145])^(a[179] & b[146])^(a[178] & b[147])^(a[177] & b[148])^(a[176] & b[149])^(a[175] & b[150])^(a[174] & b[151])^(a[173] & b[152])^(a[172] & b[153])^(a[171] & b[154])^(a[170] & b[155])^(a[169] & b[156])^(a[168] & b[157])^(a[167] & b[158])^(a[166] & b[159])^(a[165] & b[160])^(a[164] & b[161])^(a[163] & b[162])^(a[162] & b[163])^(a[161] & b[164])^(a[160] & b[165])^(a[159] & b[166])^(a[158] & b[167])^(a[157] & b[168])^(a[156] & b[169])^(a[155] & b[170])^(a[154] & b[171])^(a[153] & b[172])^(a[152] & b[173])^(a[151] & b[174])^(a[150] & b[175])^(a[149] & b[176])^(a[148] & b[177])^(a[147] & b[178])^(a[146] & b[179])^(a[145] & b[180])^(a[144] & b[181])^(a[143] & b[182])^(a[142] & b[183])^(a[141] & b[184])^(a[140] & b[185])^(a[139] & b[186])^(a[138] & b[187])^(a[137] & b[188])^(a[136] & b[189])^(a[135] & b[190])^(a[134] & b[191])^(a[133] & b[192])^(a[132] & b[193])^(a[131] & b[194])^(a[130] & b[195])^(a[129] & b[196])^(a[128] & b[197])^(a[127] & b[198])^(a[126] & b[199])^(a[125] & b[200])^(a[124] & b[201])^(a[123] & b[202])^(a[122] & b[203])^(a[121] & b[204])^(a[120] & b[205])^(a[119] & b[206])^(a[118] & b[207])^(a[117] & b[208])^(a[116] & b[209])^(a[115] & b[210])^(a[114] & b[211])^(a[113] & b[212])^(a[112] & b[213])^(a[111] & b[214])^(a[110] & b[215])^(a[109] & b[216])^(a[108] & b[217])^(a[107] & b[218])^(a[106] & b[219])^(a[105] & b[220])^(a[104] & b[221])^(a[103] & b[222])^(a[102] & b[223])^(a[101] & b[224])^(a[100] & b[225])^(a[99] & b[226])^(a[98] & b[227])^(a[97] & b[228])^(a[96] & b[229])^(a[95] & b[230])^(a[94] & b[231])^(a[93] & b[232])^(a[92] & b[233])^(a[91] & b[234])^(a[90] & b[235])^(a[89] & b[236])^(a[88] & b[237])^(a[87] & b[238])^(a[86] & b[239])^(a[85] & b[240])^(a[84] & b[241])^(a[83] & b[242])^(a[82] & b[243])^(a[81] & b[244])^(a[80] & b[245])^(a[79] & b[246])^(a[78] & b[247])^(a[77] & b[248])^(a[76] & b[249])^(a[75] & b[250])^(a[74] & b[251])^(a[73] & b[252])^(a[72] & b[253])^(a[71] & b[254])^(a[70] & b[255])^(a[69] & b[256])^(a[68] & b[257])^(a[67] & b[258])^(a[66] & b[259])^(a[65] & b[260])^(a[64] & b[261])^(a[63] & b[262])^(a[62] & b[263])^(a[61] & b[264])^(a[60] & b[265])^(a[59] & b[266])^(a[58] & b[267])^(a[57] & b[268])^(a[56] & b[269])^(a[55] & b[270])^(a[54] & b[271])^(a[53] & b[272])^(a[52] & b[273])^(a[51] & b[274])^(a[50] & b[275])^(a[49] & b[276])^(a[48] & b[277])^(a[47] & b[278])^(a[46] & b[279])^(a[45] & b[280])^(a[44] & b[281])^(a[43] & b[282])^(a[42] & b[283])^(a[41] & b[284])^(a[40] & b[285])^(a[39] & b[286])^(a[38] & b[287])^(a[37] & b[288])^(a[36] & b[289])^(a[35] & b[290])^(a[34] & b[291])^(a[33] & b[292])^(a[32] & b[293])^(a[31] & b[294])^(a[30] & b[295])^(a[29] & b[296])^(a[28] & b[297])^(a[27] & b[298])^(a[26] & b[299])^(a[25] & b[300])^(a[24] & b[301])^(a[23] & b[302])^(a[22] & b[303])^(a[21] & b[304])^(a[20] & b[305])^(a[19] & b[306])^(a[18] & b[307])^(a[17] & b[308])^(a[16] & b[309])^(a[15] & b[310])^(a[14] & b[311])^(a[13] & b[312])^(a[12] & b[313])^(a[11] & b[314])^(a[10] & b[315])^(a[9] & b[316])^(a[8] & b[317])^(a[7] & b[318])^(a[6] & b[319])^(a[5] & b[320])^(a[4] & b[321])^(a[3] & b[322])^(a[2] & b[323])^(a[1] & b[324])^(a[0] & b[325]);
assign y[326] = (a[326] & b[0])^(a[325] & b[1])^(a[324] & b[2])^(a[323] & b[3])^(a[322] & b[4])^(a[321] & b[5])^(a[320] & b[6])^(a[319] & b[7])^(a[318] & b[8])^(a[317] & b[9])^(a[316] & b[10])^(a[315] & b[11])^(a[314] & b[12])^(a[313] & b[13])^(a[312] & b[14])^(a[311] & b[15])^(a[310] & b[16])^(a[309] & b[17])^(a[308] & b[18])^(a[307] & b[19])^(a[306] & b[20])^(a[305] & b[21])^(a[304] & b[22])^(a[303] & b[23])^(a[302] & b[24])^(a[301] & b[25])^(a[300] & b[26])^(a[299] & b[27])^(a[298] & b[28])^(a[297] & b[29])^(a[296] & b[30])^(a[295] & b[31])^(a[294] & b[32])^(a[293] & b[33])^(a[292] & b[34])^(a[291] & b[35])^(a[290] & b[36])^(a[289] & b[37])^(a[288] & b[38])^(a[287] & b[39])^(a[286] & b[40])^(a[285] & b[41])^(a[284] & b[42])^(a[283] & b[43])^(a[282] & b[44])^(a[281] & b[45])^(a[280] & b[46])^(a[279] & b[47])^(a[278] & b[48])^(a[277] & b[49])^(a[276] & b[50])^(a[275] & b[51])^(a[274] & b[52])^(a[273] & b[53])^(a[272] & b[54])^(a[271] & b[55])^(a[270] & b[56])^(a[269] & b[57])^(a[268] & b[58])^(a[267] & b[59])^(a[266] & b[60])^(a[265] & b[61])^(a[264] & b[62])^(a[263] & b[63])^(a[262] & b[64])^(a[261] & b[65])^(a[260] & b[66])^(a[259] & b[67])^(a[258] & b[68])^(a[257] & b[69])^(a[256] & b[70])^(a[255] & b[71])^(a[254] & b[72])^(a[253] & b[73])^(a[252] & b[74])^(a[251] & b[75])^(a[250] & b[76])^(a[249] & b[77])^(a[248] & b[78])^(a[247] & b[79])^(a[246] & b[80])^(a[245] & b[81])^(a[244] & b[82])^(a[243] & b[83])^(a[242] & b[84])^(a[241] & b[85])^(a[240] & b[86])^(a[239] & b[87])^(a[238] & b[88])^(a[237] & b[89])^(a[236] & b[90])^(a[235] & b[91])^(a[234] & b[92])^(a[233] & b[93])^(a[232] & b[94])^(a[231] & b[95])^(a[230] & b[96])^(a[229] & b[97])^(a[228] & b[98])^(a[227] & b[99])^(a[226] & b[100])^(a[225] & b[101])^(a[224] & b[102])^(a[223] & b[103])^(a[222] & b[104])^(a[221] & b[105])^(a[220] & b[106])^(a[219] & b[107])^(a[218] & b[108])^(a[217] & b[109])^(a[216] & b[110])^(a[215] & b[111])^(a[214] & b[112])^(a[213] & b[113])^(a[212] & b[114])^(a[211] & b[115])^(a[210] & b[116])^(a[209] & b[117])^(a[208] & b[118])^(a[207] & b[119])^(a[206] & b[120])^(a[205] & b[121])^(a[204] & b[122])^(a[203] & b[123])^(a[202] & b[124])^(a[201] & b[125])^(a[200] & b[126])^(a[199] & b[127])^(a[198] & b[128])^(a[197] & b[129])^(a[196] & b[130])^(a[195] & b[131])^(a[194] & b[132])^(a[193] & b[133])^(a[192] & b[134])^(a[191] & b[135])^(a[190] & b[136])^(a[189] & b[137])^(a[188] & b[138])^(a[187] & b[139])^(a[186] & b[140])^(a[185] & b[141])^(a[184] & b[142])^(a[183] & b[143])^(a[182] & b[144])^(a[181] & b[145])^(a[180] & b[146])^(a[179] & b[147])^(a[178] & b[148])^(a[177] & b[149])^(a[176] & b[150])^(a[175] & b[151])^(a[174] & b[152])^(a[173] & b[153])^(a[172] & b[154])^(a[171] & b[155])^(a[170] & b[156])^(a[169] & b[157])^(a[168] & b[158])^(a[167] & b[159])^(a[166] & b[160])^(a[165] & b[161])^(a[164] & b[162])^(a[163] & b[163])^(a[162] & b[164])^(a[161] & b[165])^(a[160] & b[166])^(a[159] & b[167])^(a[158] & b[168])^(a[157] & b[169])^(a[156] & b[170])^(a[155] & b[171])^(a[154] & b[172])^(a[153] & b[173])^(a[152] & b[174])^(a[151] & b[175])^(a[150] & b[176])^(a[149] & b[177])^(a[148] & b[178])^(a[147] & b[179])^(a[146] & b[180])^(a[145] & b[181])^(a[144] & b[182])^(a[143] & b[183])^(a[142] & b[184])^(a[141] & b[185])^(a[140] & b[186])^(a[139] & b[187])^(a[138] & b[188])^(a[137] & b[189])^(a[136] & b[190])^(a[135] & b[191])^(a[134] & b[192])^(a[133] & b[193])^(a[132] & b[194])^(a[131] & b[195])^(a[130] & b[196])^(a[129] & b[197])^(a[128] & b[198])^(a[127] & b[199])^(a[126] & b[200])^(a[125] & b[201])^(a[124] & b[202])^(a[123] & b[203])^(a[122] & b[204])^(a[121] & b[205])^(a[120] & b[206])^(a[119] & b[207])^(a[118] & b[208])^(a[117] & b[209])^(a[116] & b[210])^(a[115] & b[211])^(a[114] & b[212])^(a[113] & b[213])^(a[112] & b[214])^(a[111] & b[215])^(a[110] & b[216])^(a[109] & b[217])^(a[108] & b[218])^(a[107] & b[219])^(a[106] & b[220])^(a[105] & b[221])^(a[104] & b[222])^(a[103] & b[223])^(a[102] & b[224])^(a[101] & b[225])^(a[100] & b[226])^(a[99] & b[227])^(a[98] & b[228])^(a[97] & b[229])^(a[96] & b[230])^(a[95] & b[231])^(a[94] & b[232])^(a[93] & b[233])^(a[92] & b[234])^(a[91] & b[235])^(a[90] & b[236])^(a[89] & b[237])^(a[88] & b[238])^(a[87] & b[239])^(a[86] & b[240])^(a[85] & b[241])^(a[84] & b[242])^(a[83] & b[243])^(a[82] & b[244])^(a[81] & b[245])^(a[80] & b[246])^(a[79] & b[247])^(a[78] & b[248])^(a[77] & b[249])^(a[76] & b[250])^(a[75] & b[251])^(a[74] & b[252])^(a[73] & b[253])^(a[72] & b[254])^(a[71] & b[255])^(a[70] & b[256])^(a[69] & b[257])^(a[68] & b[258])^(a[67] & b[259])^(a[66] & b[260])^(a[65] & b[261])^(a[64] & b[262])^(a[63] & b[263])^(a[62] & b[264])^(a[61] & b[265])^(a[60] & b[266])^(a[59] & b[267])^(a[58] & b[268])^(a[57] & b[269])^(a[56] & b[270])^(a[55] & b[271])^(a[54] & b[272])^(a[53] & b[273])^(a[52] & b[274])^(a[51] & b[275])^(a[50] & b[276])^(a[49] & b[277])^(a[48] & b[278])^(a[47] & b[279])^(a[46] & b[280])^(a[45] & b[281])^(a[44] & b[282])^(a[43] & b[283])^(a[42] & b[284])^(a[41] & b[285])^(a[40] & b[286])^(a[39] & b[287])^(a[38] & b[288])^(a[37] & b[289])^(a[36] & b[290])^(a[35] & b[291])^(a[34] & b[292])^(a[33] & b[293])^(a[32] & b[294])^(a[31] & b[295])^(a[30] & b[296])^(a[29] & b[297])^(a[28] & b[298])^(a[27] & b[299])^(a[26] & b[300])^(a[25] & b[301])^(a[24] & b[302])^(a[23] & b[303])^(a[22] & b[304])^(a[21] & b[305])^(a[20] & b[306])^(a[19] & b[307])^(a[18] & b[308])^(a[17] & b[309])^(a[16] & b[310])^(a[15] & b[311])^(a[14] & b[312])^(a[13] & b[313])^(a[12] & b[314])^(a[11] & b[315])^(a[10] & b[316])^(a[9] & b[317])^(a[8] & b[318])^(a[7] & b[319])^(a[6] & b[320])^(a[5] & b[321])^(a[4] & b[322])^(a[3] & b[323])^(a[2] & b[324])^(a[1] & b[325])^(a[0] & b[326]);
assign y[327] = (a[327] & b[0])^(a[326] & b[1])^(a[325] & b[2])^(a[324] & b[3])^(a[323] & b[4])^(a[322] & b[5])^(a[321] & b[6])^(a[320] & b[7])^(a[319] & b[8])^(a[318] & b[9])^(a[317] & b[10])^(a[316] & b[11])^(a[315] & b[12])^(a[314] & b[13])^(a[313] & b[14])^(a[312] & b[15])^(a[311] & b[16])^(a[310] & b[17])^(a[309] & b[18])^(a[308] & b[19])^(a[307] & b[20])^(a[306] & b[21])^(a[305] & b[22])^(a[304] & b[23])^(a[303] & b[24])^(a[302] & b[25])^(a[301] & b[26])^(a[300] & b[27])^(a[299] & b[28])^(a[298] & b[29])^(a[297] & b[30])^(a[296] & b[31])^(a[295] & b[32])^(a[294] & b[33])^(a[293] & b[34])^(a[292] & b[35])^(a[291] & b[36])^(a[290] & b[37])^(a[289] & b[38])^(a[288] & b[39])^(a[287] & b[40])^(a[286] & b[41])^(a[285] & b[42])^(a[284] & b[43])^(a[283] & b[44])^(a[282] & b[45])^(a[281] & b[46])^(a[280] & b[47])^(a[279] & b[48])^(a[278] & b[49])^(a[277] & b[50])^(a[276] & b[51])^(a[275] & b[52])^(a[274] & b[53])^(a[273] & b[54])^(a[272] & b[55])^(a[271] & b[56])^(a[270] & b[57])^(a[269] & b[58])^(a[268] & b[59])^(a[267] & b[60])^(a[266] & b[61])^(a[265] & b[62])^(a[264] & b[63])^(a[263] & b[64])^(a[262] & b[65])^(a[261] & b[66])^(a[260] & b[67])^(a[259] & b[68])^(a[258] & b[69])^(a[257] & b[70])^(a[256] & b[71])^(a[255] & b[72])^(a[254] & b[73])^(a[253] & b[74])^(a[252] & b[75])^(a[251] & b[76])^(a[250] & b[77])^(a[249] & b[78])^(a[248] & b[79])^(a[247] & b[80])^(a[246] & b[81])^(a[245] & b[82])^(a[244] & b[83])^(a[243] & b[84])^(a[242] & b[85])^(a[241] & b[86])^(a[240] & b[87])^(a[239] & b[88])^(a[238] & b[89])^(a[237] & b[90])^(a[236] & b[91])^(a[235] & b[92])^(a[234] & b[93])^(a[233] & b[94])^(a[232] & b[95])^(a[231] & b[96])^(a[230] & b[97])^(a[229] & b[98])^(a[228] & b[99])^(a[227] & b[100])^(a[226] & b[101])^(a[225] & b[102])^(a[224] & b[103])^(a[223] & b[104])^(a[222] & b[105])^(a[221] & b[106])^(a[220] & b[107])^(a[219] & b[108])^(a[218] & b[109])^(a[217] & b[110])^(a[216] & b[111])^(a[215] & b[112])^(a[214] & b[113])^(a[213] & b[114])^(a[212] & b[115])^(a[211] & b[116])^(a[210] & b[117])^(a[209] & b[118])^(a[208] & b[119])^(a[207] & b[120])^(a[206] & b[121])^(a[205] & b[122])^(a[204] & b[123])^(a[203] & b[124])^(a[202] & b[125])^(a[201] & b[126])^(a[200] & b[127])^(a[199] & b[128])^(a[198] & b[129])^(a[197] & b[130])^(a[196] & b[131])^(a[195] & b[132])^(a[194] & b[133])^(a[193] & b[134])^(a[192] & b[135])^(a[191] & b[136])^(a[190] & b[137])^(a[189] & b[138])^(a[188] & b[139])^(a[187] & b[140])^(a[186] & b[141])^(a[185] & b[142])^(a[184] & b[143])^(a[183] & b[144])^(a[182] & b[145])^(a[181] & b[146])^(a[180] & b[147])^(a[179] & b[148])^(a[178] & b[149])^(a[177] & b[150])^(a[176] & b[151])^(a[175] & b[152])^(a[174] & b[153])^(a[173] & b[154])^(a[172] & b[155])^(a[171] & b[156])^(a[170] & b[157])^(a[169] & b[158])^(a[168] & b[159])^(a[167] & b[160])^(a[166] & b[161])^(a[165] & b[162])^(a[164] & b[163])^(a[163] & b[164])^(a[162] & b[165])^(a[161] & b[166])^(a[160] & b[167])^(a[159] & b[168])^(a[158] & b[169])^(a[157] & b[170])^(a[156] & b[171])^(a[155] & b[172])^(a[154] & b[173])^(a[153] & b[174])^(a[152] & b[175])^(a[151] & b[176])^(a[150] & b[177])^(a[149] & b[178])^(a[148] & b[179])^(a[147] & b[180])^(a[146] & b[181])^(a[145] & b[182])^(a[144] & b[183])^(a[143] & b[184])^(a[142] & b[185])^(a[141] & b[186])^(a[140] & b[187])^(a[139] & b[188])^(a[138] & b[189])^(a[137] & b[190])^(a[136] & b[191])^(a[135] & b[192])^(a[134] & b[193])^(a[133] & b[194])^(a[132] & b[195])^(a[131] & b[196])^(a[130] & b[197])^(a[129] & b[198])^(a[128] & b[199])^(a[127] & b[200])^(a[126] & b[201])^(a[125] & b[202])^(a[124] & b[203])^(a[123] & b[204])^(a[122] & b[205])^(a[121] & b[206])^(a[120] & b[207])^(a[119] & b[208])^(a[118] & b[209])^(a[117] & b[210])^(a[116] & b[211])^(a[115] & b[212])^(a[114] & b[213])^(a[113] & b[214])^(a[112] & b[215])^(a[111] & b[216])^(a[110] & b[217])^(a[109] & b[218])^(a[108] & b[219])^(a[107] & b[220])^(a[106] & b[221])^(a[105] & b[222])^(a[104] & b[223])^(a[103] & b[224])^(a[102] & b[225])^(a[101] & b[226])^(a[100] & b[227])^(a[99] & b[228])^(a[98] & b[229])^(a[97] & b[230])^(a[96] & b[231])^(a[95] & b[232])^(a[94] & b[233])^(a[93] & b[234])^(a[92] & b[235])^(a[91] & b[236])^(a[90] & b[237])^(a[89] & b[238])^(a[88] & b[239])^(a[87] & b[240])^(a[86] & b[241])^(a[85] & b[242])^(a[84] & b[243])^(a[83] & b[244])^(a[82] & b[245])^(a[81] & b[246])^(a[80] & b[247])^(a[79] & b[248])^(a[78] & b[249])^(a[77] & b[250])^(a[76] & b[251])^(a[75] & b[252])^(a[74] & b[253])^(a[73] & b[254])^(a[72] & b[255])^(a[71] & b[256])^(a[70] & b[257])^(a[69] & b[258])^(a[68] & b[259])^(a[67] & b[260])^(a[66] & b[261])^(a[65] & b[262])^(a[64] & b[263])^(a[63] & b[264])^(a[62] & b[265])^(a[61] & b[266])^(a[60] & b[267])^(a[59] & b[268])^(a[58] & b[269])^(a[57] & b[270])^(a[56] & b[271])^(a[55] & b[272])^(a[54] & b[273])^(a[53] & b[274])^(a[52] & b[275])^(a[51] & b[276])^(a[50] & b[277])^(a[49] & b[278])^(a[48] & b[279])^(a[47] & b[280])^(a[46] & b[281])^(a[45] & b[282])^(a[44] & b[283])^(a[43] & b[284])^(a[42] & b[285])^(a[41] & b[286])^(a[40] & b[287])^(a[39] & b[288])^(a[38] & b[289])^(a[37] & b[290])^(a[36] & b[291])^(a[35] & b[292])^(a[34] & b[293])^(a[33] & b[294])^(a[32] & b[295])^(a[31] & b[296])^(a[30] & b[297])^(a[29] & b[298])^(a[28] & b[299])^(a[27] & b[300])^(a[26] & b[301])^(a[25] & b[302])^(a[24] & b[303])^(a[23] & b[304])^(a[22] & b[305])^(a[21] & b[306])^(a[20] & b[307])^(a[19] & b[308])^(a[18] & b[309])^(a[17] & b[310])^(a[16] & b[311])^(a[15] & b[312])^(a[14] & b[313])^(a[13] & b[314])^(a[12] & b[315])^(a[11] & b[316])^(a[10] & b[317])^(a[9] & b[318])^(a[8] & b[319])^(a[7] & b[320])^(a[6] & b[321])^(a[5] & b[322])^(a[4] & b[323])^(a[3] & b[324])^(a[2] & b[325])^(a[1] & b[326])^(a[0] & b[327]);
assign y[328] = (a[328] & b[0])^(a[327] & b[1])^(a[326] & b[2])^(a[325] & b[3])^(a[324] & b[4])^(a[323] & b[5])^(a[322] & b[6])^(a[321] & b[7])^(a[320] & b[8])^(a[319] & b[9])^(a[318] & b[10])^(a[317] & b[11])^(a[316] & b[12])^(a[315] & b[13])^(a[314] & b[14])^(a[313] & b[15])^(a[312] & b[16])^(a[311] & b[17])^(a[310] & b[18])^(a[309] & b[19])^(a[308] & b[20])^(a[307] & b[21])^(a[306] & b[22])^(a[305] & b[23])^(a[304] & b[24])^(a[303] & b[25])^(a[302] & b[26])^(a[301] & b[27])^(a[300] & b[28])^(a[299] & b[29])^(a[298] & b[30])^(a[297] & b[31])^(a[296] & b[32])^(a[295] & b[33])^(a[294] & b[34])^(a[293] & b[35])^(a[292] & b[36])^(a[291] & b[37])^(a[290] & b[38])^(a[289] & b[39])^(a[288] & b[40])^(a[287] & b[41])^(a[286] & b[42])^(a[285] & b[43])^(a[284] & b[44])^(a[283] & b[45])^(a[282] & b[46])^(a[281] & b[47])^(a[280] & b[48])^(a[279] & b[49])^(a[278] & b[50])^(a[277] & b[51])^(a[276] & b[52])^(a[275] & b[53])^(a[274] & b[54])^(a[273] & b[55])^(a[272] & b[56])^(a[271] & b[57])^(a[270] & b[58])^(a[269] & b[59])^(a[268] & b[60])^(a[267] & b[61])^(a[266] & b[62])^(a[265] & b[63])^(a[264] & b[64])^(a[263] & b[65])^(a[262] & b[66])^(a[261] & b[67])^(a[260] & b[68])^(a[259] & b[69])^(a[258] & b[70])^(a[257] & b[71])^(a[256] & b[72])^(a[255] & b[73])^(a[254] & b[74])^(a[253] & b[75])^(a[252] & b[76])^(a[251] & b[77])^(a[250] & b[78])^(a[249] & b[79])^(a[248] & b[80])^(a[247] & b[81])^(a[246] & b[82])^(a[245] & b[83])^(a[244] & b[84])^(a[243] & b[85])^(a[242] & b[86])^(a[241] & b[87])^(a[240] & b[88])^(a[239] & b[89])^(a[238] & b[90])^(a[237] & b[91])^(a[236] & b[92])^(a[235] & b[93])^(a[234] & b[94])^(a[233] & b[95])^(a[232] & b[96])^(a[231] & b[97])^(a[230] & b[98])^(a[229] & b[99])^(a[228] & b[100])^(a[227] & b[101])^(a[226] & b[102])^(a[225] & b[103])^(a[224] & b[104])^(a[223] & b[105])^(a[222] & b[106])^(a[221] & b[107])^(a[220] & b[108])^(a[219] & b[109])^(a[218] & b[110])^(a[217] & b[111])^(a[216] & b[112])^(a[215] & b[113])^(a[214] & b[114])^(a[213] & b[115])^(a[212] & b[116])^(a[211] & b[117])^(a[210] & b[118])^(a[209] & b[119])^(a[208] & b[120])^(a[207] & b[121])^(a[206] & b[122])^(a[205] & b[123])^(a[204] & b[124])^(a[203] & b[125])^(a[202] & b[126])^(a[201] & b[127])^(a[200] & b[128])^(a[199] & b[129])^(a[198] & b[130])^(a[197] & b[131])^(a[196] & b[132])^(a[195] & b[133])^(a[194] & b[134])^(a[193] & b[135])^(a[192] & b[136])^(a[191] & b[137])^(a[190] & b[138])^(a[189] & b[139])^(a[188] & b[140])^(a[187] & b[141])^(a[186] & b[142])^(a[185] & b[143])^(a[184] & b[144])^(a[183] & b[145])^(a[182] & b[146])^(a[181] & b[147])^(a[180] & b[148])^(a[179] & b[149])^(a[178] & b[150])^(a[177] & b[151])^(a[176] & b[152])^(a[175] & b[153])^(a[174] & b[154])^(a[173] & b[155])^(a[172] & b[156])^(a[171] & b[157])^(a[170] & b[158])^(a[169] & b[159])^(a[168] & b[160])^(a[167] & b[161])^(a[166] & b[162])^(a[165] & b[163])^(a[164] & b[164])^(a[163] & b[165])^(a[162] & b[166])^(a[161] & b[167])^(a[160] & b[168])^(a[159] & b[169])^(a[158] & b[170])^(a[157] & b[171])^(a[156] & b[172])^(a[155] & b[173])^(a[154] & b[174])^(a[153] & b[175])^(a[152] & b[176])^(a[151] & b[177])^(a[150] & b[178])^(a[149] & b[179])^(a[148] & b[180])^(a[147] & b[181])^(a[146] & b[182])^(a[145] & b[183])^(a[144] & b[184])^(a[143] & b[185])^(a[142] & b[186])^(a[141] & b[187])^(a[140] & b[188])^(a[139] & b[189])^(a[138] & b[190])^(a[137] & b[191])^(a[136] & b[192])^(a[135] & b[193])^(a[134] & b[194])^(a[133] & b[195])^(a[132] & b[196])^(a[131] & b[197])^(a[130] & b[198])^(a[129] & b[199])^(a[128] & b[200])^(a[127] & b[201])^(a[126] & b[202])^(a[125] & b[203])^(a[124] & b[204])^(a[123] & b[205])^(a[122] & b[206])^(a[121] & b[207])^(a[120] & b[208])^(a[119] & b[209])^(a[118] & b[210])^(a[117] & b[211])^(a[116] & b[212])^(a[115] & b[213])^(a[114] & b[214])^(a[113] & b[215])^(a[112] & b[216])^(a[111] & b[217])^(a[110] & b[218])^(a[109] & b[219])^(a[108] & b[220])^(a[107] & b[221])^(a[106] & b[222])^(a[105] & b[223])^(a[104] & b[224])^(a[103] & b[225])^(a[102] & b[226])^(a[101] & b[227])^(a[100] & b[228])^(a[99] & b[229])^(a[98] & b[230])^(a[97] & b[231])^(a[96] & b[232])^(a[95] & b[233])^(a[94] & b[234])^(a[93] & b[235])^(a[92] & b[236])^(a[91] & b[237])^(a[90] & b[238])^(a[89] & b[239])^(a[88] & b[240])^(a[87] & b[241])^(a[86] & b[242])^(a[85] & b[243])^(a[84] & b[244])^(a[83] & b[245])^(a[82] & b[246])^(a[81] & b[247])^(a[80] & b[248])^(a[79] & b[249])^(a[78] & b[250])^(a[77] & b[251])^(a[76] & b[252])^(a[75] & b[253])^(a[74] & b[254])^(a[73] & b[255])^(a[72] & b[256])^(a[71] & b[257])^(a[70] & b[258])^(a[69] & b[259])^(a[68] & b[260])^(a[67] & b[261])^(a[66] & b[262])^(a[65] & b[263])^(a[64] & b[264])^(a[63] & b[265])^(a[62] & b[266])^(a[61] & b[267])^(a[60] & b[268])^(a[59] & b[269])^(a[58] & b[270])^(a[57] & b[271])^(a[56] & b[272])^(a[55] & b[273])^(a[54] & b[274])^(a[53] & b[275])^(a[52] & b[276])^(a[51] & b[277])^(a[50] & b[278])^(a[49] & b[279])^(a[48] & b[280])^(a[47] & b[281])^(a[46] & b[282])^(a[45] & b[283])^(a[44] & b[284])^(a[43] & b[285])^(a[42] & b[286])^(a[41] & b[287])^(a[40] & b[288])^(a[39] & b[289])^(a[38] & b[290])^(a[37] & b[291])^(a[36] & b[292])^(a[35] & b[293])^(a[34] & b[294])^(a[33] & b[295])^(a[32] & b[296])^(a[31] & b[297])^(a[30] & b[298])^(a[29] & b[299])^(a[28] & b[300])^(a[27] & b[301])^(a[26] & b[302])^(a[25] & b[303])^(a[24] & b[304])^(a[23] & b[305])^(a[22] & b[306])^(a[21] & b[307])^(a[20] & b[308])^(a[19] & b[309])^(a[18] & b[310])^(a[17] & b[311])^(a[16] & b[312])^(a[15] & b[313])^(a[14] & b[314])^(a[13] & b[315])^(a[12] & b[316])^(a[11] & b[317])^(a[10] & b[318])^(a[9] & b[319])^(a[8] & b[320])^(a[7] & b[321])^(a[6] & b[322])^(a[5] & b[323])^(a[4] & b[324])^(a[3] & b[325])^(a[2] & b[326])^(a[1] & b[327])^(a[0] & b[328]);
assign y[329] = (a[329] & b[0])^(a[328] & b[1])^(a[327] & b[2])^(a[326] & b[3])^(a[325] & b[4])^(a[324] & b[5])^(a[323] & b[6])^(a[322] & b[7])^(a[321] & b[8])^(a[320] & b[9])^(a[319] & b[10])^(a[318] & b[11])^(a[317] & b[12])^(a[316] & b[13])^(a[315] & b[14])^(a[314] & b[15])^(a[313] & b[16])^(a[312] & b[17])^(a[311] & b[18])^(a[310] & b[19])^(a[309] & b[20])^(a[308] & b[21])^(a[307] & b[22])^(a[306] & b[23])^(a[305] & b[24])^(a[304] & b[25])^(a[303] & b[26])^(a[302] & b[27])^(a[301] & b[28])^(a[300] & b[29])^(a[299] & b[30])^(a[298] & b[31])^(a[297] & b[32])^(a[296] & b[33])^(a[295] & b[34])^(a[294] & b[35])^(a[293] & b[36])^(a[292] & b[37])^(a[291] & b[38])^(a[290] & b[39])^(a[289] & b[40])^(a[288] & b[41])^(a[287] & b[42])^(a[286] & b[43])^(a[285] & b[44])^(a[284] & b[45])^(a[283] & b[46])^(a[282] & b[47])^(a[281] & b[48])^(a[280] & b[49])^(a[279] & b[50])^(a[278] & b[51])^(a[277] & b[52])^(a[276] & b[53])^(a[275] & b[54])^(a[274] & b[55])^(a[273] & b[56])^(a[272] & b[57])^(a[271] & b[58])^(a[270] & b[59])^(a[269] & b[60])^(a[268] & b[61])^(a[267] & b[62])^(a[266] & b[63])^(a[265] & b[64])^(a[264] & b[65])^(a[263] & b[66])^(a[262] & b[67])^(a[261] & b[68])^(a[260] & b[69])^(a[259] & b[70])^(a[258] & b[71])^(a[257] & b[72])^(a[256] & b[73])^(a[255] & b[74])^(a[254] & b[75])^(a[253] & b[76])^(a[252] & b[77])^(a[251] & b[78])^(a[250] & b[79])^(a[249] & b[80])^(a[248] & b[81])^(a[247] & b[82])^(a[246] & b[83])^(a[245] & b[84])^(a[244] & b[85])^(a[243] & b[86])^(a[242] & b[87])^(a[241] & b[88])^(a[240] & b[89])^(a[239] & b[90])^(a[238] & b[91])^(a[237] & b[92])^(a[236] & b[93])^(a[235] & b[94])^(a[234] & b[95])^(a[233] & b[96])^(a[232] & b[97])^(a[231] & b[98])^(a[230] & b[99])^(a[229] & b[100])^(a[228] & b[101])^(a[227] & b[102])^(a[226] & b[103])^(a[225] & b[104])^(a[224] & b[105])^(a[223] & b[106])^(a[222] & b[107])^(a[221] & b[108])^(a[220] & b[109])^(a[219] & b[110])^(a[218] & b[111])^(a[217] & b[112])^(a[216] & b[113])^(a[215] & b[114])^(a[214] & b[115])^(a[213] & b[116])^(a[212] & b[117])^(a[211] & b[118])^(a[210] & b[119])^(a[209] & b[120])^(a[208] & b[121])^(a[207] & b[122])^(a[206] & b[123])^(a[205] & b[124])^(a[204] & b[125])^(a[203] & b[126])^(a[202] & b[127])^(a[201] & b[128])^(a[200] & b[129])^(a[199] & b[130])^(a[198] & b[131])^(a[197] & b[132])^(a[196] & b[133])^(a[195] & b[134])^(a[194] & b[135])^(a[193] & b[136])^(a[192] & b[137])^(a[191] & b[138])^(a[190] & b[139])^(a[189] & b[140])^(a[188] & b[141])^(a[187] & b[142])^(a[186] & b[143])^(a[185] & b[144])^(a[184] & b[145])^(a[183] & b[146])^(a[182] & b[147])^(a[181] & b[148])^(a[180] & b[149])^(a[179] & b[150])^(a[178] & b[151])^(a[177] & b[152])^(a[176] & b[153])^(a[175] & b[154])^(a[174] & b[155])^(a[173] & b[156])^(a[172] & b[157])^(a[171] & b[158])^(a[170] & b[159])^(a[169] & b[160])^(a[168] & b[161])^(a[167] & b[162])^(a[166] & b[163])^(a[165] & b[164])^(a[164] & b[165])^(a[163] & b[166])^(a[162] & b[167])^(a[161] & b[168])^(a[160] & b[169])^(a[159] & b[170])^(a[158] & b[171])^(a[157] & b[172])^(a[156] & b[173])^(a[155] & b[174])^(a[154] & b[175])^(a[153] & b[176])^(a[152] & b[177])^(a[151] & b[178])^(a[150] & b[179])^(a[149] & b[180])^(a[148] & b[181])^(a[147] & b[182])^(a[146] & b[183])^(a[145] & b[184])^(a[144] & b[185])^(a[143] & b[186])^(a[142] & b[187])^(a[141] & b[188])^(a[140] & b[189])^(a[139] & b[190])^(a[138] & b[191])^(a[137] & b[192])^(a[136] & b[193])^(a[135] & b[194])^(a[134] & b[195])^(a[133] & b[196])^(a[132] & b[197])^(a[131] & b[198])^(a[130] & b[199])^(a[129] & b[200])^(a[128] & b[201])^(a[127] & b[202])^(a[126] & b[203])^(a[125] & b[204])^(a[124] & b[205])^(a[123] & b[206])^(a[122] & b[207])^(a[121] & b[208])^(a[120] & b[209])^(a[119] & b[210])^(a[118] & b[211])^(a[117] & b[212])^(a[116] & b[213])^(a[115] & b[214])^(a[114] & b[215])^(a[113] & b[216])^(a[112] & b[217])^(a[111] & b[218])^(a[110] & b[219])^(a[109] & b[220])^(a[108] & b[221])^(a[107] & b[222])^(a[106] & b[223])^(a[105] & b[224])^(a[104] & b[225])^(a[103] & b[226])^(a[102] & b[227])^(a[101] & b[228])^(a[100] & b[229])^(a[99] & b[230])^(a[98] & b[231])^(a[97] & b[232])^(a[96] & b[233])^(a[95] & b[234])^(a[94] & b[235])^(a[93] & b[236])^(a[92] & b[237])^(a[91] & b[238])^(a[90] & b[239])^(a[89] & b[240])^(a[88] & b[241])^(a[87] & b[242])^(a[86] & b[243])^(a[85] & b[244])^(a[84] & b[245])^(a[83] & b[246])^(a[82] & b[247])^(a[81] & b[248])^(a[80] & b[249])^(a[79] & b[250])^(a[78] & b[251])^(a[77] & b[252])^(a[76] & b[253])^(a[75] & b[254])^(a[74] & b[255])^(a[73] & b[256])^(a[72] & b[257])^(a[71] & b[258])^(a[70] & b[259])^(a[69] & b[260])^(a[68] & b[261])^(a[67] & b[262])^(a[66] & b[263])^(a[65] & b[264])^(a[64] & b[265])^(a[63] & b[266])^(a[62] & b[267])^(a[61] & b[268])^(a[60] & b[269])^(a[59] & b[270])^(a[58] & b[271])^(a[57] & b[272])^(a[56] & b[273])^(a[55] & b[274])^(a[54] & b[275])^(a[53] & b[276])^(a[52] & b[277])^(a[51] & b[278])^(a[50] & b[279])^(a[49] & b[280])^(a[48] & b[281])^(a[47] & b[282])^(a[46] & b[283])^(a[45] & b[284])^(a[44] & b[285])^(a[43] & b[286])^(a[42] & b[287])^(a[41] & b[288])^(a[40] & b[289])^(a[39] & b[290])^(a[38] & b[291])^(a[37] & b[292])^(a[36] & b[293])^(a[35] & b[294])^(a[34] & b[295])^(a[33] & b[296])^(a[32] & b[297])^(a[31] & b[298])^(a[30] & b[299])^(a[29] & b[300])^(a[28] & b[301])^(a[27] & b[302])^(a[26] & b[303])^(a[25] & b[304])^(a[24] & b[305])^(a[23] & b[306])^(a[22] & b[307])^(a[21] & b[308])^(a[20] & b[309])^(a[19] & b[310])^(a[18] & b[311])^(a[17] & b[312])^(a[16] & b[313])^(a[15] & b[314])^(a[14] & b[315])^(a[13] & b[316])^(a[12] & b[317])^(a[11] & b[318])^(a[10] & b[319])^(a[9] & b[320])^(a[8] & b[321])^(a[7] & b[322])^(a[6] & b[323])^(a[5] & b[324])^(a[4] & b[325])^(a[3] & b[326])^(a[2] & b[327])^(a[1] & b[328])^(a[0] & b[329]);
assign y[330] = (a[330] & b[0])^(a[329] & b[1])^(a[328] & b[2])^(a[327] & b[3])^(a[326] & b[4])^(a[325] & b[5])^(a[324] & b[6])^(a[323] & b[7])^(a[322] & b[8])^(a[321] & b[9])^(a[320] & b[10])^(a[319] & b[11])^(a[318] & b[12])^(a[317] & b[13])^(a[316] & b[14])^(a[315] & b[15])^(a[314] & b[16])^(a[313] & b[17])^(a[312] & b[18])^(a[311] & b[19])^(a[310] & b[20])^(a[309] & b[21])^(a[308] & b[22])^(a[307] & b[23])^(a[306] & b[24])^(a[305] & b[25])^(a[304] & b[26])^(a[303] & b[27])^(a[302] & b[28])^(a[301] & b[29])^(a[300] & b[30])^(a[299] & b[31])^(a[298] & b[32])^(a[297] & b[33])^(a[296] & b[34])^(a[295] & b[35])^(a[294] & b[36])^(a[293] & b[37])^(a[292] & b[38])^(a[291] & b[39])^(a[290] & b[40])^(a[289] & b[41])^(a[288] & b[42])^(a[287] & b[43])^(a[286] & b[44])^(a[285] & b[45])^(a[284] & b[46])^(a[283] & b[47])^(a[282] & b[48])^(a[281] & b[49])^(a[280] & b[50])^(a[279] & b[51])^(a[278] & b[52])^(a[277] & b[53])^(a[276] & b[54])^(a[275] & b[55])^(a[274] & b[56])^(a[273] & b[57])^(a[272] & b[58])^(a[271] & b[59])^(a[270] & b[60])^(a[269] & b[61])^(a[268] & b[62])^(a[267] & b[63])^(a[266] & b[64])^(a[265] & b[65])^(a[264] & b[66])^(a[263] & b[67])^(a[262] & b[68])^(a[261] & b[69])^(a[260] & b[70])^(a[259] & b[71])^(a[258] & b[72])^(a[257] & b[73])^(a[256] & b[74])^(a[255] & b[75])^(a[254] & b[76])^(a[253] & b[77])^(a[252] & b[78])^(a[251] & b[79])^(a[250] & b[80])^(a[249] & b[81])^(a[248] & b[82])^(a[247] & b[83])^(a[246] & b[84])^(a[245] & b[85])^(a[244] & b[86])^(a[243] & b[87])^(a[242] & b[88])^(a[241] & b[89])^(a[240] & b[90])^(a[239] & b[91])^(a[238] & b[92])^(a[237] & b[93])^(a[236] & b[94])^(a[235] & b[95])^(a[234] & b[96])^(a[233] & b[97])^(a[232] & b[98])^(a[231] & b[99])^(a[230] & b[100])^(a[229] & b[101])^(a[228] & b[102])^(a[227] & b[103])^(a[226] & b[104])^(a[225] & b[105])^(a[224] & b[106])^(a[223] & b[107])^(a[222] & b[108])^(a[221] & b[109])^(a[220] & b[110])^(a[219] & b[111])^(a[218] & b[112])^(a[217] & b[113])^(a[216] & b[114])^(a[215] & b[115])^(a[214] & b[116])^(a[213] & b[117])^(a[212] & b[118])^(a[211] & b[119])^(a[210] & b[120])^(a[209] & b[121])^(a[208] & b[122])^(a[207] & b[123])^(a[206] & b[124])^(a[205] & b[125])^(a[204] & b[126])^(a[203] & b[127])^(a[202] & b[128])^(a[201] & b[129])^(a[200] & b[130])^(a[199] & b[131])^(a[198] & b[132])^(a[197] & b[133])^(a[196] & b[134])^(a[195] & b[135])^(a[194] & b[136])^(a[193] & b[137])^(a[192] & b[138])^(a[191] & b[139])^(a[190] & b[140])^(a[189] & b[141])^(a[188] & b[142])^(a[187] & b[143])^(a[186] & b[144])^(a[185] & b[145])^(a[184] & b[146])^(a[183] & b[147])^(a[182] & b[148])^(a[181] & b[149])^(a[180] & b[150])^(a[179] & b[151])^(a[178] & b[152])^(a[177] & b[153])^(a[176] & b[154])^(a[175] & b[155])^(a[174] & b[156])^(a[173] & b[157])^(a[172] & b[158])^(a[171] & b[159])^(a[170] & b[160])^(a[169] & b[161])^(a[168] & b[162])^(a[167] & b[163])^(a[166] & b[164])^(a[165] & b[165])^(a[164] & b[166])^(a[163] & b[167])^(a[162] & b[168])^(a[161] & b[169])^(a[160] & b[170])^(a[159] & b[171])^(a[158] & b[172])^(a[157] & b[173])^(a[156] & b[174])^(a[155] & b[175])^(a[154] & b[176])^(a[153] & b[177])^(a[152] & b[178])^(a[151] & b[179])^(a[150] & b[180])^(a[149] & b[181])^(a[148] & b[182])^(a[147] & b[183])^(a[146] & b[184])^(a[145] & b[185])^(a[144] & b[186])^(a[143] & b[187])^(a[142] & b[188])^(a[141] & b[189])^(a[140] & b[190])^(a[139] & b[191])^(a[138] & b[192])^(a[137] & b[193])^(a[136] & b[194])^(a[135] & b[195])^(a[134] & b[196])^(a[133] & b[197])^(a[132] & b[198])^(a[131] & b[199])^(a[130] & b[200])^(a[129] & b[201])^(a[128] & b[202])^(a[127] & b[203])^(a[126] & b[204])^(a[125] & b[205])^(a[124] & b[206])^(a[123] & b[207])^(a[122] & b[208])^(a[121] & b[209])^(a[120] & b[210])^(a[119] & b[211])^(a[118] & b[212])^(a[117] & b[213])^(a[116] & b[214])^(a[115] & b[215])^(a[114] & b[216])^(a[113] & b[217])^(a[112] & b[218])^(a[111] & b[219])^(a[110] & b[220])^(a[109] & b[221])^(a[108] & b[222])^(a[107] & b[223])^(a[106] & b[224])^(a[105] & b[225])^(a[104] & b[226])^(a[103] & b[227])^(a[102] & b[228])^(a[101] & b[229])^(a[100] & b[230])^(a[99] & b[231])^(a[98] & b[232])^(a[97] & b[233])^(a[96] & b[234])^(a[95] & b[235])^(a[94] & b[236])^(a[93] & b[237])^(a[92] & b[238])^(a[91] & b[239])^(a[90] & b[240])^(a[89] & b[241])^(a[88] & b[242])^(a[87] & b[243])^(a[86] & b[244])^(a[85] & b[245])^(a[84] & b[246])^(a[83] & b[247])^(a[82] & b[248])^(a[81] & b[249])^(a[80] & b[250])^(a[79] & b[251])^(a[78] & b[252])^(a[77] & b[253])^(a[76] & b[254])^(a[75] & b[255])^(a[74] & b[256])^(a[73] & b[257])^(a[72] & b[258])^(a[71] & b[259])^(a[70] & b[260])^(a[69] & b[261])^(a[68] & b[262])^(a[67] & b[263])^(a[66] & b[264])^(a[65] & b[265])^(a[64] & b[266])^(a[63] & b[267])^(a[62] & b[268])^(a[61] & b[269])^(a[60] & b[270])^(a[59] & b[271])^(a[58] & b[272])^(a[57] & b[273])^(a[56] & b[274])^(a[55] & b[275])^(a[54] & b[276])^(a[53] & b[277])^(a[52] & b[278])^(a[51] & b[279])^(a[50] & b[280])^(a[49] & b[281])^(a[48] & b[282])^(a[47] & b[283])^(a[46] & b[284])^(a[45] & b[285])^(a[44] & b[286])^(a[43] & b[287])^(a[42] & b[288])^(a[41] & b[289])^(a[40] & b[290])^(a[39] & b[291])^(a[38] & b[292])^(a[37] & b[293])^(a[36] & b[294])^(a[35] & b[295])^(a[34] & b[296])^(a[33] & b[297])^(a[32] & b[298])^(a[31] & b[299])^(a[30] & b[300])^(a[29] & b[301])^(a[28] & b[302])^(a[27] & b[303])^(a[26] & b[304])^(a[25] & b[305])^(a[24] & b[306])^(a[23] & b[307])^(a[22] & b[308])^(a[21] & b[309])^(a[20] & b[310])^(a[19] & b[311])^(a[18] & b[312])^(a[17] & b[313])^(a[16] & b[314])^(a[15] & b[315])^(a[14] & b[316])^(a[13] & b[317])^(a[12] & b[318])^(a[11] & b[319])^(a[10] & b[320])^(a[9] & b[321])^(a[8] & b[322])^(a[7] & b[323])^(a[6] & b[324])^(a[5] & b[325])^(a[4] & b[326])^(a[3] & b[327])^(a[2] & b[328])^(a[1] & b[329])^(a[0] & b[330]);
assign y[331] = (a[331] & b[0])^(a[330] & b[1])^(a[329] & b[2])^(a[328] & b[3])^(a[327] & b[4])^(a[326] & b[5])^(a[325] & b[6])^(a[324] & b[7])^(a[323] & b[8])^(a[322] & b[9])^(a[321] & b[10])^(a[320] & b[11])^(a[319] & b[12])^(a[318] & b[13])^(a[317] & b[14])^(a[316] & b[15])^(a[315] & b[16])^(a[314] & b[17])^(a[313] & b[18])^(a[312] & b[19])^(a[311] & b[20])^(a[310] & b[21])^(a[309] & b[22])^(a[308] & b[23])^(a[307] & b[24])^(a[306] & b[25])^(a[305] & b[26])^(a[304] & b[27])^(a[303] & b[28])^(a[302] & b[29])^(a[301] & b[30])^(a[300] & b[31])^(a[299] & b[32])^(a[298] & b[33])^(a[297] & b[34])^(a[296] & b[35])^(a[295] & b[36])^(a[294] & b[37])^(a[293] & b[38])^(a[292] & b[39])^(a[291] & b[40])^(a[290] & b[41])^(a[289] & b[42])^(a[288] & b[43])^(a[287] & b[44])^(a[286] & b[45])^(a[285] & b[46])^(a[284] & b[47])^(a[283] & b[48])^(a[282] & b[49])^(a[281] & b[50])^(a[280] & b[51])^(a[279] & b[52])^(a[278] & b[53])^(a[277] & b[54])^(a[276] & b[55])^(a[275] & b[56])^(a[274] & b[57])^(a[273] & b[58])^(a[272] & b[59])^(a[271] & b[60])^(a[270] & b[61])^(a[269] & b[62])^(a[268] & b[63])^(a[267] & b[64])^(a[266] & b[65])^(a[265] & b[66])^(a[264] & b[67])^(a[263] & b[68])^(a[262] & b[69])^(a[261] & b[70])^(a[260] & b[71])^(a[259] & b[72])^(a[258] & b[73])^(a[257] & b[74])^(a[256] & b[75])^(a[255] & b[76])^(a[254] & b[77])^(a[253] & b[78])^(a[252] & b[79])^(a[251] & b[80])^(a[250] & b[81])^(a[249] & b[82])^(a[248] & b[83])^(a[247] & b[84])^(a[246] & b[85])^(a[245] & b[86])^(a[244] & b[87])^(a[243] & b[88])^(a[242] & b[89])^(a[241] & b[90])^(a[240] & b[91])^(a[239] & b[92])^(a[238] & b[93])^(a[237] & b[94])^(a[236] & b[95])^(a[235] & b[96])^(a[234] & b[97])^(a[233] & b[98])^(a[232] & b[99])^(a[231] & b[100])^(a[230] & b[101])^(a[229] & b[102])^(a[228] & b[103])^(a[227] & b[104])^(a[226] & b[105])^(a[225] & b[106])^(a[224] & b[107])^(a[223] & b[108])^(a[222] & b[109])^(a[221] & b[110])^(a[220] & b[111])^(a[219] & b[112])^(a[218] & b[113])^(a[217] & b[114])^(a[216] & b[115])^(a[215] & b[116])^(a[214] & b[117])^(a[213] & b[118])^(a[212] & b[119])^(a[211] & b[120])^(a[210] & b[121])^(a[209] & b[122])^(a[208] & b[123])^(a[207] & b[124])^(a[206] & b[125])^(a[205] & b[126])^(a[204] & b[127])^(a[203] & b[128])^(a[202] & b[129])^(a[201] & b[130])^(a[200] & b[131])^(a[199] & b[132])^(a[198] & b[133])^(a[197] & b[134])^(a[196] & b[135])^(a[195] & b[136])^(a[194] & b[137])^(a[193] & b[138])^(a[192] & b[139])^(a[191] & b[140])^(a[190] & b[141])^(a[189] & b[142])^(a[188] & b[143])^(a[187] & b[144])^(a[186] & b[145])^(a[185] & b[146])^(a[184] & b[147])^(a[183] & b[148])^(a[182] & b[149])^(a[181] & b[150])^(a[180] & b[151])^(a[179] & b[152])^(a[178] & b[153])^(a[177] & b[154])^(a[176] & b[155])^(a[175] & b[156])^(a[174] & b[157])^(a[173] & b[158])^(a[172] & b[159])^(a[171] & b[160])^(a[170] & b[161])^(a[169] & b[162])^(a[168] & b[163])^(a[167] & b[164])^(a[166] & b[165])^(a[165] & b[166])^(a[164] & b[167])^(a[163] & b[168])^(a[162] & b[169])^(a[161] & b[170])^(a[160] & b[171])^(a[159] & b[172])^(a[158] & b[173])^(a[157] & b[174])^(a[156] & b[175])^(a[155] & b[176])^(a[154] & b[177])^(a[153] & b[178])^(a[152] & b[179])^(a[151] & b[180])^(a[150] & b[181])^(a[149] & b[182])^(a[148] & b[183])^(a[147] & b[184])^(a[146] & b[185])^(a[145] & b[186])^(a[144] & b[187])^(a[143] & b[188])^(a[142] & b[189])^(a[141] & b[190])^(a[140] & b[191])^(a[139] & b[192])^(a[138] & b[193])^(a[137] & b[194])^(a[136] & b[195])^(a[135] & b[196])^(a[134] & b[197])^(a[133] & b[198])^(a[132] & b[199])^(a[131] & b[200])^(a[130] & b[201])^(a[129] & b[202])^(a[128] & b[203])^(a[127] & b[204])^(a[126] & b[205])^(a[125] & b[206])^(a[124] & b[207])^(a[123] & b[208])^(a[122] & b[209])^(a[121] & b[210])^(a[120] & b[211])^(a[119] & b[212])^(a[118] & b[213])^(a[117] & b[214])^(a[116] & b[215])^(a[115] & b[216])^(a[114] & b[217])^(a[113] & b[218])^(a[112] & b[219])^(a[111] & b[220])^(a[110] & b[221])^(a[109] & b[222])^(a[108] & b[223])^(a[107] & b[224])^(a[106] & b[225])^(a[105] & b[226])^(a[104] & b[227])^(a[103] & b[228])^(a[102] & b[229])^(a[101] & b[230])^(a[100] & b[231])^(a[99] & b[232])^(a[98] & b[233])^(a[97] & b[234])^(a[96] & b[235])^(a[95] & b[236])^(a[94] & b[237])^(a[93] & b[238])^(a[92] & b[239])^(a[91] & b[240])^(a[90] & b[241])^(a[89] & b[242])^(a[88] & b[243])^(a[87] & b[244])^(a[86] & b[245])^(a[85] & b[246])^(a[84] & b[247])^(a[83] & b[248])^(a[82] & b[249])^(a[81] & b[250])^(a[80] & b[251])^(a[79] & b[252])^(a[78] & b[253])^(a[77] & b[254])^(a[76] & b[255])^(a[75] & b[256])^(a[74] & b[257])^(a[73] & b[258])^(a[72] & b[259])^(a[71] & b[260])^(a[70] & b[261])^(a[69] & b[262])^(a[68] & b[263])^(a[67] & b[264])^(a[66] & b[265])^(a[65] & b[266])^(a[64] & b[267])^(a[63] & b[268])^(a[62] & b[269])^(a[61] & b[270])^(a[60] & b[271])^(a[59] & b[272])^(a[58] & b[273])^(a[57] & b[274])^(a[56] & b[275])^(a[55] & b[276])^(a[54] & b[277])^(a[53] & b[278])^(a[52] & b[279])^(a[51] & b[280])^(a[50] & b[281])^(a[49] & b[282])^(a[48] & b[283])^(a[47] & b[284])^(a[46] & b[285])^(a[45] & b[286])^(a[44] & b[287])^(a[43] & b[288])^(a[42] & b[289])^(a[41] & b[290])^(a[40] & b[291])^(a[39] & b[292])^(a[38] & b[293])^(a[37] & b[294])^(a[36] & b[295])^(a[35] & b[296])^(a[34] & b[297])^(a[33] & b[298])^(a[32] & b[299])^(a[31] & b[300])^(a[30] & b[301])^(a[29] & b[302])^(a[28] & b[303])^(a[27] & b[304])^(a[26] & b[305])^(a[25] & b[306])^(a[24] & b[307])^(a[23] & b[308])^(a[22] & b[309])^(a[21] & b[310])^(a[20] & b[311])^(a[19] & b[312])^(a[18] & b[313])^(a[17] & b[314])^(a[16] & b[315])^(a[15] & b[316])^(a[14] & b[317])^(a[13] & b[318])^(a[12] & b[319])^(a[11] & b[320])^(a[10] & b[321])^(a[9] & b[322])^(a[8] & b[323])^(a[7] & b[324])^(a[6] & b[325])^(a[5] & b[326])^(a[4] & b[327])^(a[3] & b[328])^(a[2] & b[329])^(a[1] & b[330])^(a[0] & b[331]);
assign y[332] = (a[332] & b[0])^(a[331] & b[1])^(a[330] & b[2])^(a[329] & b[3])^(a[328] & b[4])^(a[327] & b[5])^(a[326] & b[6])^(a[325] & b[7])^(a[324] & b[8])^(a[323] & b[9])^(a[322] & b[10])^(a[321] & b[11])^(a[320] & b[12])^(a[319] & b[13])^(a[318] & b[14])^(a[317] & b[15])^(a[316] & b[16])^(a[315] & b[17])^(a[314] & b[18])^(a[313] & b[19])^(a[312] & b[20])^(a[311] & b[21])^(a[310] & b[22])^(a[309] & b[23])^(a[308] & b[24])^(a[307] & b[25])^(a[306] & b[26])^(a[305] & b[27])^(a[304] & b[28])^(a[303] & b[29])^(a[302] & b[30])^(a[301] & b[31])^(a[300] & b[32])^(a[299] & b[33])^(a[298] & b[34])^(a[297] & b[35])^(a[296] & b[36])^(a[295] & b[37])^(a[294] & b[38])^(a[293] & b[39])^(a[292] & b[40])^(a[291] & b[41])^(a[290] & b[42])^(a[289] & b[43])^(a[288] & b[44])^(a[287] & b[45])^(a[286] & b[46])^(a[285] & b[47])^(a[284] & b[48])^(a[283] & b[49])^(a[282] & b[50])^(a[281] & b[51])^(a[280] & b[52])^(a[279] & b[53])^(a[278] & b[54])^(a[277] & b[55])^(a[276] & b[56])^(a[275] & b[57])^(a[274] & b[58])^(a[273] & b[59])^(a[272] & b[60])^(a[271] & b[61])^(a[270] & b[62])^(a[269] & b[63])^(a[268] & b[64])^(a[267] & b[65])^(a[266] & b[66])^(a[265] & b[67])^(a[264] & b[68])^(a[263] & b[69])^(a[262] & b[70])^(a[261] & b[71])^(a[260] & b[72])^(a[259] & b[73])^(a[258] & b[74])^(a[257] & b[75])^(a[256] & b[76])^(a[255] & b[77])^(a[254] & b[78])^(a[253] & b[79])^(a[252] & b[80])^(a[251] & b[81])^(a[250] & b[82])^(a[249] & b[83])^(a[248] & b[84])^(a[247] & b[85])^(a[246] & b[86])^(a[245] & b[87])^(a[244] & b[88])^(a[243] & b[89])^(a[242] & b[90])^(a[241] & b[91])^(a[240] & b[92])^(a[239] & b[93])^(a[238] & b[94])^(a[237] & b[95])^(a[236] & b[96])^(a[235] & b[97])^(a[234] & b[98])^(a[233] & b[99])^(a[232] & b[100])^(a[231] & b[101])^(a[230] & b[102])^(a[229] & b[103])^(a[228] & b[104])^(a[227] & b[105])^(a[226] & b[106])^(a[225] & b[107])^(a[224] & b[108])^(a[223] & b[109])^(a[222] & b[110])^(a[221] & b[111])^(a[220] & b[112])^(a[219] & b[113])^(a[218] & b[114])^(a[217] & b[115])^(a[216] & b[116])^(a[215] & b[117])^(a[214] & b[118])^(a[213] & b[119])^(a[212] & b[120])^(a[211] & b[121])^(a[210] & b[122])^(a[209] & b[123])^(a[208] & b[124])^(a[207] & b[125])^(a[206] & b[126])^(a[205] & b[127])^(a[204] & b[128])^(a[203] & b[129])^(a[202] & b[130])^(a[201] & b[131])^(a[200] & b[132])^(a[199] & b[133])^(a[198] & b[134])^(a[197] & b[135])^(a[196] & b[136])^(a[195] & b[137])^(a[194] & b[138])^(a[193] & b[139])^(a[192] & b[140])^(a[191] & b[141])^(a[190] & b[142])^(a[189] & b[143])^(a[188] & b[144])^(a[187] & b[145])^(a[186] & b[146])^(a[185] & b[147])^(a[184] & b[148])^(a[183] & b[149])^(a[182] & b[150])^(a[181] & b[151])^(a[180] & b[152])^(a[179] & b[153])^(a[178] & b[154])^(a[177] & b[155])^(a[176] & b[156])^(a[175] & b[157])^(a[174] & b[158])^(a[173] & b[159])^(a[172] & b[160])^(a[171] & b[161])^(a[170] & b[162])^(a[169] & b[163])^(a[168] & b[164])^(a[167] & b[165])^(a[166] & b[166])^(a[165] & b[167])^(a[164] & b[168])^(a[163] & b[169])^(a[162] & b[170])^(a[161] & b[171])^(a[160] & b[172])^(a[159] & b[173])^(a[158] & b[174])^(a[157] & b[175])^(a[156] & b[176])^(a[155] & b[177])^(a[154] & b[178])^(a[153] & b[179])^(a[152] & b[180])^(a[151] & b[181])^(a[150] & b[182])^(a[149] & b[183])^(a[148] & b[184])^(a[147] & b[185])^(a[146] & b[186])^(a[145] & b[187])^(a[144] & b[188])^(a[143] & b[189])^(a[142] & b[190])^(a[141] & b[191])^(a[140] & b[192])^(a[139] & b[193])^(a[138] & b[194])^(a[137] & b[195])^(a[136] & b[196])^(a[135] & b[197])^(a[134] & b[198])^(a[133] & b[199])^(a[132] & b[200])^(a[131] & b[201])^(a[130] & b[202])^(a[129] & b[203])^(a[128] & b[204])^(a[127] & b[205])^(a[126] & b[206])^(a[125] & b[207])^(a[124] & b[208])^(a[123] & b[209])^(a[122] & b[210])^(a[121] & b[211])^(a[120] & b[212])^(a[119] & b[213])^(a[118] & b[214])^(a[117] & b[215])^(a[116] & b[216])^(a[115] & b[217])^(a[114] & b[218])^(a[113] & b[219])^(a[112] & b[220])^(a[111] & b[221])^(a[110] & b[222])^(a[109] & b[223])^(a[108] & b[224])^(a[107] & b[225])^(a[106] & b[226])^(a[105] & b[227])^(a[104] & b[228])^(a[103] & b[229])^(a[102] & b[230])^(a[101] & b[231])^(a[100] & b[232])^(a[99] & b[233])^(a[98] & b[234])^(a[97] & b[235])^(a[96] & b[236])^(a[95] & b[237])^(a[94] & b[238])^(a[93] & b[239])^(a[92] & b[240])^(a[91] & b[241])^(a[90] & b[242])^(a[89] & b[243])^(a[88] & b[244])^(a[87] & b[245])^(a[86] & b[246])^(a[85] & b[247])^(a[84] & b[248])^(a[83] & b[249])^(a[82] & b[250])^(a[81] & b[251])^(a[80] & b[252])^(a[79] & b[253])^(a[78] & b[254])^(a[77] & b[255])^(a[76] & b[256])^(a[75] & b[257])^(a[74] & b[258])^(a[73] & b[259])^(a[72] & b[260])^(a[71] & b[261])^(a[70] & b[262])^(a[69] & b[263])^(a[68] & b[264])^(a[67] & b[265])^(a[66] & b[266])^(a[65] & b[267])^(a[64] & b[268])^(a[63] & b[269])^(a[62] & b[270])^(a[61] & b[271])^(a[60] & b[272])^(a[59] & b[273])^(a[58] & b[274])^(a[57] & b[275])^(a[56] & b[276])^(a[55] & b[277])^(a[54] & b[278])^(a[53] & b[279])^(a[52] & b[280])^(a[51] & b[281])^(a[50] & b[282])^(a[49] & b[283])^(a[48] & b[284])^(a[47] & b[285])^(a[46] & b[286])^(a[45] & b[287])^(a[44] & b[288])^(a[43] & b[289])^(a[42] & b[290])^(a[41] & b[291])^(a[40] & b[292])^(a[39] & b[293])^(a[38] & b[294])^(a[37] & b[295])^(a[36] & b[296])^(a[35] & b[297])^(a[34] & b[298])^(a[33] & b[299])^(a[32] & b[300])^(a[31] & b[301])^(a[30] & b[302])^(a[29] & b[303])^(a[28] & b[304])^(a[27] & b[305])^(a[26] & b[306])^(a[25] & b[307])^(a[24] & b[308])^(a[23] & b[309])^(a[22] & b[310])^(a[21] & b[311])^(a[20] & b[312])^(a[19] & b[313])^(a[18] & b[314])^(a[17] & b[315])^(a[16] & b[316])^(a[15] & b[317])^(a[14] & b[318])^(a[13] & b[319])^(a[12] & b[320])^(a[11] & b[321])^(a[10] & b[322])^(a[9] & b[323])^(a[8] & b[324])^(a[7] & b[325])^(a[6] & b[326])^(a[5] & b[327])^(a[4] & b[328])^(a[3] & b[329])^(a[2] & b[330])^(a[1] & b[331])^(a[0] & b[332]);
assign y[333] = (a[333] & b[0])^(a[332] & b[1])^(a[331] & b[2])^(a[330] & b[3])^(a[329] & b[4])^(a[328] & b[5])^(a[327] & b[6])^(a[326] & b[7])^(a[325] & b[8])^(a[324] & b[9])^(a[323] & b[10])^(a[322] & b[11])^(a[321] & b[12])^(a[320] & b[13])^(a[319] & b[14])^(a[318] & b[15])^(a[317] & b[16])^(a[316] & b[17])^(a[315] & b[18])^(a[314] & b[19])^(a[313] & b[20])^(a[312] & b[21])^(a[311] & b[22])^(a[310] & b[23])^(a[309] & b[24])^(a[308] & b[25])^(a[307] & b[26])^(a[306] & b[27])^(a[305] & b[28])^(a[304] & b[29])^(a[303] & b[30])^(a[302] & b[31])^(a[301] & b[32])^(a[300] & b[33])^(a[299] & b[34])^(a[298] & b[35])^(a[297] & b[36])^(a[296] & b[37])^(a[295] & b[38])^(a[294] & b[39])^(a[293] & b[40])^(a[292] & b[41])^(a[291] & b[42])^(a[290] & b[43])^(a[289] & b[44])^(a[288] & b[45])^(a[287] & b[46])^(a[286] & b[47])^(a[285] & b[48])^(a[284] & b[49])^(a[283] & b[50])^(a[282] & b[51])^(a[281] & b[52])^(a[280] & b[53])^(a[279] & b[54])^(a[278] & b[55])^(a[277] & b[56])^(a[276] & b[57])^(a[275] & b[58])^(a[274] & b[59])^(a[273] & b[60])^(a[272] & b[61])^(a[271] & b[62])^(a[270] & b[63])^(a[269] & b[64])^(a[268] & b[65])^(a[267] & b[66])^(a[266] & b[67])^(a[265] & b[68])^(a[264] & b[69])^(a[263] & b[70])^(a[262] & b[71])^(a[261] & b[72])^(a[260] & b[73])^(a[259] & b[74])^(a[258] & b[75])^(a[257] & b[76])^(a[256] & b[77])^(a[255] & b[78])^(a[254] & b[79])^(a[253] & b[80])^(a[252] & b[81])^(a[251] & b[82])^(a[250] & b[83])^(a[249] & b[84])^(a[248] & b[85])^(a[247] & b[86])^(a[246] & b[87])^(a[245] & b[88])^(a[244] & b[89])^(a[243] & b[90])^(a[242] & b[91])^(a[241] & b[92])^(a[240] & b[93])^(a[239] & b[94])^(a[238] & b[95])^(a[237] & b[96])^(a[236] & b[97])^(a[235] & b[98])^(a[234] & b[99])^(a[233] & b[100])^(a[232] & b[101])^(a[231] & b[102])^(a[230] & b[103])^(a[229] & b[104])^(a[228] & b[105])^(a[227] & b[106])^(a[226] & b[107])^(a[225] & b[108])^(a[224] & b[109])^(a[223] & b[110])^(a[222] & b[111])^(a[221] & b[112])^(a[220] & b[113])^(a[219] & b[114])^(a[218] & b[115])^(a[217] & b[116])^(a[216] & b[117])^(a[215] & b[118])^(a[214] & b[119])^(a[213] & b[120])^(a[212] & b[121])^(a[211] & b[122])^(a[210] & b[123])^(a[209] & b[124])^(a[208] & b[125])^(a[207] & b[126])^(a[206] & b[127])^(a[205] & b[128])^(a[204] & b[129])^(a[203] & b[130])^(a[202] & b[131])^(a[201] & b[132])^(a[200] & b[133])^(a[199] & b[134])^(a[198] & b[135])^(a[197] & b[136])^(a[196] & b[137])^(a[195] & b[138])^(a[194] & b[139])^(a[193] & b[140])^(a[192] & b[141])^(a[191] & b[142])^(a[190] & b[143])^(a[189] & b[144])^(a[188] & b[145])^(a[187] & b[146])^(a[186] & b[147])^(a[185] & b[148])^(a[184] & b[149])^(a[183] & b[150])^(a[182] & b[151])^(a[181] & b[152])^(a[180] & b[153])^(a[179] & b[154])^(a[178] & b[155])^(a[177] & b[156])^(a[176] & b[157])^(a[175] & b[158])^(a[174] & b[159])^(a[173] & b[160])^(a[172] & b[161])^(a[171] & b[162])^(a[170] & b[163])^(a[169] & b[164])^(a[168] & b[165])^(a[167] & b[166])^(a[166] & b[167])^(a[165] & b[168])^(a[164] & b[169])^(a[163] & b[170])^(a[162] & b[171])^(a[161] & b[172])^(a[160] & b[173])^(a[159] & b[174])^(a[158] & b[175])^(a[157] & b[176])^(a[156] & b[177])^(a[155] & b[178])^(a[154] & b[179])^(a[153] & b[180])^(a[152] & b[181])^(a[151] & b[182])^(a[150] & b[183])^(a[149] & b[184])^(a[148] & b[185])^(a[147] & b[186])^(a[146] & b[187])^(a[145] & b[188])^(a[144] & b[189])^(a[143] & b[190])^(a[142] & b[191])^(a[141] & b[192])^(a[140] & b[193])^(a[139] & b[194])^(a[138] & b[195])^(a[137] & b[196])^(a[136] & b[197])^(a[135] & b[198])^(a[134] & b[199])^(a[133] & b[200])^(a[132] & b[201])^(a[131] & b[202])^(a[130] & b[203])^(a[129] & b[204])^(a[128] & b[205])^(a[127] & b[206])^(a[126] & b[207])^(a[125] & b[208])^(a[124] & b[209])^(a[123] & b[210])^(a[122] & b[211])^(a[121] & b[212])^(a[120] & b[213])^(a[119] & b[214])^(a[118] & b[215])^(a[117] & b[216])^(a[116] & b[217])^(a[115] & b[218])^(a[114] & b[219])^(a[113] & b[220])^(a[112] & b[221])^(a[111] & b[222])^(a[110] & b[223])^(a[109] & b[224])^(a[108] & b[225])^(a[107] & b[226])^(a[106] & b[227])^(a[105] & b[228])^(a[104] & b[229])^(a[103] & b[230])^(a[102] & b[231])^(a[101] & b[232])^(a[100] & b[233])^(a[99] & b[234])^(a[98] & b[235])^(a[97] & b[236])^(a[96] & b[237])^(a[95] & b[238])^(a[94] & b[239])^(a[93] & b[240])^(a[92] & b[241])^(a[91] & b[242])^(a[90] & b[243])^(a[89] & b[244])^(a[88] & b[245])^(a[87] & b[246])^(a[86] & b[247])^(a[85] & b[248])^(a[84] & b[249])^(a[83] & b[250])^(a[82] & b[251])^(a[81] & b[252])^(a[80] & b[253])^(a[79] & b[254])^(a[78] & b[255])^(a[77] & b[256])^(a[76] & b[257])^(a[75] & b[258])^(a[74] & b[259])^(a[73] & b[260])^(a[72] & b[261])^(a[71] & b[262])^(a[70] & b[263])^(a[69] & b[264])^(a[68] & b[265])^(a[67] & b[266])^(a[66] & b[267])^(a[65] & b[268])^(a[64] & b[269])^(a[63] & b[270])^(a[62] & b[271])^(a[61] & b[272])^(a[60] & b[273])^(a[59] & b[274])^(a[58] & b[275])^(a[57] & b[276])^(a[56] & b[277])^(a[55] & b[278])^(a[54] & b[279])^(a[53] & b[280])^(a[52] & b[281])^(a[51] & b[282])^(a[50] & b[283])^(a[49] & b[284])^(a[48] & b[285])^(a[47] & b[286])^(a[46] & b[287])^(a[45] & b[288])^(a[44] & b[289])^(a[43] & b[290])^(a[42] & b[291])^(a[41] & b[292])^(a[40] & b[293])^(a[39] & b[294])^(a[38] & b[295])^(a[37] & b[296])^(a[36] & b[297])^(a[35] & b[298])^(a[34] & b[299])^(a[33] & b[300])^(a[32] & b[301])^(a[31] & b[302])^(a[30] & b[303])^(a[29] & b[304])^(a[28] & b[305])^(a[27] & b[306])^(a[26] & b[307])^(a[25] & b[308])^(a[24] & b[309])^(a[23] & b[310])^(a[22] & b[311])^(a[21] & b[312])^(a[20] & b[313])^(a[19] & b[314])^(a[18] & b[315])^(a[17] & b[316])^(a[16] & b[317])^(a[15] & b[318])^(a[14] & b[319])^(a[13] & b[320])^(a[12] & b[321])^(a[11] & b[322])^(a[10] & b[323])^(a[9] & b[324])^(a[8] & b[325])^(a[7] & b[326])^(a[6] & b[327])^(a[5] & b[328])^(a[4] & b[329])^(a[3] & b[330])^(a[2] & b[331])^(a[1] & b[332])^(a[0] & b[333]);
assign y[334] = (a[334] & b[0])^(a[333] & b[1])^(a[332] & b[2])^(a[331] & b[3])^(a[330] & b[4])^(a[329] & b[5])^(a[328] & b[6])^(a[327] & b[7])^(a[326] & b[8])^(a[325] & b[9])^(a[324] & b[10])^(a[323] & b[11])^(a[322] & b[12])^(a[321] & b[13])^(a[320] & b[14])^(a[319] & b[15])^(a[318] & b[16])^(a[317] & b[17])^(a[316] & b[18])^(a[315] & b[19])^(a[314] & b[20])^(a[313] & b[21])^(a[312] & b[22])^(a[311] & b[23])^(a[310] & b[24])^(a[309] & b[25])^(a[308] & b[26])^(a[307] & b[27])^(a[306] & b[28])^(a[305] & b[29])^(a[304] & b[30])^(a[303] & b[31])^(a[302] & b[32])^(a[301] & b[33])^(a[300] & b[34])^(a[299] & b[35])^(a[298] & b[36])^(a[297] & b[37])^(a[296] & b[38])^(a[295] & b[39])^(a[294] & b[40])^(a[293] & b[41])^(a[292] & b[42])^(a[291] & b[43])^(a[290] & b[44])^(a[289] & b[45])^(a[288] & b[46])^(a[287] & b[47])^(a[286] & b[48])^(a[285] & b[49])^(a[284] & b[50])^(a[283] & b[51])^(a[282] & b[52])^(a[281] & b[53])^(a[280] & b[54])^(a[279] & b[55])^(a[278] & b[56])^(a[277] & b[57])^(a[276] & b[58])^(a[275] & b[59])^(a[274] & b[60])^(a[273] & b[61])^(a[272] & b[62])^(a[271] & b[63])^(a[270] & b[64])^(a[269] & b[65])^(a[268] & b[66])^(a[267] & b[67])^(a[266] & b[68])^(a[265] & b[69])^(a[264] & b[70])^(a[263] & b[71])^(a[262] & b[72])^(a[261] & b[73])^(a[260] & b[74])^(a[259] & b[75])^(a[258] & b[76])^(a[257] & b[77])^(a[256] & b[78])^(a[255] & b[79])^(a[254] & b[80])^(a[253] & b[81])^(a[252] & b[82])^(a[251] & b[83])^(a[250] & b[84])^(a[249] & b[85])^(a[248] & b[86])^(a[247] & b[87])^(a[246] & b[88])^(a[245] & b[89])^(a[244] & b[90])^(a[243] & b[91])^(a[242] & b[92])^(a[241] & b[93])^(a[240] & b[94])^(a[239] & b[95])^(a[238] & b[96])^(a[237] & b[97])^(a[236] & b[98])^(a[235] & b[99])^(a[234] & b[100])^(a[233] & b[101])^(a[232] & b[102])^(a[231] & b[103])^(a[230] & b[104])^(a[229] & b[105])^(a[228] & b[106])^(a[227] & b[107])^(a[226] & b[108])^(a[225] & b[109])^(a[224] & b[110])^(a[223] & b[111])^(a[222] & b[112])^(a[221] & b[113])^(a[220] & b[114])^(a[219] & b[115])^(a[218] & b[116])^(a[217] & b[117])^(a[216] & b[118])^(a[215] & b[119])^(a[214] & b[120])^(a[213] & b[121])^(a[212] & b[122])^(a[211] & b[123])^(a[210] & b[124])^(a[209] & b[125])^(a[208] & b[126])^(a[207] & b[127])^(a[206] & b[128])^(a[205] & b[129])^(a[204] & b[130])^(a[203] & b[131])^(a[202] & b[132])^(a[201] & b[133])^(a[200] & b[134])^(a[199] & b[135])^(a[198] & b[136])^(a[197] & b[137])^(a[196] & b[138])^(a[195] & b[139])^(a[194] & b[140])^(a[193] & b[141])^(a[192] & b[142])^(a[191] & b[143])^(a[190] & b[144])^(a[189] & b[145])^(a[188] & b[146])^(a[187] & b[147])^(a[186] & b[148])^(a[185] & b[149])^(a[184] & b[150])^(a[183] & b[151])^(a[182] & b[152])^(a[181] & b[153])^(a[180] & b[154])^(a[179] & b[155])^(a[178] & b[156])^(a[177] & b[157])^(a[176] & b[158])^(a[175] & b[159])^(a[174] & b[160])^(a[173] & b[161])^(a[172] & b[162])^(a[171] & b[163])^(a[170] & b[164])^(a[169] & b[165])^(a[168] & b[166])^(a[167] & b[167])^(a[166] & b[168])^(a[165] & b[169])^(a[164] & b[170])^(a[163] & b[171])^(a[162] & b[172])^(a[161] & b[173])^(a[160] & b[174])^(a[159] & b[175])^(a[158] & b[176])^(a[157] & b[177])^(a[156] & b[178])^(a[155] & b[179])^(a[154] & b[180])^(a[153] & b[181])^(a[152] & b[182])^(a[151] & b[183])^(a[150] & b[184])^(a[149] & b[185])^(a[148] & b[186])^(a[147] & b[187])^(a[146] & b[188])^(a[145] & b[189])^(a[144] & b[190])^(a[143] & b[191])^(a[142] & b[192])^(a[141] & b[193])^(a[140] & b[194])^(a[139] & b[195])^(a[138] & b[196])^(a[137] & b[197])^(a[136] & b[198])^(a[135] & b[199])^(a[134] & b[200])^(a[133] & b[201])^(a[132] & b[202])^(a[131] & b[203])^(a[130] & b[204])^(a[129] & b[205])^(a[128] & b[206])^(a[127] & b[207])^(a[126] & b[208])^(a[125] & b[209])^(a[124] & b[210])^(a[123] & b[211])^(a[122] & b[212])^(a[121] & b[213])^(a[120] & b[214])^(a[119] & b[215])^(a[118] & b[216])^(a[117] & b[217])^(a[116] & b[218])^(a[115] & b[219])^(a[114] & b[220])^(a[113] & b[221])^(a[112] & b[222])^(a[111] & b[223])^(a[110] & b[224])^(a[109] & b[225])^(a[108] & b[226])^(a[107] & b[227])^(a[106] & b[228])^(a[105] & b[229])^(a[104] & b[230])^(a[103] & b[231])^(a[102] & b[232])^(a[101] & b[233])^(a[100] & b[234])^(a[99] & b[235])^(a[98] & b[236])^(a[97] & b[237])^(a[96] & b[238])^(a[95] & b[239])^(a[94] & b[240])^(a[93] & b[241])^(a[92] & b[242])^(a[91] & b[243])^(a[90] & b[244])^(a[89] & b[245])^(a[88] & b[246])^(a[87] & b[247])^(a[86] & b[248])^(a[85] & b[249])^(a[84] & b[250])^(a[83] & b[251])^(a[82] & b[252])^(a[81] & b[253])^(a[80] & b[254])^(a[79] & b[255])^(a[78] & b[256])^(a[77] & b[257])^(a[76] & b[258])^(a[75] & b[259])^(a[74] & b[260])^(a[73] & b[261])^(a[72] & b[262])^(a[71] & b[263])^(a[70] & b[264])^(a[69] & b[265])^(a[68] & b[266])^(a[67] & b[267])^(a[66] & b[268])^(a[65] & b[269])^(a[64] & b[270])^(a[63] & b[271])^(a[62] & b[272])^(a[61] & b[273])^(a[60] & b[274])^(a[59] & b[275])^(a[58] & b[276])^(a[57] & b[277])^(a[56] & b[278])^(a[55] & b[279])^(a[54] & b[280])^(a[53] & b[281])^(a[52] & b[282])^(a[51] & b[283])^(a[50] & b[284])^(a[49] & b[285])^(a[48] & b[286])^(a[47] & b[287])^(a[46] & b[288])^(a[45] & b[289])^(a[44] & b[290])^(a[43] & b[291])^(a[42] & b[292])^(a[41] & b[293])^(a[40] & b[294])^(a[39] & b[295])^(a[38] & b[296])^(a[37] & b[297])^(a[36] & b[298])^(a[35] & b[299])^(a[34] & b[300])^(a[33] & b[301])^(a[32] & b[302])^(a[31] & b[303])^(a[30] & b[304])^(a[29] & b[305])^(a[28] & b[306])^(a[27] & b[307])^(a[26] & b[308])^(a[25] & b[309])^(a[24] & b[310])^(a[23] & b[311])^(a[22] & b[312])^(a[21] & b[313])^(a[20] & b[314])^(a[19] & b[315])^(a[18] & b[316])^(a[17] & b[317])^(a[16] & b[318])^(a[15] & b[319])^(a[14] & b[320])^(a[13] & b[321])^(a[12] & b[322])^(a[11] & b[323])^(a[10] & b[324])^(a[9] & b[325])^(a[8] & b[326])^(a[7] & b[327])^(a[6] & b[328])^(a[5] & b[329])^(a[4] & b[330])^(a[3] & b[331])^(a[2] & b[332])^(a[1] & b[333])^(a[0] & b[334]);
assign y[335] = (a[335] & b[0])^(a[334] & b[1])^(a[333] & b[2])^(a[332] & b[3])^(a[331] & b[4])^(a[330] & b[5])^(a[329] & b[6])^(a[328] & b[7])^(a[327] & b[8])^(a[326] & b[9])^(a[325] & b[10])^(a[324] & b[11])^(a[323] & b[12])^(a[322] & b[13])^(a[321] & b[14])^(a[320] & b[15])^(a[319] & b[16])^(a[318] & b[17])^(a[317] & b[18])^(a[316] & b[19])^(a[315] & b[20])^(a[314] & b[21])^(a[313] & b[22])^(a[312] & b[23])^(a[311] & b[24])^(a[310] & b[25])^(a[309] & b[26])^(a[308] & b[27])^(a[307] & b[28])^(a[306] & b[29])^(a[305] & b[30])^(a[304] & b[31])^(a[303] & b[32])^(a[302] & b[33])^(a[301] & b[34])^(a[300] & b[35])^(a[299] & b[36])^(a[298] & b[37])^(a[297] & b[38])^(a[296] & b[39])^(a[295] & b[40])^(a[294] & b[41])^(a[293] & b[42])^(a[292] & b[43])^(a[291] & b[44])^(a[290] & b[45])^(a[289] & b[46])^(a[288] & b[47])^(a[287] & b[48])^(a[286] & b[49])^(a[285] & b[50])^(a[284] & b[51])^(a[283] & b[52])^(a[282] & b[53])^(a[281] & b[54])^(a[280] & b[55])^(a[279] & b[56])^(a[278] & b[57])^(a[277] & b[58])^(a[276] & b[59])^(a[275] & b[60])^(a[274] & b[61])^(a[273] & b[62])^(a[272] & b[63])^(a[271] & b[64])^(a[270] & b[65])^(a[269] & b[66])^(a[268] & b[67])^(a[267] & b[68])^(a[266] & b[69])^(a[265] & b[70])^(a[264] & b[71])^(a[263] & b[72])^(a[262] & b[73])^(a[261] & b[74])^(a[260] & b[75])^(a[259] & b[76])^(a[258] & b[77])^(a[257] & b[78])^(a[256] & b[79])^(a[255] & b[80])^(a[254] & b[81])^(a[253] & b[82])^(a[252] & b[83])^(a[251] & b[84])^(a[250] & b[85])^(a[249] & b[86])^(a[248] & b[87])^(a[247] & b[88])^(a[246] & b[89])^(a[245] & b[90])^(a[244] & b[91])^(a[243] & b[92])^(a[242] & b[93])^(a[241] & b[94])^(a[240] & b[95])^(a[239] & b[96])^(a[238] & b[97])^(a[237] & b[98])^(a[236] & b[99])^(a[235] & b[100])^(a[234] & b[101])^(a[233] & b[102])^(a[232] & b[103])^(a[231] & b[104])^(a[230] & b[105])^(a[229] & b[106])^(a[228] & b[107])^(a[227] & b[108])^(a[226] & b[109])^(a[225] & b[110])^(a[224] & b[111])^(a[223] & b[112])^(a[222] & b[113])^(a[221] & b[114])^(a[220] & b[115])^(a[219] & b[116])^(a[218] & b[117])^(a[217] & b[118])^(a[216] & b[119])^(a[215] & b[120])^(a[214] & b[121])^(a[213] & b[122])^(a[212] & b[123])^(a[211] & b[124])^(a[210] & b[125])^(a[209] & b[126])^(a[208] & b[127])^(a[207] & b[128])^(a[206] & b[129])^(a[205] & b[130])^(a[204] & b[131])^(a[203] & b[132])^(a[202] & b[133])^(a[201] & b[134])^(a[200] & b[135])^(a[199] & b[136])^(a[198] & b[137])^(a[197] & b[138])^(a[196] & b[139])^(a[195] & b[140])^(a[194] & b[141])^(a[193] & b[142])^(a[192] & b[143])^(a[191] & b[144])^(a[190] & b[145])^(a[189] & b[146])^(a[188] & b[147])^(a[187] & b[148])^(a[186] & b[149])^(a[185] & b[150])^(a[184] & b[151])^(a[183] & b[152])^(a[182] & b[153])^(a[181] & b[154])^(a[180] & b[155])^(a[179] & b[156])^(a[178] & b[157])^(a[177] & b[158])^(a[176] & b[159])^(a[175] & b[160])^(a[174] & b[161])^(a[173] & b[162])^(a[172] & b[163])^(a[171] & b[164])^(a[170] & b[165])^(a[169] & b[166])^(a[168] & b[167])^(a[167] & b[168])^(a[166] & b[169])^(a[165] & b[170])^(a[164] & b[171])^(a[163] & b[172])^(a[162] & b[173])^(a[161] & b[174])^(a[160] & b[175])^(a[159] & b[176])^(a[158] & b[177])^(a[157] & b[178])^(a[156] & b[179])^(a[155] & b[180])^(a[154] & b[181])^(a[153] & b[182])^(a[152] & b[183])^(a[151] & b[184])^(a[150] & b[185])^(a[149] & b[186])^(a[148] & b[187])^(a[147] & b[188])^(a[146] & b[189])^(a[145] & b[190])^(a[144] & b[191])^(a[143] & b[192])^(a[142] & b[193])^(a[141] & b[194])^(a[140] & b[195])^(a[139] & b[196])^(a[138] & b[197])^(a[137] & b[198])^(a[136] & b[199])^(a[135] & b[200])^(a[134] & b[201])^(a[133] & b[202])^(a[132] & b[203])^(a[131] & b[204])^(a[130] & b[205])^(a[129] & b[206])^(a[128] & b[207])^(a[127] & b[208])^(a[126] & b[209])^(a[125] & b[210])^(a[124] & b[211])^(a[123] & b[212])^(a[122] & b[213])^(a[121] & b[214])^(a[120] & b[215])^(a[119] & b[216])^(a[118] & b[217])^(a[117] & b[218])^(a[116] & b[219])^(a[115] & b[220])^(a[114] & b[221])^(a[113] & b[222])^(a[112] & b[223])^(a[111] & b[224])^(a[110] & b[225])^(a[109] & b[226])^(a[108] & b[227])^(a[107] & b[228])^(a[106] & b[229])^(a[105] & b[230])^(a[104] & b[231])^(a[103] & b[232])^(a[102] & b[233])^(a[101] & b[234])^(a[100] & b[235])^(a[99] & b[236])^(a[98] & b[237])^(a[97] & b[238])^(a[96] & b[239])^(a[95] & b[240])^(a[94] & b[241])^(a[93] & b[242])^(a[92] & b[243])^(a[91] & b[244])^(a[90] & b[245])^(a[89] & b[246])^(a[88] & b[247])^(a[87] & b[248])^(a[86] & b[249])^(a[85] & b[250])^(a[84] & b[251])^(a[83] & b[252])^(a[82] & b[253])^(a[81] & b[254])^(a[80] & b[255])^(a[79] & b[256])^(a[78] & b[257])^(a[77] & b[258])^(a[76] & b[259])^(a[75] & b[260])^(a[74] & b[261])^(a[73] & b[262])^(a[72] & b[263])^(a[71] & b[264])^(a[70] & b[265])^(a[69] & b[266])^(a[68] & b[267])^(a[67] & b[268])^(a[66] & b[269])^(a[65] & b[270])^(a[64] & b[271])^(a[63] & b[272])^(a[62] & b[273])^(a[61] & b[274])^(a[60] & b[275])^(a[59] & b[276])^(a[58] & b[277])^(a[57] & b[278])^(a[56] & b[279])^(a[55] & b[280])^(a[54] & b[281])^(a[53] & b[282])^(a[52] & b[283])^(a[51] & b[284])^(a[50] & b[285])^(a[49] & b[286])^(a[48] & b[287])^(a[47] & b[288])^(a[46] & b[289])^(a[45] & b[290])^(a[44] & b[291])^(a[43] & b[292])^(a[42] & b[293])^(a[41] & b[294])^(a[40] & b[295])^(a[39] & b[296])^(a[38] & b[297])^(a[37] & b[298])^(a[36] & b[299])^(a[35] & b[300])^(a[34] & b[301])^(a[33] & b[302])^(a[32] & b[303])^(a[31] & b[304])^(a[30] & b[305])^(a[29] & b[306])^(a[28] & b[307])^(a[27] & b[308])^(a[26] & b[309])^(a[25] & b[310])^(a[24] & b[311])^(a[23] & b[312])^(a[22] & b[313])^(a[21] & b[314])^(a[20] & b[315])^(a[19] & b[316])^(a[18] & b[317])^(a[17] & b[318])^(a[16] & b[319])^(a[15] & b[320])^(a[14] & b[321])^(a[13] & b[322])^(a[12] & b[323])^(a[11] & b[324])^(a[10] & b[325])^(a[9] & b[326])^(a[8] & b[327])^(a[7] & b[328])^(a[6] & b[329])^(a[5] & b[330])^(a[4] & b[331])^(a[3] & b[332])^(a[2] & b[333])^(a[1] & b[334])^(a[0] & b[335]);
assign y[336] = (a[336] & b[0])^(a[335] & b[1])^(a[334] & b[2])^(a[333] & b[3])^(a[332] & b[4])^(a[331] & b[5])^(a[330] & b[6])^(a[329] & b[7])^(a[328] & b[8])^(a[327] & b[9])^(a[326] & b[10])^(a[325] & b[11])^(a[324] & b[12])^(a[323] & b[13])^(a[322] & b[14])^(a[321] & b[15])^(a[320] & b[16])^(a[319] & b[17])^(a[318] & b[18])^(a[317] & b[19])^(a[316] & b[20])^(a[315] & b[21])^(a[314] & b[22])^(a[313] & b[23])^(a[312] & b[24])^(a[311] & b[25])^(a[310] & b[26])^(a[309] & b[27])^(a[308] & b[28])^(a[307] & b[29])^(a[306] & b[30])^(a[305] & b[31])^(a[304] & b[32])^(a[303] & b[33])^(a[302] & b[34])^(a[301] & b[35])^(a[300] & b[36])^(a[299] & b[37])^(a[298] & b[38])^(a[297] & b[39])^(a[296] & b[40])^(a[295] & b[41])^(a[294] & b[42])^(a[293] & b[43])^(a[292] & b[44])^(a[291] & b[45])^(a[290] & b[46])^(a[289] & b[47])^(a[288] & b[48])^(a[287] & b[49])^(a[286] & b[50])^(a[285] & b[51])^(a[284] & b[52])^(a[283] & b[53])^(a[282] & b[54])^(a[281] & b[55])^(a[280] & b[56])^(a[279] & b[57])^(a[278] & b[58])^(a[277] & b[59])^(a[276] & b[60])^(a[275] & b[61])^(a[274] & b[62])^(a[273] & b[63])^(a[272] & b[64])^(a[271] & b[65])^(a[270] & b[66])^(a[269] & b[67])^(a[268] & b[68])^(a[267] & b[69])^(a[266] & b[70])^(a[265] & b[71])^(a[264] & b[72])^(a[263] & b[73])^(a[262] & b[74])^(a[261] & b[75])^(a[260] & b[76])^(a[259] & b[77])^(a[258] & b[78])^(a[257] & b[79])^(a[256] & b[80])^(a[255] & b[81])^(a[254] & b[82])^(a[253] & b[83])^(a[252] & b[84])^(a[251] & b[85])^(a[250] & b[86])^(a[249] & b[87])^(a[248] & b[88])^(a[247] & b[89])^(a[246] & b[90])^(a[245] & b[91])^(a[244] & b[92])^(a[243] & b[93])^(a[242] & b[94])^(a[241] & b[95])^(a[240] & b[96])^(a[239] & b[97])^(a[238] & b[98])^(a[237] & b[99])^(a[236] & b[100])^(a[235] & b[101])^(a[234] & b[102])^(a[233] & b[103])^(a[232] & b[104])^(a[231] & b[105])^(a[230] & b[106])^(a[229] & b[107])^(a[228] & b[108])^(a[227] & b[109])^(a[226] & b[110])^(a[225] & b[111])^(a[224] & b[112])^(a[223] & b[113])^(a[222] & b[114])^(a[221] & b[115])^(a[220] & b[116])^(a[219] & b[117])^(a[218] & b[118])^(a[217] & b[119])^(a[216] & b[120])^(a[215] & b[121])^(a[214] & b[122])^(a[213] & b[123])^(a[212] & b[124])^(a[211] & b[125])^(a[210] & b[126])^(a[209] & b[127])^(a[208] & b[128])^(a[207] & b[129])^(a[206] & b[130])^(a[205] & b[131])^(a[204] & b[132])^(a[203] & b[133])^(a[202] & b[134])^(a[201] & b[135])^(a[200] & b[136])^(a[199] & b[137])^(a[198] & b[138])^(a[197] & b[139])^(a[196] & b[140])^(a[195] & b[141])^(a[194] & b[142])^(a[193] & b[143])^(a[192] & b[144])^(a[191] & b[145])^(a[190] & b[146])^(a[189] & b[147])^(a[188] & b[148])^(a[187] & b[149])^(a[186] & b[150])^(a[185] & b[151])^(a[184] & b[152])^(a[183] & b[153])^(a[182] & b[154])^(a[181] & b[155])^(a[180] & b[156])^(a[179] & b[157])^(a[178] & b[158])^(a[177] & b[159])^(a[176] & b[160])^(a[175] & b[161])^(a[174] & b[162])^(a[173] & b[163])^(a[172] & b[164])^(a[171] & b[165])^(a[170] & b[166])^(a[169] & b[167])^(a[168] & b[168])^(a[167] & b[169])^(a[166] & b[170])^(a[165] & b[171])^(a[164] & b[172])^(a[163] & b[173])^(a[162] & b[174])^(a[161] & b[175])^(a[160] & b[176])^(a[159] & b[177])^(a[158] & b[178])^(a[157] & b[179])^(a[156] & b[180])^(a[155] & b[181])^(a[154] & b[182])^(a[153] & b[183])^(a[152] & b[184])^(a[151] & b[185])^(a[150] & b[186])^(a[149] & b[187])^(a[148] & b[188])^(a[147] & b[189])^(a[146] & b[190])^(a[145] & b[191])^(a[144] & b[192])^(a[143] & b[193])^(a[142] & b[194])^(a[141] & b[195])^(a[140] & b[196])^(a[139] & b[197])^(a[138] & b[198])^(a[137] & b[199])^(a[136] & b[200])^(a[135] & b[201])^(a[134] & b[202])^(a[133] & b[203])^(a[132] & b[204])^(a[131] & b[205])^(a[130] & b[206])^(a[129] & b[207])^(a[128] & b[208])^(a[127] & b[209])^(a[126] & b[210])^(a[125] & b[211])^(a[124] & b[212])^(a[123] & b[213])^(a[122] & b[214])^(a[121] & b[215])^(a[120] & b[216])^(a[119] & b[217])^(a[118] & b[218])^(a[117] & b[219])^(a[116] & b[220])^(a[115] & b[221])^(a[114] & b[222])^(a[113] & b[223])^(a[112] & b[224])^(a[111] & b[225])^(a[110] & b[226])^(a[109] & b[227])^(a[108] & b[228])^(a[107] & b[229])^(a[106] & b[230])^(a[105] & b[231])^(a[104] & b[232])^(a[103] & b[233])^(a[102] & b[234])^(a[101] & b[235])^(a[100] & b[236])^(a[99] & b[237])^(a[98] & b[238])^(a[97] & b[239])^(a[96] & b[240])^(a[95] & b[241])^(a[94] & b[242])^(a[93] & b[243])^(a[92] & b[244])^(a[91] & b[245])^(a[90] & b[246])^(a[89] & b[247])^(a[88] & b[248])^(a[87] & b[249])^(a[86] & b[250])^(a[85] & b[251])^(a[84] & b[252])^(a[83] & b[253])^(a[82] & b[254])^(a[81] & b[255])^(a[80] & b[256])^(a[79] & b[257])^(a[78] & b[258])^(a[77] & b[259])^(a[76] & b[260])^(a[75] & b[261])^(a[74] & b[262])^(a[73] & b[263])^(a[72] & b[264])^(a[71] & b[265])^(a[70] & b[266])^(a[69] & b[267])^(a[68] & b[268])^(a[67] & b[269])^(a[66] & b[270])^(a[65] & b[271])^(a[64] & b[272])^(a[63] & b[273])^(a[62] & b[274])^(a[61] & b[275])^(a[60] & b[276])^(a[59] & b[277])^(a[58] & b[278])^(a[57] & b[279])^(a[56] & b[280])^(a[55] & b[281])^(a[54] & b[282])^(a[53] & b[283])^(a[52] & b[284])^(a[51] & b[285])^(a[50] & b[286])^(a[49] & b[287])^(a[48] & b[288])^(a[47] & b[289])^(a[46] & b[290])^(a[45] & b[291])^(a[44] & b[292])^(a[43] & b[293])^(a[42] & b[294])^(a[41] & b[295])^(a[40] & b[296])^(a[39] & b[297])^(a[38] & b[298])^(a[37] & b[299])^(a[36] & b[300])^(a[35] & b[301])^(a[34] & b[302])^(a[33] & b[303])^(a[32] & b[304])^(a[31] & b[305])^(a[30] & b[306])^(a[29] & b[307])^(a[28] & b[308])^(a[27] & b[309])^(a[26] & b[310])^(a[25] & b[311])^(a[24] & b[312])^(a[23] & b[313])^(a[22] & b[314])^(a[21] & b[315])^(a[20] & b[316])^(a[19] & b[317])^(a[18] & b[318])^(a[17] & b[319])^(a[16] & b[320])^(a[15] & b[321])^(a[14] & b[322])^(a[13] & b[323])^(a[12] & b[324])^(a[11] & b[325])^(a[10] & b[326])^(a[9] & b[327])^(a[8] & b[328])^(a[7] & b[329])^(a[6] & b[330])^(a[5] & b[331])^(a[4] & b[332])^(a[3] & b[333])^(a[2] & b[334])^(a[1] & b[335])^(a[0] & b[336]);
assign y[337] = (a[337] & b[0])^(a[336] & b[1])^(a[335] & b[2])^(a[334] & b[3])^(a[333] & b[4])^(a[332] & b[5])^(a[331] & b[6])^(a[330] & b[7])^(a[329] & b[8])^(a[328] & b[9])^(a[327] & b[10])^(a[326] & b[11])^(a[325] & b[12])^(a[324] & b[13])^(a[323] & b[14])^(a[322] & b[15])^(a[321] & b[16])^(a[320] & b[17])^(a[319] & b[18])^(a[318] & b[19])^(a[317] & b[20])^(a[316] & b[21])^(a[315] & b[22])^(a[314] & b[23])^(a[313] & b[24])^(a[312] & b[25])^(a[311] & b[26])^(a[310] & b[27])^(a[309] & b[28])^(a[308] & b[29])^(a[307] & b[30])^(a[306] & b[31])^(a[305] & b[32])^(a[304] & b[33])^(a[303] & b[34])^(a[302] & b[35])^(a[301] & b[36])^(a[300] & b[37])^(a[299] & b[38])^(a[298] & b[39])^(a[297] & b[40])^(a[296] & b[41])^(a[295] & b[42])^(a[294] & b[43])^(a[293] & b[44])^(a[292] & b[45])^(a[291] & b[46])^(a[290] & b[47])^(a[289] & b[48])^(a[288] & b[49])^(a[287] & b[50])^(a[286] & b[51])^(a[285] & b[52])^(a[284] & b[53])^(a[283] & b[54])^(a[282] & b[55])^(a[281] & b[56])^(a[280] & b[57])^(a[279] & b[58])^(a[278] & b[59])^(a[277] & b[60])^(a[276] & b[61])^(a[275] & b[62])^(a[274] & b[63])^(a[273] & b[64])^(a[272] & b[65])^(a[271] & b[66])^(a[270] & b[67])^(a[269] & b[68])^(a[268] & b[69])^(a[267] & b[70])^(a[266] & b[71])^(a[265] & b[72])^(a[264] & b[73])^(a[263] & b[74])^(a[262] & b[75])^(a[261] & b[76])^(a[260] & b[77])^(a[259] & b[78])^(a[258] & b[79])^(a[257] & b[80])^(a[256] & b[81])^(a[255] & b[82])^(a[254] & b[83])^(a[253] & b[84])^(a[252] & b[85])^(a[251] & b[86])^(a[250] & b[87])^(a[249] & b[88])^(a[248] & b[89])^(a[247] & b[90])^(a[246] & b[91])^(a[245] & b[92])^(a[244] & b[93])^(a[243] & b[94])^(a[242] & b[95])^(a[241] & b[96])^(a[240] & b[97])^(a[239] & b[98])^(a[238] & b[99])^(a[237] & b[100])^(a[236] & b[101])^(a[235] & b[102])^(a[234] & b[103])^(a[233] & b[104])^(a[232] & b[105])^(a[231] & b[106])^(a[230] & b[107])^(a[229] & b[108])^(a[228] & b[109])^(a[227] & b[110])^(a[226] & b[111])^(a[225] & b[112])^(a[224] & b[113])^(a[223] & b[114])^(a[222] & b[115])^(a[221] & b[116])^(a[220] & b[117])^(a[219] & b[118])^(a[218] & b[119])^(a[217] & b[120])^(a[216] & b[121])^(a[215] & b[122])^(a[214] & b[123])^(a[213] & b[124])^(a[212] & b[125])^(a[211] & b[126])^(a[210] & b[127])^(a[209] & b[128])^(a[208] & b[129])^(a[207] & b[130])^(a[206] & b[131])^(a[205] & b[132])^(a[204] & b[133])^(a[203] & b[134])^(a[202] & b[135])^(a[201] & b[136])^(a[200] & b[137])^(a[199] & b[138])^(a[198] & b[139])^(a[197] & b[140])^(a[196] & b[141])^(a[195] & b[142])^(a[194] & b[143])^(a[193] & b[144])^(a[192] & b[145])^(a[191] & b[146])^(a[190] & b[147])^(a[189] & b[148])^(a[188] & b[149])^(a[187] & b[150])^(a[186] & b[151])^(a[185] & b[152])^(a[184] & b[153])^(a[183] & b[154])^(a[182] & b[155])^(a[181] & b[156])^(a[180] & b[157])^(a[179] & b[158])^(a[178] & b[159])^(a[177] & b[160])^(a[176] & b[161])^(a[175] & b[162])^(a[174] & b[163])^(a[173] & b[164])^(a[172] & b[165])^(a[171] & b[166])^(a[170] & b[167])^(a[169] & b[168])^(a[168] & b[169])^(a[167] & b[170])^(a[166] & b[171])^(a[165] & b[172])^(a[164] & b[173])^(a[163] & b[174])^(a[162] & b[175])^(a[161] & b[176])^(a[160] & b[177])^(a[159] & b[178])^(a[158] & b[179])^(a[157] & b[180])^(a[156] & b[181])^(a[155] & b[182])^(a[154] & b[183])^(a[153] & b[184])^(a[152] & b[185])^(a[151] & b[186])^(a[150] & b[187])^(a[149] & b[188])^(a[148] & b[189])^(a[147] & b[190])^(a[146] & b[191])^(a[145] & b[192])^(a[144] & b[193])^(a[143] & b[194])^(a[142] & b[195])^(a[141] & b[196])^(a[140] & b[197])^(a[139] & b[198])^(a[138] & b[199])^(a[137] & b[200])^(a[136] & b[201])^(a[135] & b[202])^(a[134] & b[203])^(a[133] & b[204])^(a[132] & b[205])^(a[131] & b[206])^(a[130] & b[207])^(a[129] & b[208])^(a[128] & b[209])^(a[127] & b[210])^(a[126] & b[211])^(a[125] & b[212])^(a[124] & b[213])^(a[123] & b[214])^(a[122] & b[215])^(a[121] & b[216])^(a[120] & b[217])^(a[119] & b[218])^(a[118] & b[219])^(a[117] & b[220])^(a[116] & b[221])^(a[115] & b[222])^(a[114] & b[223])^(a[113] & b[224])^(a[112] & b[225])^(a[111] & b[226])^(a[110] & b[227])^(a[109] & b[228])^(a[108] & b[229])^(a[107] & b[230])^(a[106] & b[231])^(a[105] & b[232])^(a[104] & b[233])^(a[103] & b[234])^(a[102] & b[235])^(a[101] & b[236])^(a[100] & b[237])^(a[99] & b[238])^(a[98] & b[239])^(a[97] & b[240])^(a[96] & b[241])^(a[95] & b[242])^(a[94] & b[243])^(a[93] & b[244])^(a[92] & b[245])^(a[91] & b[246])^(a[90] & b[247])^(a[89] & b[248])^(a[88] & b[249])^(a[87] & b[250])^(a[86] & b[251])^(a[85] & b[252])^(a[84] & b[253])^(a[83] & b[254])^(a[82] & b[255])^(a[81] & b[256])^(a[80] & b[257])^(a[79] & b[258])^(a[78] & b[259])^(a[77] & b[260])^(a[76] & b[261])^(a[75] & b[262])^(a[74] & b[263])^(a[73] & b[264])^(a[72] & b[265])^(a[71] & b[266])^(a[70] & b[267])^(a[69] & b[268])^(a[68] & b[269])^(a[67] & b[270])^(a[66] & b[271])^(a[65] & b[272])^(a[64] & b[273])^(a[63] & b[274])^(a[62] & b[275])^(a[61] & b[276])^(a[60] & b[277])^(a[59] & b[278])^(a[58] & b[279])^(a[57] & b[280])^(a[56] & b[281])^(a[55] & b[282])^(a[54] & b[283])^(a[53] & b[284])^(a[52] & b[285])^(a[51] & b[286])^(a[50] & b[287])^(a[49] & b[288])^(a[48] & b[289])^(a[47] & b[290])^(a[46] & b[291])^(a[45] & b[292])^(a[44] & b[293])^(a[43] & b[294])^(a[42] & b[295])^(a[41] & b[296])^(a[40] & b[297])^(a[39] & b[298])^(a[38] & b[299])^(a[37] & b[300])^(a[36] & b[301])^(a[35] & b[302])^(a[34] & b[303])^(a[33] & b[304])^(a[32] & b[305])^(a[31] & b[306])^(a[30] & b[307])^(a[29] & b[308])^(a[28] & b[309])^(a[27] & b[310])^(a[26] & b[311])^(a[25] & b[312])^(a[24] & b[313])^(a[23] & b[314])^(a[22] & b[315])^(a[21] & b[316])^(a[20] & b[317])^(a[19] & b[318])^(a[18] & b[319])^(a[17] & b[320])^(a[16] & b[321])^(a[15] & b[322])^(a[14] & b[323])^(a[13] & b[324])^(a[12] & b[325])^(a[11] & b[326])^(a[10] & b[327])^(a[9] & b[328])^(a[8] & b[329])^(a[7] & b[330])^(a[6] & b[331])^(a[5] & b[332])^(a[4] & b[333])^(a[3] & b[334])^(a[2] & b[335])^(a[1] & b[336])^(a[0] & b[337]);
assign y[338] = (a[338] & b[0])^(a[337] & b[1])^(a[336] & b[2])^(a[335] & b[3])^(a[334] & b[4])^(a[333] & b[5])^(a[332] & b[6])^(a[331] & b[7])^(a[330] & b[8])^(a[329] & b[9])^(a[328] & b[10])^(a[327] & b[11])^(a[326] & b[12])^(a[325] & b[13])^(a[324] & b[14])^(a[323] & b[15])^(a[322] & b[16])^(a[321] & b[17])^(a[320] & b[18])^(a[319] & b[19])^(a[318] & b[20])^(a[317] & b[21])^(a[316] & b[22])^(a[315] & b[23])^(a[314] & b[24])^(a[313] & b[25])^(a[312] & b[26])^(a[311] & b[27])^(a[310] & b[28])^(a[309] & b[29])^(a[308] & b[30])^(a[307] & b[31])^(a[306] & b[32])^(a[305] & b[33])^(a[304] & b[34])^(a[303] & b[35])^(a[302] & b[36])^(a[301] & b[37])^(a[300] & b[38])^(a[299] & b[39])^(a[298] & b[40])^(a[297] & b[41])^(a[296] & b[42])^(a[295] & b[43])^(a[294] & b[44])^(a[293] & b[45])^(a[292] & b[46])^(a[291] & b[47])^(a[290] & b[48])^(a[289] & b[49])^(a[288] & b[50])^(a[287] & b[51])^(a[286] & b[52])^(a[285] & b[53])^(a[284] & b[54])^(a[283] & b[55])^(a[282] & b[56])^(a[281] & b[57])^(a[280] & b[58])^(a[279] & b[59])^(a[278] & b[60])^(a[277] & b[61])^(a[276] & b[62])^(a[275] & b[63])^(a[274] & b[64])^(a[273] & b[65])^(a[272] & b[66])^(a[271] & b[67])^(a[270] & b[68])^(a[269] & b[69])^(a[268] & b[70])^(a[267] & b[71])^(a[266] & b[72])^(a[265] & b[73])^(a[264] & b[74])^(a[263] & b[75])^(a[262] & b[76])^(a[261] & b[77])^(a[260] & b[78])^(a[259] & b[79])^(a[258] & b[80])^(a[257] & b[81])^(a[256] & b[82])^(a[255] & b[83])^(a[254] & b[84])^(a[253] & b[85])^(a[252] & b[86])^(a[251] & b[87])^(a[250] & b[88])^(a[249] & b[89])^(a[248] & b[90])^(a[247] & b[91])^(a[246] & b[92])^(a[245] & b[93])^(a[244] & b[94])^(a[243] & b[95])^(a[242] & b[96])^(a[241] & b[97])^(a[240] & b[98])^(a[239] & b[99])^(a[238] & b[100])^(a[237] & b[101])^(a[236] & b[102])^(a[235] & b[103])^(a[234] & b[104])^(a[233] & b[105])^(a[232] & b[106])^(a[231] & b[107])^(a[230] & b[108])^(a[229] & b[109])^(a[228] & b[110])^(a[227] & b[111])^(a[226] & b[112])^(a[225] & b[113])^(a[224] & b[114])^(a[223] & b[115])^(a[222] & b[116])^(a[221] & b[117])^(a[220] & b[118])^(a[219] & b[119])^(a[218] & b[120])^(a[217] & b[121])^(a[216] & b[122])^(a[215] & b[123])^(a[214] & b[124])^(a[213] & b[125])^(a[212] & b[126])^(a[211] & b[127])^(a[210] & b[128])^(a[209] & b[129])^(a[208] & b[130])^(a[207] & b[131])^(a[206] & b[132])^(a[205] & b[133])^(a[204] & b[134])^(a[203] & b[135])^(a[202] & b[136])^(a[201] & b[137])^(a[200] & b[138])^(a[199] & b[139])^(a[198] & b[140])^(a[197] & b[141])^(a[196] & b[142])^(a[195] & b[143])^(a[194] & b[144])^(a[193] & b[145])^(a[192] & b[146])^(a[191] & b[147])^(a[190] & b[148])^(a[189] & b[149])^(a[188] & b[150])^(a[187] & b[151])^(a[186] & b[152])^(a[185] & b[153])^(a[184] & b[154])^(a[183] & b[155])^(a[182] & b[156])^(a[181] & b[157])^(a[180] & b[158])^(a[179] & b[159])^(a[178] & b[160])^(a[177] & b[161])^(a[176] & b[162])^(a[175] & b[163])^(a[174] & b[164])^(a[173] & b[165])^(a[172] & b[166])^(a[171] & b[167])^(a[170] & b[168])^(a[169] & b[169])^(a[168] & b[170])^(a[167] & b[171])^(a[166] & b[172])^(a[165] & b[173])^(a[164] & b[174])^(a[163] & b[175])^(a[162] & b[176])^(a[161] & b[177])^(a[160] & b[178])^(a[159] & b[179])^(a[158] & b[180])^(a[157] & b[181])^(a[156] & b[182])^(a[155] & b[183])^(a[154] & b[184])^(a[153] & b[185])^(a[152] & b[186])^(a[151] & b[187])^(a[150] & b[188])^(a[149] & b[189])^(a[148] & b[190])^(a[147] & b[191])^(a[146] & b[192])^(a[145] & b[193])^(a[144] & b[194])^(a[143] & b[195])^(a[142] & b[196])^(a[141] & b[197])^(a[140] & b[198])^(a[139] & b[199])^(a[138] & b[200])^(a[137] & b[201])^(a[136] & b[202])^(a[135] & b[203])^(a[134] & b[204])^(a[133] & b[205])^(a[132] & b[206])^(a[131] & b[207])^(a[130] & b[208])^(a[129] & b[209])^(a[128] & b[210])^(a[127] & b[211])^(a[126] & b[212])^(a[125] & b[213])^(a[124] & b[214])^(a[123] & b[215])^(a[122] & b[216])^(a[121] & b[217])^(a[120] & b[218])^(a[119] & b[219])^(a[118] & b[220])^(a[117] & b[221])^(a[116] & b[222])^(a[115] & b[223])^(a[114] & b[224])^(a[113] & b[225])^(a[112] & b[226])^(a[111] & b[227])^(a[110] & b[228])^(a[109] & b[229])^(a[108] & b[230])^(a[107] & b[231])^(a[106] & b[232])^(a[105] & b[233])^(a[104] & b[234])^(a[103] & b[235])^(a[102] & b[236])^(a[101] & b[237])^(a[100] & b[238])^(a[99] & b[239])^(a[98] & b[240])^(a[97] & b[241])^(a[96] & b[242])^(a[95] & b[243])^(a[94] & b[244])^(a[93] & b[245])^(a[92] & b[246])^(a[91] & b[247])^(a[90] & b[248])^(a[89] & b[249])^(a[88] & b[250])^(a[87] & b[251])^(a[86] & b[252])^(a[85] & b[253])^(a[84] & b[254])^(a[83] & b[255])^(a[82] & b[256])^(a[81] & b[257])^(a[80] & b[258])^(a[79] & b[259])^(a[78] & b[260])^(a[77] & b[261])^(a[76] & b[262])^(a[75] & b[263])^(a[74] & b[264])^(a[73] & b[265])^(a[72] & b[266])^(a[71] & b[267])^(a[70] & b[268])^(a[69] & b[269])^(a[68] & b[270])^(a[67] & b[271])^(a[66] & b[272])^(a[65] & b[273])^(a[64] & b[274])^(a[63] & b[275])^(a[62] & b[276])^(a[61] & b[277])^(a[60] & b[278])^(a[59] & b[279])^(a[58] & b[280])^(a[57] & b[281])^(a[56] & b[282])^(a[55] & b[283])^(a[54] & b[284])^(a[53] & b[285])^(a[52] & b[286])^(a[51] & b[287])^(a[50] & b[288])^(a[49] & b[289])^(a[48] & b[290])^(a[47] & b[291])^(a[46] & b[292])^(a[45] & b[293])^(a[44] & b[294])^(a[43] & b[295])^(a[42] & b[296])^(a[41] & b[297])^(a[40] & b[298])^(a[39] & b[299])^(a[38] & b[300])^(a[37] & b[301])^(a[36] & b[302])^(a[35] & b[303])^(a[34] & b[304])^(a[33] & b[305])^(a[32] & b[306])^(a[31] & b[307])^(a[30] & b[308])^(a[29] & b[309])^(a[28] & b[310])^(a[27] & b[311])^(a[26] & b[312])^(a[25] & b[313])^(a[24] & b[314])^(a[23] & b[315])^(a[22] & b[316])^(a[21] & b[317])^(a[20] & b[318])^(a[19] & b[319])^(a[18] & b[320])^(a[17] & b[321])^(a[16] & b[322])^(a[15] & b[323])^(a[14] & b[324])^(a[13] & b[325])^(a[12] & b[326])^(a[11] & b[327])^(a[10] & b[328])^(a[9] & b[329])^(a[8] & b[330])^(a[7] & b[331])^(a[6] & b[332])^(a[5] & b[333])^(a[4] & b[334])^(a[3] & b[335])^(a[2] & b[336])^(a[1] & b[337])^(a[0] & b[338]);
assign y[339] = (a[339] & b[0])^(a[338] & b[1])^(a[337] & b[2])^(a[336] & b[3])^(a[335] & b[4])^(a[334] & b[5])^(a[333] & b[6])^(a[332] & b[7])^(a[331] & b[8])^(a[330] & b[9])^(a[329] & b[10])^(a[328] & b[11])^(a[327] & b[12])^(a[326] & b[13])^(a[325] & b[14])^(a[324] & b[15])^(a[323] & b[16])^(a[322] & b[17])^(a[321] & b[18])^(a[320] & b[19])^(a[319] & b[20])^(a[318] & b[21])^(a[317] & b[22])^(a[316] & b[23])^(a[315] & b[24])^(a[314] & b[25])^(a[313] & b[26])^(a[312] & b[27])^(a[311] & b[28])^(a[310] & b[29])^(a[309] & b[30])^(a[308] & b[31])^(a[307] & b[32])^(a[306] & b[33])^(a[305] & b[34])^(a[304] & b[35])^(a[303] & b[36])^(a[302] & b[37])^(a[301] & b[38])^(a[300] & b[39])^(a[299] & b[40])^(a[298] & b[41])^(a[297] & b[42])^(a[296] & b[43])^(a[295] & b[44])^(a[294] & b[45])^(a[293] & b[46])^(a[292] & b[47])^(a[291] & b[48])^(a[290] & b[49])^(a[289] & b[50])^(a[288] & b[51])^(a[287] & b[52])^(a[286] & b[53])^(a[285] & b[54])^(a[284] & b[55])^(a[283] & b[56])^(a[282] & b[57])^(a[281] & b[58])^(a[280] & b[59])^(a[279] & b[60])^(a[278] & b[61])^(a[277] & b[62])^(a[276] & b[63])^(a[275] & b[64])^(a[274] & b[65])^(a[273] & b[66])^(a[272] & b[67])^(a[271] & b[68])^(a[270] & b[69])^(a[269] & b[70])^(a[268] & b[71])^(a[267] & b[72])^(a[266] & b[73])^(a[265] & b[74])^(a[264] & b[75])^(a[263] & b[76])^(a[262] & b[77])^(a[261] & b[78])^(a[260] & b[79])^(a[259] & b[80])^(a[258] & b[81])^(a[257] & b[82])^(a[256] & b[83])^(a[255] & b[84])^(a[254] & b[85])^(a[253] & b[86])^(a[252] & b[87])^(a[251] & b[88])^(a[250] & b[89])^(a[249] & b[90])^(a[248] & b[91])^(a[247] & b[92])^(a[246] & b[93])^(a[245] & b[94])^(a[244] & b[95])^(a[243] & b[96])^(a[242] & b[97])^(a[241] & b[98])^(a[240] & b[99])^(a[239] & b[100])^(a[238] & b[101])^(a[237] & b[102])^(a[236] & b[103])^(a[235] & b[104])^(a[234] & b[105])^(a[233] & b[106])^(a[232] & b[107])^(a[231] & b[108])^(a[230] & b[109])^(a[229] & b[110])^(a[228] & b[111])^(a[227] & b[112])^(a[226] & b[113])^(a[225] & b[114])^(a[224] & b[115])^(a[223] & b[116])^(a[222] & b[117])^(a[221] & b[118])^(a[220] & b[119])^(a[219] & b[120])^(a[218] & b[121])^(a[217] & b[122])^(a[216] & b[123])^(a[215] & b[124])^(a[214] & b[125])^(a[213] & b[126])^(a[212] & b[127])^(a[211] & b[128])^(a[210] & b[129])^(a[209] & b[130])^(a[208] & b[131])^(a[207] & b[132])^(a[206] & b[133])^(a[205] & b[134])^(a[204] & b[135])^(a[203] & b[136])^(a[202] & b[137])^(a[201] & b[138])^(a[200] & b[139])^(a[199] & b[140])^(a[198] & b[141])^(a[197] & b[142])^(a[196] & b[143])^(a[195] & b[144])^(a[194] & b[145])^(a[193] & b[146])^(a[192] & b[147])^(a[191] & b[148])^(a[190] & b[149])^(a[189] & b[150])^(a[188] & b[151])^(a[187] & b[152])^(a[186] & b[153])^(a[185] & b[154])^(a[184] & b[155])^(a[183] & b[156])^(a[182] & b[157])^(a[181] & b[158])^(a[180] & b[159])^(a[179] & b[160])^(a[178] & b[161])^(a[177] & b[162])^(a[176] & b[163])^(a[175] & b[164])^(a[174] & b[165])^(a[173] & b[166])^(a[172] & b[167])^(a[171] & b[168])^(a[170] & b[169])^(a[169] & b[170])^(a[168] & b[171])^(a[167] & b[172])^(a[166] & b[173])^(a[165] & b[174])^(a[164] & b[175])^(a[163] & b[176])^(a[162] & b[177])^(a[161] & b[178])^(a[160] & b[179])^(a[159] & b[180])^(a[158] & b[181])^(a[157] & b[182])^(a[156] & b[183])^(a[155] & b[184])^(a[154] & b[185])^(a[153] & b[186])^(a[152] & b[187])^(a[151] & b[188])^(a[150] & b[189])^(a[149] & b[190])^(a[148] & b[191])^(a[147] & b[192])^(a[146] & b[193])^(a[145] & b[194])^(a[144] & b[195])^(a[143] & b[196])^(a[142] & b[197])^(a[141] & b[198])^(a[140] & b[199])^(a[139] & b[200])^(a[138] & b[201])^(a[137] & b[202])^(a[136] & b[203])^(a[135] & b[204])^(a[134] & b[205])^(a[133] & b[206])^(a[132] & b[207])^(a[131] & b[208])^(a[130] & b[209])^(a[129] & b[210])^(a[128] & b[211])^(a[127] & b[212])^(a[126] & b[213])^(a[125] & b[214])^(a[124] & b[215])^(a[123] & b[216])^(a[122] & b[217])^(a[121] & b[218])^(a[120] & b[219])^(a[119] & b[220])^(a[118] & b[221])^(a[117] & b[222])^(a[116] & b[223])^(a[115] & b[224])^(a[114] & b[225])^(a[113] & b[226])^(a[112] & b[227])^(a[111] & b[228])^(a[110] & b[229])^(a[109] & b[230])^(a[108] & b[231])^(a[107] & b[232])^(a[106] & b[233])^(a[105] & b[234])^(a[104] & b[235])^(a[103] & b[236])^(a[102] & b[237])^(a[101] & b[238])^(a[100] & b[239])^(a[99] & b[240])^(a[98] & b[241])^(a[97] & b[242])^(a[96] & b[243])^(a[95] & b[244])^(a[94] & b[245])^(a[93] & b[246])^(a[92] & b[247])^(a[91] & b[248])^(a[90] & b[249])^(a[89] & b[250])^(a[88] & b[251])^(a[87] & b[252])^(a[86] & b[253])^(a[85] & b[254])^(a[84] & b[255])^(a[83] & b[256])^(a[82] & b[257])^(a[81] & b[258])^(a[80] & b[259])^(a[79] & b[260])^(a[78] & b[261])^(a[77] & b[262])^(a[76] & b[263])^(a[75] & b[264])^(a[74] & b[265])^(a[73] & b[266])^(a[72] & b[267])^(a[71] & b[268])^(a[70] & b[269])^(a[69] & b[270])^(a[68] & b[271])^(a[67] & b[272])^(a[66] & b[273])^(a[65] & b[274])^(a[64] & b[275])^(a[63] & b[276])^(a[62] & b[277])^(a[61] & b[278])^(a[60] & b[279])^(a[59] & b[280])^(a[58] & b[281])^(a[57] & b[282])^(a[56] & b[283])^(a[55] & b[284])^(a[54] & b[285])^(a[53] & b[286])^(a[52] & b[287])^(a[51] & b[288])^(a[50] & b[289])^(a[49] & b[290])^(a[48] & b[291])^(a[47] & b[292])^(a[46] & b[293])^(a[45] & b[294])^(a[44] & b[295])^(a[43] & b[296])^(a[42] & b[297])^(a[41] & b[298])^(a[40] & b[299])^(a[39] & b[300])^(a[38] & b[301])^(a[37] & b[302])^(a[36] & b[303])^(a[35] & b[304])^(a[34] & b[305])^(a[33] & b[306])^(a[32] & b[307])^(a[31] & b[308])^(a[30] & b[309])^(a[29] & b[310])^(a[28] & b[311])^(a[27] & b[312])^(a[26] & b[313])^(a[25] & b[314])^(a[24] & b[315])^(a[23] & b[316])^(a[22] & b[317])^(a[21] & b[318])^(a[20] & b[319])^(a[19] & b[320])^(a[18] & b[321])^(a[17] & b[322])^(a[16] & b[323])^(a[15] & b[324])^(a[14] & b[325])^(a[13] & b[326])^(a[12] & b[327])^(a[11] & b[328])^(a[10] & b[329])^(a[9] & b[330])^(a[8] & b[331])^(a[7] & b[332])^(a[6] & b[333])^(a[5] & b[334])^(a[4] & b[335])^(a[3] & b[336])^(a[2] & b[337])^(a[1] & b[338])^(a[0] & b[339]);
assign y[340] = (a[340] & b[0])^(a[339] & b[1])^(a[338] & b[2])^(a[337] & b[3])^(a[336] & b[4])^(a[335] & b[5])^(a[334] & b[6])^(a[333] & b[7])^(a[332] & b[8])^(a[331] & b[9])^(a[330] & b[10])^(a[329] & b[11])^(a[328] & b[12])^(a[327] & b[13])^(a[326] & b[14])^(a[325] & b[15])^(a[324] & b[16])^(a[323] & b[17])^(a[322] & b[18])^(a[321] & b[19])^(a[320] & b[20])^(a[319] & b[21])^(a[318] & b[22])^(a[317] & b[23])^(a[316] & b[24])^(a[315] & b[25])^(a[314] & b[26])^(a[313] & b[27])^(a[312] & b[28])^(a[311] & b[29])^(a[310] & b[30])^(a[309] & b[31])^(a[308] & b[32])^(a[307] & b[33])^(a[306] & b[34])^(a[305] & b[35])^(a[304] & b[36])^(a[303] & b[37])^(a[302] & b[38])^(a[301] & b[39])^(a[300] & b[40])^(a[299] & b[41])^(a[298] & b[42])^(a[297] & b[43])^(a[296] & b[44])^(a[295] & b[45])^(a[294] & b[46])^(a[293] & b[47])^(a[292] & b[48])^(a[291] & b[49])^(a[290] & b[50])^(a[289] & b[51])^(a[288] & b[52])^(a[287] & b[53])^(a[286] & b[54])^(a[285] & b[55])^(a[284] & b[56])^(a[283] & b[57])^(a[282] & b[58])^(a[281] & b[59])^(a[280] & b[60])^(a[279] & b[61])^(a[278] & b[62])^(a[277] & b[63])^(a[276] & b[64])^(a[275] & b[65])^(a[274] & b[66])^(a[273] & b[67])^(a[272] & b[68])^(a[271] & b[69])^(a[270] & b[70])^(a[269] & b[71])^(a[268] & b[72])^(a[267] & b[73])^(a[266] & b[74])^(a[265] & b[75])^(a[264] & b[76])^(a[263] & b[77])^(a[262] & b[78])^(a[261] & b[79])^(a[260] & b[80])^(a[259] & b[81])^(a[258] & b[82])^(a[257] & b[83])^(a[256] & b[84])^(a[255] & b[85])^(a[254] & b[86])^(a[253] & b[87])^(a[252] & b[88])^(a[251] & b[89])^(a[250] & b[90])^(a[249] & b[91])^(a[248] & b[92])^(a[247] & b[93])^(a[246] & b[94])^(a[245] & b[95])^(a[244] & b[96])^(a[243] & b[97])^(a[242] & b[98])^(a[241] & b[99])^(a[240] & b[100])^(a[239] & b[101])^(a[238] & b[102])^(a[237] & b[103])^(a[236] & b[104])^(a[235] & b[105])^(a[234] & b[106])^(a[233] & b[107])^(a[232] & b[108])^(a[231] & b[109])^(a[230] & b[110])^(a[229] & b[111])^(a[228] & b[112])^(a[227] & b[113])^(a[226] & b[114])^(a[225] & b[115])^(a[224] & b[116])^(a[223] & b[117])^(a[222] & b[118])^(a[221] & b[119])^(a[220] & b[120])^(a[219] & b[121])^(a[218] & b[122])^(a[217] & b[123])^(a[216] & b[124])^(a[215] & b[125])^(a[214] & b[126])^(a[213] & b[127])^(a[212] & b[128])^(a[211] & b[129])^(a[210] & b[130])^(a[209] & b[131])^(a[208] & b[132])^(a[207] & b[133])^(a[206] & b[134])^(a[205] & b[135])^(a[204] & b[136])^(a[203] & b[137])^(a[202] & b[138])^(a[201] & b[139])^(a[200] & b[140])^(a[199] & b[141])^(a[198] & b[142])^(a[197] & b[143])^(a[196] & b[144])^(a[195] & b[145])^(a[194] & b[146])^(a[193] & b[147])^(a[192] & b[148])^(a[191] & b[149])^(a[190] & b[150])^(a[189] & b[151])^(a[188] & b[152])^(a[187] & b[153])^(a[186] & b[154])^(a[185] & b[155])^(a[184] & b[156])^(a[183] & b[157])^(a[182] & b[158])^(a[181] & b[159])^(a[180] & b[160])^(a[179] & b[161])^(a[178] & b[162])^(a[177] & b[163])^(a[176] & b[164])^(a[175] & b[165])^(a[174] & b[166])^(a[173] & b[167])^(a[172] & b[168])^(a[171] & b[169])^(a[170] & b[170])^(a[169] & b[171])^(a[168] & b[172])^(a[167] & b[173])^(a[166] & b[174])^(a[165] & b[175])^(a[164] & b[176])^(a[163] & b[177])^(a[162] & b[178])^(a[161] & b[179])^(a[160] & b[180])^(a[159] & b[181])^(a[158] & b[182])^(a[157] & b[183])^(a[156] & b[184])^(a[155] & b[185])^(a[154] & b[186])^(a[153] & b[187])^(a[152] & b[188])^(a[151] & b[189])^(a[150] & b[190])^(a[149] & b[191])^(a[148] & b[192])^(a[147] & b[193])^(a[146] & b[194])^(a[145] & b[195])^(a[144] & b[196])^(a[143] & b[197])^(a[142] & b[198])^(a[141] & b[199])^(a[140] & b[200])^(a[139] & b[201])^(a[138] & b[202])^(a[137] & b[203])^(a[136] & b[204])^(a[135] & b[205])^(a[134] & b[206])^(a[133] & b[207])^(a[132] & b[208])^(a[131] & b[209])^(a[130] & b[210])^(a[129] & b[211])^(a[128] & b[212])^(a[127] & b[213])^(a[126] & b[214])^(a[125] & b[215])^(a[124] & b[216])^(a[123] & b[217])^(a[122] & b[218])^(a[121] & b[219])^(a[120] & b[220])^(a[119] & b[221])^(a[118] & b[222])^(a[117] & b[223])^(a[116] & b[224])^(a[115] & b[225])^(a[114] & b[226])^(a[113] & b[227])^(a[112] & b[228])^(a[111] & b[229])^(a[110] & b[230])^(a[109] & b[231])^(a[108] & b[232])^(a[107] & b[233])^(a[106] & b[234])^(a[105] & b[235])^(a[104] & b[236])^(a[103] & b[237])^(a[102] & b[238])^(a[101] & b[239])^(a[100] & b[240])^(a[99] & b[241])^(a[98] & b[242])^(a[97] & b[243])^(a[96] & b[244])^(a[95] & b[245])^(a[94] & b[246])^(a[93] & b[247])^(a[92] & b[248])^(a[91] & b[249])^(a[90] & b[250])^(a[89] & b[251])^(a[88] & b[252])^(a[87] & b[253])^(a[86] & b[254])^(a[85] & b[255])^(a[84] & b[256])^(a[83] & b[257])^(a[82] & b[258])^(a[81] & b[259])^(a[80] & b[260])^(a[79] & b[261])^(a[78] & b[262])^(a[77] & b[263])^(a[76] & b[264])^(a[75] & b[265])^(a[74] & b[266])^(a[73] & b[267])^(a[72] & b[268])^(a[71] & b[269])^(a[70] & b[270])^(a[69] & b[271])^(a[68] & b[272])^(a[67] & b[273])^(a[66] & b[274])^(a[65] & b[275])^(a[64] & b[276])^(a[63] & b[277])^(a[62] & b[278])^(a[61] & b[279])^(a[60] & b[280])^(a[59] & b[281])^(a[58] & b[282])^(a[57] & b[283])^(a[56] & b[284])^(a[55] & b[285])^(a[54] & b[286])^(a[53] & b[287])^(a[52] & b[288])^(a[51] & b[289])^(a[50] & b[290])^(a[49] & b[291])^(a[48] & b[292])^(a[47] & b[293])^(a[46] & b[294])^(a[45] & b[295])^(a[44] & b[296])^(a[43] & b[297])^(a[42] & b[298])^(a[41] & b[299])^(a[40] & b[300])^(a[39] & b[301])^(a[38] & b[302])^(a[37] & b[303])^(a[36] & b[304])^(a[35] & b[305])^(a[34] & b[306])^(a[33] & b[307])^(a[32] & b[308])^(a[31] & b[309])^(a[30] & b[310])^(a[29] & b[311])^(a[28] & b[312])^(a[27] & b[313])^(a[26] & b[314])^(a[25] & b[315])^(a[24] & b[316])^(a[23] & b[317])^(a[22] & b[318])^(a[21] & b[319])^(a[20] & b[320])^(a[19] & b[321])^(a[18] & b[322])^(a[17] & b[323])^(a[16] & b[324])^(a[15] & b[325])^(a[14] & b[326])^(a[13] & b[327])^(a[12] & b[328])^(a[11] & b[329])^(a[10] & b[330])^(a[9] & b[331])^(a[8] & b[332])^(a[7] & b[333])^(a[6] & b[334])^(a[5] & b[335])^(a[4] & b[336])^(a[3] & b[337])^(a[2] & b[338])^(a[1] & b[339])^(a[0] & b[340]);
assign y[341] = (a[341] & b[0])^(a[340] & b[1])^(a[339] & b[2])^(a[338] & b[3])^(a[337] & b[4])^(a[336] & b[5])^(a[335] & b[6])^(a[334] & b[7])^(a[333] & b[8])^(a[332] & b[9])^(a[331] & b[10])^(a[330] & b[11])^(a[329] & b[12])^(a[328] & b[13])^(a[327] & b[14])^(a[326] & b[15])^(a[325] & b[16])^(a[324] & b[17])^(a[323] & b[18])^(a[322] & b[19])^(a[321] & b[20])^(a[320] & b[21])^(a[319] & b[22])^(a[318] & b[23])^(a[317] & b[24])^(a[316] & b[25])^(a[315] & b[26])^(a[314] & b[27])^(a[313] & b[28])^(a[312] & b[29])^(a[311] & b[30])^(a[310] & b[31])^(a[309] & b[32])^(a[308] & b[33])^(a[307] & b[34])^(a[306] & b[35])^(a[305] & b[36])^(a[304] & b[37])^(a[303] & b[38])^(a[302] & b[39])^(a[301] & b[40])^(a[300] & b[41])^(a[299] & b[42])^(a[298] & b[43])^(a[297] & b[44])^(a[296] & b[45])^(a[295] & b[46])^(a[294] & b[47])^(a[293] & b[48])^(a[292] & b[49])^(a[291] & b[50])^(a[290] & b[51])^(a[289] & b[52])^(a[288] & b[53])^(a[287] & b[54])^(a[286] & b[55])^(a[285] & b[56])^(a[284] & b[57])^(a[283] & b[58])^(a[282] & b[59])^(a[281] & b[60])^(a[280] & b[61])^(a[279] & b[62])^(a[278] & b[63])^(a[277] & b[64])^(a[276] & b[65])^(a[275] & b[66])^(a[274] & b[67])^(a[273] & b[68])^(a[272] & b[69])^(a[271] & b[70])^(a[270] & b[71])^(a[269] & b[72])^(a[268] & b[73])^(a[267] & b[74])^(a[266] & b[75])^(a[265] & b[76])^(a[264] & b[77])^(a[263] & b[78])^(a[262] & b[79])^(a[261] & b[80])^(a[260] & b[81])^(a[259] & b[82])^(a[258] & b[83])^(a[257] & b[84])^(a[256] & b[85])^(a[255] & b[86])^(a[254] & b[87])^(a[253] & b[88])^(a[252] & b[89])^(a[251] & b[90])^(a[250] & b[91])^(a[249] & b[92])^(a[248] & b[93])^(a[247] & b[94])^(a[246] & b[95])^(a[245] & b[96])^(a[244] & b[97])^(a[243] & b[98])^(a[242] & b[99])^(a[241] & b[100])^(a[240] & b[101])^(a[239] & b[102])^(a[238] & b[103])^(a[237] & b[104])^(a[236] & b[105])^(a[235] & b[106])^(a[234] & b[107])^(a[233] & b[108])^(a[232] & b[109])^(a[231] & b[110])^(a[230] & b[111])^(a[229] & b[112])^(a[228] & b[113])^(a[227] & b[114])^(a[226] & b[115])^(a[225] & b[116])^(a[224] & b[117])^(a[223] & b[118])^(a[222] & b[119])^(a[221] & b[120])^(a[220] & b[121])^(a[219] & b[122])^(a[218] & b[123])^(a[217] & b[124])^(a[216] & b[125])^(a[215] & b[126])^(a[214] & b[127])^(a[213] & b[128])^(a[212] & b[129])^(a[211] & b[130])^(a[210] & b[131])^(a[209] & b[132])^(a[208] & b[133])^(a[207] & b[134])^(a[206] & b[135])^(a[205] & b[136])^(a[204] & b[137])^(a[203] & b[138])^(a[202] & b[139])^(a[201] & b[140])^(a[200] & b[141])^(a[199] & b[142])^(a[198] & b[143])^(a[197] & b[144])^(a[196] & b[145])^(a[195] & b[146])^(a[194] & b[147])^(a[193] & b[148])^(a[192] & b[149])^(a[191] & b[150])^(a[190] & b[151])^(a[189] & b[152])^(a[188] & b[153])^(a[187] & b[154])^(a[186] & b[155])^(a[185] & b[156])^(a[184] & b[157])^(a[183] & b[158])^(a[182] & b[159])^(a[181] & b[160])^(a[180] & b[161])^(a[179] & b[162])^(a[178] & b[163])^(a[177] & b[164])^(a[176] & b[165])^(a[175] & b[166])^(a[174] & b[167])^(a[173] & b[168])^(a[172] & b[169])^(a[171] & b[170])^(a[170] & b[171])^(a[169] & b[172])^(a[168] & b[173])^(a[167] & b[174])^(a[166] & b[175])^(a[165] & b[176])^(a[164] & b[177])^(a[163] & b[178])^(a[162] & b[179])^(a[161] & b[180])^(a[160] & b[181])^(a[159] & b[182])^(a[158] & b[183])^(a[157] & b[184])^(a[156] & b[185])^(a[155] & b[186])^(a[154] & b[187])^(a[153] & b[188])^(a[152] & b[189])^(a[151] & b[190])^(a[150] & b[191])^(a[149] & b[192])^(a[148] & b[193])^(a[147] & b[194])^(a[146] & b[195])^(a[145] & b[196])^(a[144] & b[197])^(a[143] & b[198])^(a[142] & b[199])^(a[141] & b[200])^(a[140] & b[201])^(a[139] & b[202])^(a[138] & b[203])^(a[137] & b[204])^(a[136] & b[205])^(a[135] & b[206])^(a[134] & b[207])^(a[133] & b[208])^(a[132] & b[209])^(a[131] & b[210])^(a[130] & b[211])^(a[129] & b[212])^(a[128] & b[213])^(a[127] & b[214])^(a[126] & b[215])^(a[125] & b[216])^(a[124] & b[217])^(a[123] & b[218])^(a[122] & b[219])^(a[121] & b[220])^(a[120] & b[221])^(a[119] & b[222])^(a[118] & b[223])^(a[117] & b[224])^(a[116] & b[225])^(a[115] & b[226])^(a[114] & b[227])^(a[113] & b[228])^(a[112] & b[229])^(a[111] & b[230])^(a[110] & b[231])^(a[109] & b[232])^(a[108] & b[233])^(a[107] & b[234])^(a[106] & b[235])^(a[105] & b[236])^(a[104] & b[237])^(a[103] & b[238])^(a[102] & b[239])^(a[101] & b[240])^(a[100] & b[241])^(a[99] & b[242])^(a[98] & b[243])^(a[97] & b[244])^(a[96] & b[245])^(a[95] & b[246])^(a[94] & b[247])^(a[93] & b[248])^(a[92] & b[249])^(a[91] & b[250])^(a[90] & b[251])^(a[89] & b[252])^(a[88] & b[253])^(a[87] & b[254])^(a[86] & b[255])^(a[85] & b[256])^(a[84] & b[257])^(a[83] & b[258])^(a[82] & b[259])^(a[81] & b[260])^(a[80] & b[261])^(a[79] & b[262])^(a[78] & b[263])^(a[77] & b[264])^(a[76] & b[265])^(a[75] & b[266])^(a[74] & b[267])^(a[73] & b[268])^(a[72] & b[269])^(a[71] & b[270])^(a[70] & b[271])^(a[69] & b[272])^(a[68] & b[273])^(a[67] & b[274])^(a[66] & b[275])^(a[65] & b[276])^(a[64] & b[277])^(a[63] & b[278])^(a[62] & b[279])^(a[61] & b[280])^(a[60] & b[281])^(a[59] & b[282])^(a[58] & b[283])^(a[57] & b[284])^(a[56] & b[285])^(a[55] & b[286])^(a[54] & b[287])^(a[53] & b[288])^(a[52] & b[289])^(a[51] & b[290])^(a[50] & b[291])^(a[49] & b[292])^(a[48] & b[293])^(a[47] & b[294])^(a[46] & b[295])^(a[45] & b[296])^(a[44] & b[297])^(a[43] & b[298])^(a[42] & b[299])^(a[41] & b[300])^(a[40] & b[301])^(a[39] & b[302])^(a[38] & b[303])^(a[37] & b[304])^(a[36] & b[305])^(a[35] & b[306])^(a[34] & b[307])^(a[33] & b[308])^(a[32] & b[309])^(a[31] & b[310])^(a[30] & b[311])^(a[29] & b[312])^(a[28] & b[313])^(a[27] & b[314])^(a[26] & b[315])^(a[25] & b[316])^(a[24] & b[317])^(a[23] & b[318])^(a[22] & b[319])^(a[21] & b[320])^(a[20] & b[321])^(a[19] & b[322])^(a[18] & b[323])^(a[17] & b[324])^(a[16] & b[325])^(a[15] & b[326])^(a[14] & b[327])^(a[13] & b[328])^(a[12] & b[329])^(a[11] & b[330])^(a[10] & b[331])^(a[9] & b[332])^(a[8] & b[333])^(a[7] & b[334])^(a[6] & b[335])^(a[5] & b[336])^(a[4] & b[337])^(a[3] & b[338])^(a[2] & b[339])^(a[1] & b[340])^(a[0] & b[341]);
assign y[342] = (a[342] & b[0])^(a[341] & b[1])^(a[340] & b[2])^(a[339] & b[3])^(a[338] & b[4])^(a[337] & b[5])^(a[336] & b[6])^(a[335] & b[7])^(a[334] & b[8])^(a[333] & b[9])^(a[332] & b[10])^(a[331] & b[11])^(a[330] & b[12])^(a[329] & b[13])^(a[328] & b[14])^(a[327] & b[15])^(a[326] & b[16])^(a[325] & b[17])^(a[324] & b[18])^(a[323] & b[19])^(a[322] & b[20])^(a[321] & b[21])^(a[320] & b[22])^(a[319] & b[23])^(a[318] & b[24])^(a[317] & b[25])^(a[316] & b[26])^(a[315] & b[27])^(a[314] & b[28])^(a[313] & b[29])^(a[312] & b[30])^(a[311] & b[31])^(a[310] & b[32])^(a[309] & b[33])^(a[308] & b[34])^(a[307] & b[35])^(a[306] & b[36])^(a[305] & b[37])^(a[304] & b[38])^(a[303] & b[39])^(a[302] & b[40])^(a[301] & b[41])^(a[300] & b[42])^(a[299] & b[43])^(a[298] & b[44])^(a[297] & b[45])^(a[296] & b[46])^(a[295] & b[47])^(a[294] & b[48])^(a[293] & b[49])^(a[292] & b[50])^(a[291] & b[51])^(a[290] & b[52])^(a[289] & b[53])^(a[288] & b[54])^(a[287] & b[55])^(a[286] & b[56])^(a[285] & b[57])^(a[284] & b[58])^(a[283] & b[59])^(a[282] & b[60])^(a[281] & b[61])^(a[280] & b[62])^(a[279] & b[63])^(a[278] & b[64])^(a[277] & b[65])^(a[276] & b[66])^(a[275] & b[67])^(a[274] & b[68])^(a[273] & b[69])^(a[272] & b[70])^(a[271] & b[71])^(a[270] & b[72])^(a[269] & b[73])^(a[268] & b[74])^(a[267] & b[75])^(a[266] & b[76])^(a[265] & b[77])^(a[264] & b[78])^(a[263] & b[79])^(a[262] & b[80])^(a[261] & b[81])^(a[260] & b[82])^(a[259] & b[83])^(a[258] & b[84])^(a[257] & b[85])^(a[256] & b[86])^(a[255] & b[87])^(a[254] & b[88])^(a[253] & b[89])^(a[252] & b[90])^(a[251] & b[91])^(a[250] & b[92])^(a[249] & b[93])^(a[248] & b[94])^(a[247] & b[95])^(a[246] & b[96])^(a[245] & b[97])^(a[244] & b[98])^(a[243] & b[99])^(a[242] & b[100])^(a[241] & b[101])^(a[240] & b[102])^(a[239] & b[103])^(a[238] & b[104])^(a[237] & b[105])^(a[236] & b[106])^(a[235] & b[107])^(a[234] & b[108])^(a[233] & b[109])^(a[232] & b[110])^(a[231] & b[111])^(a[230] & b[112])^(a[229] & b[113])^(a[228] & b[114])^(a[227] & b[115])^(a[226] & b[116])^(a[225] & b[117])^(a[224] & b[118])^(a[223] & b[119])^(a[222] & b[120])^(a[221] & b[121])^(a[220] & b[122])^(a[219] & b[123])^(a[218] & b[124])^(a[217] & b[125])^(a[216] & b[126])^(a[215] & b[127])^(a[214] & b[128])^(a[213] & b[129])^(a[212] & b[130])^(a[211] & b[131])^(a[210] & b[132])^(a[209] & b[133])^(a[208] & b[134])^(a[207] & b[135])^(a[206] & b[136])^(a[205] & b[137])^(a[204] & b[138])^(a[203] & b[139])^(a[202] & b[140])^(a[201] & b[141])^(a[200] & b[142])^(a[199] & b[143])^(a[198] & b[144])^(a[197] & b[145])^(a[196] & b[146])^(a[195] & b[147])^(a[194] & b[148])^(a[193] & b[149])^(a[192] & b[150])^(a[191] & b[151])^(a[190] & b[152])^(a[189] & b[153])^(a[188] & b[154])^(a[187] & b[155])^(a[186] & b[156])^(a[185] & b[157])^(a[184] & b[158])^(a[183] & b[159])^(a[182] & b[160])^(a[181] & b[161])^(a[180] & b[162])^(a[179] & b[163])^(a[178] & b[164])^(a[177] & b[165])^(a[176] & b[166])^(a[175] & b[167])^(a[174] & b[168])^(a[173] & b[169])^(a[172] & b[170])^(a[171] & b[171])^(a[170] & b[172])^(a[169] & b[173])^(a[168] & b[174])^(a[167] & b[175])^(a[166] & b[176])^(a[165] & b[177])^(a[164] & b[178])^(a[163] & b[179])^(a[162] & b[180])^(a[161] & b[181])^(a[160] & b[182])^(a[159] & b[183])^(a[158] & b[184])^(a[157] & b[185])^(a[156] & b[186])^(a[155] & b[187])^(a[154] & b[188])^(a[153] & b[189])^(a[152] & b[190])^(a[151] & b[191])^(a[150] & b[192])^(a[149] & b[193])^(a[148] & b[194])^(a[147] & b[195])^(a[146] & b[196])^(a[145] & b[197])^(a[144] & b[198])^(a[143] & b[199])^(a[142] & b[200])^(a[141] & b[201])^(a[140] & b[202])^(a[139] & b[203])^(a[138] & b[204])^(a[137] & b[205])^(a[136] & b[206])^(a[135] & b[207])^(a[134] & b[208])^(a[133] & b[209])^(a[132] & b[210])^(a[131] & b[211])^(a[130] & b[212])^(a[129] & b[213])^(a[128] & b[214])^(a[127] & b[215])^(a[126] & b[216])^(a[125] & b[217])^(a[124] & b[218])^(a[123] & b[219])^(a[122] & b[220])^(a[121] & b[221])^(a[120] & b[222])^(a[119] & b[223])^(a[118] & b[224])^(a[117] & b[225])^(a[116] & b[226])^(a[115] & b[227])^(a[114] & b[228])^(a[113] & b[229])^(a[112] & b[230])^(a[111] & b[231])^(a[110] & b[232])^(a[109] & b[233])^(a[108] & b[234])^(a[107] & b[235])^(a[106] & b[236])^(a[105] & b[237])^(a[104] & b[238])^(a[103] & b[239])^(a[102] & b[240])^(a[101] & b[241])^(a[100] & b[242])^(a[99] & b[243])^(a[98] & b[244])^(a[97] & b[245])^(a[96] & b[246])^(a[95] & b[247])^(a[94] & b[248])^(a[93] & b[249])^(a[92] & b[250])^(a[91] & b[251])^(a[90] & b[252])^(a[89] & b[253])^(a[88] & b[254])^(a[87] & b[255])^(a[86] & b[256])^(a[85] & b[257])^(a[84] & b[258])^(a[83] & b[259])^(a[82] & b[260])^(a[81] & b[261])^(a[80] & b[262])^(a[79] & b[263])^(a[78] & b[264])^(a[77] & b[265])^(a[76] & b[266])^(a[75] & b[267])^(a[74] & b[268])^(a[73] & b[269])^(a[72] & b[270])^(a[71] & b[271])^(a[70] & b[272])^(a[69] & b[273])^(a[68] & b[274])^(a[67] & b[275])^(a[66] & b[276])^(a[65] & b[277])^(a[64] & b[278])^(a[63] & b[279])^(a[62] & b[280])^(a[61] & b[281])^(a[60] & b[282])^(a[59] & b[283])^(a[58] & b[284])^(a[57] & b[285])^(a[56] & b[286])^(a[55] & b[287])^(a[54] & b[288])^(a[53] & b[289])^(a[52] & b[290])^(a[51] & b[291])^(a[50] & b[292])^(a[49] & b[293])^(a[48] & b[294])^(a[47] & b[295])^(a[46] & b[296])^(a[45] & b[297])^(a[44] & b[298])^(a[43] & b[299])^(a[42] & b[300])^(a[41] & b[301])^(a[40] & b[302])^(a[39] & b[303])^(a[38] & b[304])^(a[37] & b[305])^(a[36] & b[306])^(a[35] & b[307])^(a[34] & b[308])^(a[33] & b[309])^(a[32] & b[310])^(a[31] & b[311])^(a[30] & b[312])^(a[29] & b[313])^(a[28] & b[314])^(a[27] & b[315])^(a[26] & b[316])^(a[25] & b[317])^(a[24] & b[318])^(a[23] & b[319])^(a[22] & b[320])^(a[21] & b[321])^(a[20] & b[322])^(a[19] & b[323])^(a[18] & b[324])^(a[17] & b[325])^(a[16] & b[326])^(a[15] & b[327])^(a[14] & b[328])^(a[13] & b[329])^(a[12] & b[330])^(a[11] & b[331])^(a[10] & b[332])^(a[9] & b[333])^(a[8] & b[334])^(a[7] & b[335])^(a[6] & b[336])^(a[5] & b[337])^(a[4] & b[338])^(a[3] & b[339])^(a[2] & b[340])^(a[1] & b[341])^(a[0] & b[342]);
assign y[343] = (a[343] & b[0])^(a[342] & b[1])^(a[341] & b[2])^(a[340] & b[3])^(a[339] & b[4])^(a[338] & b[5])^(a[337] & b[6])^(a[336] & b[7])^(a[335] & b[8])^(a[334] & b[9])^(a[333] & b[10])^(a[332] & b[11])^(a[331] & b[12])^(a[330] & b[13])^(a[329] & b[14])^(a[328] & b[15])^(a[327] & b[16])^(a[326] & b[17])^(a[325] & b[18])^(a[324] & b[19])^(a[323] & b[20])^(a[322] & b[21])^(a[321] & b[22])^(a[320] & b[23])^(a[319] & b[24])^(a[318] & b[25])^(a[317] & b[26])^(a[316] & b[27])^(a[315] & b[28])^(a[314] & b[29])^(a[313] & b[30])^(a[312] & b[31])^(a[311] & b[32])^(a[310] & b[33])^(a[309] & b[34])^(a[308] & b[35])^(a[307] & b[36])^(a[306] & b[37])^(a[305] & b[38])^(a[304] & b[39])^(a[303] & b[40])^(a[302] & b[41])^(a[301] & b[42])^(a[300] & b[43])^(a[299] & b[44])^(a[298] & b[45])^(a[297] & b[46])^(a[296] & b[47])^(a[295] & b[48])^(a[294] & b[49])^(a[293] & b[50])^(a[292] & b[51])^(a[291] & b[52])^(a[290] & b[53])^(a[289] & b[54])^(a[288] & b[55])^(a[287] & b[56])^(a[286] & b[57])^(a[285] & b[58])^(a[284] & b[59])^(a[283] & b[60])^(a[282] & b[61])^(a[281] & b[62])^(a[280] & b[63])^(a[279] & b[64])^(a[278] & b[65])^(a[277] & b[66])^(a[276] & b[67])^(a[275] & b[68])^(a[274] & b[69])^(a[273] & b[70])^(a[272] & b[71])^(a[271] & b[72])^(a[270] & b[73])^(a[269] & b[74])^(a[268] & b[75])^(a[267] & b[76])^(a[266] & b[77])^(a[265] & b[78])^(a[264] & b[79])^(a[263] & b[80])^(a[262] & b[81])^(a[261] & b[82])^(a[260] & b[83])^(a[259] & b[84])^(a[258] & b[85])^(a[257] & b[86])^(a[256] & b[87])^(a[255] & b[88])^(a[254] & b[89])^(a[253] & b[90])^(a[252] & b[91])^(a[251] & b[92])^(a[250] & b[93])^(a[249] & b[94])^(a[248] & b[95])^(a[247] & b[96])^(a[246] & b[97])^(a[245] & b[98])^(a[244] & b[99])^(a[243] & b[100])^(a[242] & b[101])^(a[241] & b[102])^(a[240] & b[103])^(a[239] & b[104])^(a[238] & b[105])^(a[237] & b[106])^(a[236] & b[107])^(a[235] & b[108])^(a[234] & b[109])^(a[233] & b[110])^(a[232] & b[111])^(a[231] & b[112])^(a[230] & b[113])^(a[229] & b[114])^(a[228] & b[115])^(a[227] & b[116])^(a[226] & b[117])^(a[225] & b[118])^(a[224] & b[119])^(a[223] & b[120])^(a[222] & b[121])^(a[221] & b[122])^(a[220] & b[123])^(a[219] & b[124])^(a[218] & b[125])^(a[217] & b[126])^(a[216] & b[127])^(a[215] & b[128])^(a[214] & b[129])^(a[213] & b[130])^(a[212] & b[131])^(a[211] & b[132])^(a[210] & b[133])^(a[209] & b[134])^(a[208] & b[135])^(a[207] & b[136])^(a[206] & b[137])^(a[205] & b[138])^(a[204] & b[139])^(a[203] & b[140])^(a[202] & b[141])^(a[201] & b[142])^(a[200] & b[143])^(a[199] & b[144])^(a[198] & b[145])^(a[197] & b[146])^(a[196] & b[147])^(a[195] & b[148])^(a[194] & b[149])^(a[193] & b[150])^(a[192] & b[151])^(a[191] & b[152])^(a[190] & b[153])^(a[189] & b[154])^(a[188] & b[155])^(a[187] & b[156])^(a[186] & b[157])^(a[185] & b[158])^(a[184] & b[159])^(a[183] & b[160])^(a[182] & b[161])^(a[181] & b[162])^(a[180] & b[163])^(a[179] & b[164])^(a[178] & b[165])^(a[177] & b[166])^(a[176] & b[167])^(a[175] & b[168])^(a[174] & b[169])^(a[173] & b[170])^(a[172] & b[171])^(a[171] & b[172])^(a[170] & b[173])^(a[169] & b[174])^(a[168] & b[175])^(a[167] & b[176])^(a[166] & b[177])^(a[165] & b[178])^(a[164] & b[179])^(a[163] & b[180])^(a[162] & b[181])^(a[161] & b[182])^(a[160] & b[183])^(a[159] & b[184])^(a[158] & b[185])^(a[157] & b[186])^(a[156] & b[187])^(a[155] & b[188])^(a[154] & b[189])^(a[153] & b[190])^(a[152] & b[191])^(a[151] & b[192])^(a[150] & b[193])^(a[149] & b[194])^(a[148] & b[195])^(a[147] & b[196])^(a[146] & b[197])^(a[145] & b[198])^(a[144] & b[199])^(a[143] & b[200])^(a[142] & b[201])^(a[141] & b[202])^(a[140] & b[203])^(a[139] & b[204])^(a[138] & b[205])^(a[137] & b[206])^(a[136] & b[207])^(a[135] & b[208])^(a[134] & b[209])^(a[133] & b[210])^(a[132] & b[211])^(a[131] & b[212])^(a[130] & b[213])^(a[129] & b[214])^(a[128] & b[215])^(a[127] & b[216])^(a[126] & b[217])^(a[125] & b[218])^(a[124] & b[219])^(a[123] & b[220])^(a[122] & b[221])^(a[121] & b[222])^(a[120] & b[223])^(a[119] & b[224])^(a[118] & b[225])^(a[117] & b[226])^(a[116] & b[227])^(a[115] & b[228])^(a[114] & b[229])^(a[113] & b[230])^(a[112] & b[231])^(a[111] & b[232])^(a[110] & b[233])^(a[109] & b[234])^(a[108] & b[235])^(a[107] & b[236])^(a[106] & b[237])^(a[105] & b[238])^(a[104] & b[239])^(a[103] & b[240])^(a[102] & b[241])^(a[101] & b[242])^(a[100] & b[243])^(a[99] & b[244])^(a[98] & b[245])^(a[97] & b[246])^(a[96] & b[247])^(a[95] & b[248])^(a[94] & b[249])^(a[93] & b[250])^(a[92] & b[251])^(a[91] & b[252])^(a[90] & b[253])^(a[89] & b[254])^(a[88] & b[255])^(a[87] & b[256])^(a[86] & b[257])^(a[85] & b[258])^(a[84] & b[259])^(a[83] & b[260])^(a[82] & b[261])^(a[81] & b[262])^(a[80] & b[263])^(a[79] & b[264])^(a[78] & b[265])^(a[77] & b[266])^(a[76] & b[267])^(a[75] & b[268])^(a[74] & b[269])^(a[73] & b[270])^(a[72] & b[271])^(a[71] & b[272])^(a[70] & b[273])^(a[69] & b[274])^(a[68] & b[275])^(a[67] & b[276])^(a[66] & b[277])^(a[65] & b[278])^(a[64] & b[279])^(a[63] & b[280])^(a[62] & b[281])^(a[61] & b[282])^(a[60] & b[283])^(a[59] & b[284])^(a[58] & b[285])^(a[57] & b[286])^(a[56] & b[287])^(a[55] & b[288])^(a[54] & b[289])^(a[53] & b[290])^(a[52] & b[291])^(a[51] & b[292])^(a[50] & b[293])^(a[49] & b[294])^(a[48] & b[295])^(a[47] & b[296])^(a[46] & b[297])^(a[45] & b[298])^(a[44] & b[299])^(a[43] & b[300])^(a[42] & b[301])^(a[41] & b[302])^(a[40] & b[303])^(a[39] & b[304])^(a[38] & b[305])^(a[37] & b[306])^(a[36] & b[307])^(a[35] & b[308])^(a[34] & b[309])^(a[33] & b[310])^(a[32] & b[311])^(a[31] & b[312])^(a[30] & b[313])^(a[29] & b[314])^(a[28] & b[315])^(a[27] & b[316])^(a[26] & b[317])^(a[25] & b[318])^(a[24] & b[319])^(a[23] & b[320])^(a[22] & b[321])^(a[21] & b[322])^(a[20] & b[323])^(a[19] & b[324])^(a[18] & b[325])^(a[17] & b[326])^(a[16] & b[327])^(a[15] & b[328])^(a[14] & b[329])^(a[13] & b[330])^(a[12] & b[331])^(a[11] & b[332])^(a[10] & b[333])^(a[9] & b[334])^(a[8] & b[335])^(a[7] & b[336])^(a[6] & b[337])^(a[5] & b[338])^(a[4] & b[339])^(a[3] & b[340])^(a[2] & b[341])^(a[1] & b[342])^(a[0] & b[343]);
assign y[344] = (a[344] & b[0])^(a[343] & b[1])^(a[342] & b[2])^(a[341] & b[3])^(a[340] & b[4])^(a[339] & b[5])^(a[338] & b[6])^(a[337] & b[7])^(a[336] & b[8])^(a[335] & b[9])^(a[334] & b[10])^(a[333] & b[11])^(a[332] & b[12])^(a[331] & b[13])^(a[330] & b[14])^(a[329] & b[15])^(a[328] & b[16])^(a[327] & b[17])^(a[326] & b[18])^(a[325] & b[19])^(a[324] & b[20])^(a[323] & b[21])^(a[322] & b[22])^(a[321] & b[23])^(a[320] & b[24])^(a[319] & b[25])^(a[318] & b[26])^(a[317] & b[27])^(a[316] & b[28])^(a[315] & b[29])^(a[314] & b[30])^(a[313] & b[31])^(a[312] & b[32])^(a[311] & b[33])^(a[310] & b[34])^(a[309] & b[35])^(a[308] & b[36])^(a[307] & b[37])^(a[306] & b[38])^(a[305] & b[39])^(a[304] & b[40])^(a[303] & b[41])^(a[302] & b[42])^(a[301] & b[43])^(a[300] & b[44])^(a[299] & b[45])^(a[298] & b[46])^(a[297] & b[47])^(a[296] & b[48])^(a[295] & b[49])^(a[294] & b[50])^(a[293] & b[51])^(a[292] & b[52])^(a[291] & b[53])^(a[290] & b[54])^(a[289] & b[55])^(a[288] & b[56])^(a[287] & b[57])^(a[286] & b[58])^(a[285] & b[59])^(a[284] & b[60])^(a[283] & b[61])^(a[282] & b[62])^(a[281] & b[63])^(a[280] & b[64])^(a[279] & b[65])^(a[278] & b[66])^(a[277] & b[67])^(a[276] & b[68])^(a[275] & b[69])^(a[274] & b[70])^(a[273] & b[71])^(a[272] & b[72])^(a[271] & b[73])^(a[270] & b[74])^(a[269] & b[75])^(a[268] & b[76])^(a[267] & b[77])^(a[266] & b[78])^(a[265] & b[79])^(a[264] & b[80])^(a[263] & b[81])^(a[262] & b[82])^(a[261] & b[83])^(a[260] & b[84])^(a[259] & b[85])^(a[258] & b[86])^(a[257] & b[87])^(a[256] & b[88])^(a[255] & b[89])^(a[254] & b[90])^(a[253] & b[91])^(a[252] & b[92])^(a[251] & b[93])^(a[250] & b[94])^(a[249] & b[95])^(a[248] & b[96])^(a[247] & b[97])^(a[246] & b[98])^(a[245] & b[99])^(a[244] & b[100])^(a[243] & b[101])^(a[242] & b[102])^(a[241] & b[103])^(a[240] & b[104])^(a[239] & b[105])^(a[238] & b[106])^(a[237] & b[107])^(a[236] & b[108])^(a[235] & b[109])^(a[234] & b[110])^(a[233] & b[111])^(a[232] & b[112])^(a[231] & b[113])^(a[230] & b[114])^(a[229] & b[115])^(a[228] & b[116])^(a[227] & b[117])^(a[226] & b[118])^(a[225] & b[119])^(a[224] & b[120])^(a[223] & b[121])^(a[222] & b[122])^(a[221] & b[123])^(a[220] & b[124])^(a[219] & b[125])^(a[218] & b[126])^(a[217] & b[127])^(a[216] & b[128])^(a[215] & b[129])^(a[214] & b[130])^(a[213] & b[131])^(a[212] & b[132])^(a[211] & b[133])^(a[210] & b[134])^(a[209] & b[135])^(a[208] & b[136])^(a[207] & b[137])^(a[206] & b[138])^(a[205] & b[139])^(a[204] & b[140])^(a[203] & b[141])^(a[202] & b[142])^(a[201] & b[143])^(a[200] & b[144])^(a[199] & b[145])^(a[198] & b[146])^(a[197] & b[147])^(a[196] & b[148])^(a[195] & b[149])^(a[194] & b[150])^(a[193] & b[151])^(a[192] & b[152])^(a[191] & b[153])^(a[190] & b[154])^(a[189] & b[155])^(a[188] & b[156])^(a[187] & b[157])^(a[186] & b[158])^(a[185] & b[159])^(a[184] & b[160])^(a[183] & b[161])^(a[182] & b[162])^(a[181] & b[163])^(a[180] & b[164])^(a[179] & b[165])^(a[178] & b[166])^(a[177] & b[167])^(a[176] & b[168])^(a[175] & b[169])^(a[174] & b[170])^(a[173] & b[171])^(a[172] & b[172])^(a[171] & b[173])^(a[170] & b[174])^(a[169] & b[175])^(a[168] & b[176])^(a[167] & b[177])^(a[166] & b[178])^(a[165] & b[179])^(a[164] & b[180])^(a[163] & b[181])^(a[162] & b[182])^(a[161] & b[183])^(a[160] & b[184])^(a[159] & b[185])^(a[158] & b[186])^(a[157] & b[187])^(a[156] & b[188])^(a[155] & b[189])^(a[154] & b[190])^(a[153] & b[191])^(a[152] & b[192])^(a[151] & b[193])^(a[150] & b[194])^(a[149] & b[195])^(a[148] & b[196])^(a[147] & b[197])^(a[146] & b[198])^(a[145] & b[199])^(a[144] & b[200])^(a[143] & b[201])^(a[142] & b[202])^(a[141] & b[203])^(a[140] & b[204])^(a[139] & b[205])^(a[138] & b[206])^(a[137] & b[207])^(a[136] & b[208])^(a[135] & b[209])^(a[134] & b[210])^(a[133] & b[211])^(a[132] & b[212])^(a[131] & b[213])^(a[130] & b[214])^(a[129] & b[215])^(a[128] & b[216])^(a[127] & b[217])^(a[126] & b[218])^(a[125] & b[219])^(a[124] & b[220])^(a[123] & b[221])^(a[122] & b[222])^(a[121] & b[223])^(a[120] & b[224])^(a[119] & b[225])^(a[118] & b[226])^(a[117] & b[227])^(a[116] & b[228])^(a[115] & b[229])^(a[114] & b[230])^(a[113] & b[231])^(a[112] & b[232])^(a[111] & b[233])^(a[110] & b[234])^(a[109] & b[235])^(a[108] & b[236])^(a[107] & b[237])^(a[106] & b[238])^(a[105] & b[239])^(a[104] & b[240])^(a[103] & b[241])^(a[102] & b[242])^(a[101] & b[243])^(a[100] & b[244])^(a[99] & b[245])^(a[98] & b[246])^(a[97] & b[247])^(a[96] & b[248])^(a[95] & b[249])^(a[94] & b[250])^(a[93] & b[251])^(a[92] & b[252])^(a[91] & b[253])^(a[90] & b[254])^(a[89] & b[255])^(a[88] & b[256])^(a[87] & b[257])^(a[86] & b[258])^(a[85] & b[259])^(a[84] & b[260])^(a[83] & b[261])^(a[82] & b[262])^(a[81] & b[263])^(a[80] & b[264])^(a[79] & b[265])^(a[78] & b[266])^(a[77] & b[267])^(a[76] & b[268])^(a[75] & b[269])^(a[74] & b[270])^(a[73] & b[271])^(a[72] & b[272])^(a[71] & b[273])^(a[70] & b[274])^(a[69] & b[275])^(a[68] & b[276])^(a[67] & b[277])^(a[66] & b[278])^(a[65] & b[279])^(a[64] & b[280])^(a[63] & b[281])^(a[62] & b[282])^(a[61] & b[283])^(a[60] & b[284])^(a[59] & b[285])^(a[58] & b[286])^(a[57] & b[287])^(a[56] & b[288])^(a[55] & b[289])^(a[54] & b[290])^(a[53] & b[291])^(a[52] & b[292])^(a[51] & b[293])^(a[50] & b[294])^(a[49] & b[295])^(a[48] & b[296])^(a[47] & b[297])^(a[46] & b[298])^(a[45] & b[299])^(a[44] & b[300])^(a[43] & b[301])^(a[42] & b[302])^(a[41] & b[303])^(a[40] & b[304])^(a[39] & b[305])^(a[38] & b[306])^(a[37] & b[307])^(a[36] & b[308])^(a[35] & b[309])^(a[34] & b[310])^(a[33] & b[311])^(a[32] & b[312])^(a[31] & b[313])^(a[30] & b[314])^(a[29] & b[315])^(a[28] & b[316])^(a[27] & b[317])^(a[26] & b[318])^(a[25] & b[319])^(a[24] & b[320])^(a[23] & b[321])^(a[22] & b[322])^(a[21] & b[323])^(a[20] & b[324])^(a[19] & b[325])^(a[18] & b[326])^(a[17] & b[327])^(a[16] & b[328])^(a[15] & b[329])^(a[14] & b[330])^(a[13] & b[331])^(a[12] & b[332])^(a[11] & b[333])^(a[10] & b[334])^(a[9] & b[335])^(a[8] & b[336])^(a[7] & b[337])^(a[6] & b[338])^(a[5] & b[339])^(a[4] & b[340])^(a[3] & b[341])^(a[2] & b[342])^(a[1] & b[343])^(a[0] & b[344]);
assign y[345] = (a[345] & b[0])^(a[344] & b[1])^(a[343] & b[2])^(a[342] & b[3])^(a[341] & b[4])^(a[340] & b[5])^(a[339] & b[6])^(a[338] & b[7])^(a[337] & b[8])^(a[336] & b[9])^(a[335] & b[10])^(a[334] & b[11])^(a[333] & b[12])^(a[332] & b[13])^(a[331] & b[14])^(a[330] & b[15])^(a[329] & b[16])^(a[328] & b[17])^(a[327] & b[18])^(a[326] & b[19])^(a[325] & b[20])^(a[324] & b[21])^(a[323] & b[22])^(a[322] & b[23])^(a[321] & b[24])^(a[320] & b[25])^(a[319] & b[26])^(a[318] & b[27])^(a[317] & b[28])^(a[316] & b[29])^(a[315] & b[30])^(a[314] & b[31])^(a[313] & b[32])^(a[312] & b[33])^(a[311] & b[34])^(a[310] & b[35])^(a[309] & b[36])^(a[308] & b[37])^(a[307] & b[38])^(a[306] & b[39])^(a[305] & b[40])^(a[304] & b[41])^(a[303] & b[42])^(a[302] & b[43])^(a[301] & b[44])^(a[300] & b[45])^(a[299] & b[46])^(a[298] & b[47])^(a[297] & b[48])^(a[296] & b[49])^(a[295] & b[50])^(a[294] & b[51])^(a[293] & b[52])^(a[292] & b[53])^(a[291] & b[54])^(a[290] & b[55])^(a[289] & b[56])^(a[288] & b[57])^(a[287] & b[58])^(a[286] & b[59])^(a[285] & b[60])^(a[284] & b[61])^(a[283] & b[62])^(a[282] & b[63])^(a[281] & b[64])^(a[280] & b[65])^(a[279] & b[66])^(a[278] & b[67])^(a[277] & b[68])^(a[276] & b[69])^(a[275] & b[70])^(a[274] & b[71])^(a[273] & b[72])^(a[272] & b[73])^(a[271] & b[74])^(a[270] & b[75])^(a[269] & b[76])^(a[268] & b[77])^(a[267] & b[78])^(a[266] & b[79])^(a[265] & b[80])^(a[264] & b[81])^(a[263] & b[82])^(a[262] & b[83])^(a[261] & b[84])^(a[260] & b[85])^(a[259] & b[86])^(a[258] & b[87])^(a[257] & b[88])^(a[256] & b[89])^(a[255] & b[90])^(a[254] & b[91])^(a[253] & b[92])^(a[252] & b[93])^(a[251] & b[94])^(a[250] & b[95])^(a[249] & b[96])^(a[248] & b[97])^(a[247] & b[98])^(a[246] & b[99])^(a[245] & b[100])^(a[244] & b[101])^(a[243] & b[102])^(a[242] & b[103])^(a[241] & b[104])^(a[240] & b[105])^(a[239] & b[106])^(a[238] & b[107])^(a[237] & b[108])^(a[236] & b[109])^(a[235] & b[110])^(a[234] & b[111])^(a[233] & b[112])^(a[232] & b[113])^(a[231] & b[114])^(a[230] & b[115])^(a[229] & b[116])^(a[228] & b[117])^(a[227] & b[118])^(a[226] & b[119])^(a[225] & b[120])^(a[224] & b[121])^(a[223] & b[122])^(a[222] & b[123])^(a[221] & b[124])^(a[220] & b[125])^(a[219] & b[126])^(a[218] & b[127])^(a[217] & b[128])^(a[216] & b[129])^(a[215] & b[130])^(a[214] & b[131])^(a[213] & b[132])^(a[212] & b[133])^(a[211] & b[134])^(a[210] & b[135])^(a[209] & b[136])^(a[208] & b[137])^(a[207] & b[138])^(a[206] & b[139])^(a[205] & b[140])^(a[204] & b[141])^(a[203] & b[142])^(a[202] & b[143])^(a[201] & b[144])^(a[200] & b[145])^(a[199] & b[146])^(a[198] & b[147])^(a[197] & b[148])^(a[196] & b[149])^(a[195] & b[150])^(a[194] & b[151])^(a[193] & b[152])^(a[192] & b[153])^(a[191] & b[154])^(a[190] & b[155])^(a[189] & b[156])^(a[188] & b[157])^(a[187] & b[158])^(a[186] & b[159])^(a[185] & b[160])^(a[184] & b[161])^(a[183] & b[162])^(a[182] & b[163])^(a[181] & b[164])^(a[180] & b[165])^(a[179] & b[166])^(a[178] & b[167])^(a[177] & b[168])^(a[176] & b[169])^(a[175] & b[170])^(a[174] & b[171])^(a[173] & b[172])^(a[172] & b[173])^(a[171] & b[174])^(a[170] & b[175])^(a[169] & b[176])^(a[168] & b[177])^(a[167] & b[178])^(a[166] & b[179])^(a[165] & b[180])^(a[164] & b[181])^(a[163] & b[182])^(a[162] & b[183])^(a[161] & b[184])^(a[160] & b[185])^(a[159] & b[186])^(a[158] & b[187])^(a[157] & b[188])^(a[156] & b[189])^(a[155] & b[190])^(a[154] & b[191])^(a[153] & b[192])^(a[152] & b[193])^(a[151] & b[194])^(a[150] & b[195])^(a[149] & b[196])^(a[148] & b[197])^(a[147] & b[198])^(a[146] & b[199])^(a[145] & b[200])^(a[144] & b[201])^(a[143] & b[202])^(a[142] & b[203])^(a[141] & b[204])^(a[140] & b[205])^(a[139] & b[206])^(a[138] & b[207])^(a[137] & b[208])^(a[136] & b[209])^(a[135] & b[210])^(a[134] & b[211])^(a[133] & b[212])^(a[132] & b[213])^(a[131] & b[214])^(a[130] & b[215])^(a[129] & b[216])^(a[128] & b[217])^(a[127] & b[218])^(a[126] & b[219])^(a[125] & b[220])^(a[124] & b[221])^(a[123] & b[222])^(a[122] & b[223])^(a[121] & b[224])^(a[120] & b[225])^(a[119] & b[226])^(a[118] & b[227])^(a[117] & b[228])^(a[116] & b[229])^(a[115] & b[230])^(a[114] & b[231])^(a[113] & b[232])^(a[112] & b[233])^(a[111] & b[234])^(a[110] & b[235])^(a[109] & b[236])^(a[108] & b[237])^(a[107] & b[238])^(a[106] & b[239])^(a[105] & b[240])^(a[104] & b[241])^(a[103] & b[242])^(a[102] & b[243])^(a[101] & b[244])^(a[100] & b[245])^(a[99] & b[246])^(a[98] & b[247])^(a[97] & b[248])^(a[96] & b[249])^(a[95] & b[250])^(a[94] & b[251])^(a[93] & b[252])^(a[92] & b[253])^(a[91] & b[254])^(a[90] & b[255])^(a[89] & b[256])^(a[88] & b[257])^(a[87] & b[258])^(a[86] & b[259])^(a[85] & b[260])^(a[84] & b[261])^(a[83] & b[262])^(a[82] & b[263])^(a[81] & b[264])^(a[80] & b[265])^(a[79] & b[266])^(a[78] & b[267])^(a[77] & b[268])^(a[76] & b[269])^(a[75] & b[270])^(a[74] & b[271])^(a[73] & b[272])^(a[72] & b[273])^(a[71] & b[274])^(a[70] & b[275])^(a[69] & b[276])^(a[68] & b[277])^(a[67] & b[278])^(a[66] & b[279])^(a[65] & b[280])^(a[64] & b[281])^(a[63] & b[282])^(a[62] & b[283])^(a[61] & b[284])^(a[60] & b[285])^(a[59] & b[286])^(a[58] & b[287])^(a[57] & b[288])^(a[56] & b[289])^(a[55] & b[290])^(a[54] & b[291])^(a[53] & b[292])^(a[52] & b[293])^(a[51] & b[294])^(a[50] & b[295])^(a[49] & b[296])^(a[48] & b[297])^(a[47] & b[298])^(a[46] & b[299])^(a[45] & b[300])^(a[44] & b[301])^(a[43] & b[302])^(a[42] & b[303])^(a[41] & b[304])^(a[40] & b[305])^(a[39] & b[306])^(a[38] & b[307])^(a[37] & b[308])^(a[36] & b[309])^(a[35] & b[310])^(a[34] & b[311])^(a[33] & b[312])^(a[32] & b[313])^(a[31] & b[314])^(a[30] & b[315])^(a[29] & b[316])^(a[28] & b[317])^(a[27] & b[318])^(a[26] & b[319])^(a[25] & b[320])^(a[24] & b[321])^(a[23] & b[322])^(a[22] & b[323])^(a[21] & b[324])^(a[20] & b[325])^(a[19] & b[326])^(a[18] & b[327])^(a[17] & b[328])^(a[16] & b[329])^(a[15] & b[330])^(a[14] & b[331])^(a[13] & b[332])^(a[12] & b[333])^(a[11] & b[334])^(a[10] & b[335])^(a[9] & b[336])^(a[8] & b[337])^(a[7] & b[338])^(a[6] & b[339])^(a[5] & b[340])^(a[4] & b[341])^(a[3] & b[342])^(a[2] & b[343])^(a[1] & b[344])^(a[0] & b[345]);
assign y[346] = (a[346] & b[0])^(a[345] & b[1])^(a[344] & b[2])^(a[343] & b[3])^(a[342] & b[4])^(a[341] & b[5])^(a[340] & b[6])^(a[339] & b[7])^(a[338] & b[8])^(a[337] & b[9])^(a[336] & b[10])^(a[335] & b[11])^(a[334] & b[12])^(a[333] & b[13])^(a[332] & b[14])^(a[331] & b[15])^(a[330] & b[16])^(a[329] & b[17])^(a[328] & b[18])^(a[327] & b[19])^(a[326] & b[20])^(a[325] & b[21])^(a[324] & b[22])^(a[323] & b[23])^(a[322] & b[24])^(a[321] & b[25])^(a[320] & b[26])^(a[319] & b[27])^(a[318] & b[28])^(a[317] & b[29])^(a[316] & b[30])^(a[315] & b[31])^(a[314] & b[32])^(a[313] & b[33])^(a[312] & b[34])^(a[311] & b[35])^(a[310] & b[36])^(a[309] & b[37])^(a[308] & b[38])^(a[307] & b[39])^(a[306] & b[40])^(a[305] & b[41])^(a[304] & b[42])^(a[303] & b[43])^(a[302] & b[44])^(a[301] & b[45])^(a[300] & b[46])^(a[299] & b[47])^(a[298] & b[48])^(a[297] & b[49])^(a[296] & b[50])^(a[295] & b[51])^(a[294] & b[52])^(a[293] & b[53])^(a[292] & b[54])^(a[291] & b[55])^(a[290] & b[56])^(a[289] & b[57])^(a[288] & b[58])^(a[287] & b[59])^(a[286] & b[60])^(a[285] & b[61])^(a[284] & b[62])^(a[283] & b[63])^(a[282] & b[64])^(a[281] & b[65])^(a[280] & b[66])^(a[279] & b[67])^(a[278] & b[68])^(a[277] & b[69])^(a[276] & b[70])^(a[275] & b[71])^(a[274] & b[72])^(a[273] & b[73])^(a[272] & b[74])^(a[271] & b[75])^(a[270] & b[76])^(a[269] & b[77])^(a[268] & b[78])^(a[267] & b[79])^(a[266] & b[80])^(a[265] & b[81])^(a[264] & b[82])^(a[263] & b[83])^(a[262] & b[84])^(a[261] & b[85])^(a[260] & b[86])^(a[259] & b[87])^(a[258] & b[88])^(a[257] & b[89])^(a[256] & b[90])^(a[255] & b[91])^(a[254] & b[92])^(a[253] & b[93])^(a[252] & b[94])^(a[251] & b[95])^(a[250] & b[96])^(a[249] & b[97])^(a[248] & b[98])^(a[247] & b[99])^(a[246] & b[100])^(a[245] & b[101])^(a[244] & b[102])^(a[243] & b[103])^(a[242] & b[104])^(a[241] & b[105])^(a[240] & b[106])^(a[239] & b[107])^(a[238] & b[108])^(a[237] & b[109])^(a[236] & b[110])^(a[235] & b[111])^(a[234] & b[112])^(a[233] & b[113])^(a[232] & b[114])^(a[231] & b[115])^(a[230] & b[116])^(a[229] & b[117])^(a[228] & b[118])^(a[227] & b[119])^(a[226] & b[120])^(a[225] & b[121])^(a[224] & b[122])^(a[223] & b[123])^(a[222] & b[124])^(a[221] & b[125])^(a[220] & b[126])^(a[219] & b[127])^(a[218] & b[128])^(a[217] & b[129])^(a[216] & b[130])^(a[215] & b[131])^(a[214] & b[132])^(a[213] & b[133])^(a[212] & b[134])^(a[211] & b[135])^(a[210] & b[136])^(a[209] & b[137])^(a[208] & b[138])^(a[207] & b[139])^(a[206] & b[140])^(a[205] & b[141])^(a[204] & b[142])^(a[203] & b[143])^(a[202] & b[144])^(a[201] & b[145])^(a[200] & b[146])^(a[199] & b[147])^(a[198] & b[148])^(a[197] & b[149])^(a[196] & b[150])^(a[195] & b[151])^(a[194] & b[152])^(a[193] & b[153])^(a[192] & b[154])^(a[191] & b[155])^(a[190] & b[156])^(a[189] & b[157])^(a[188] & b[158])^(a[187] & b[159])^(a[186] & b[160])^(a[185] & b[161])^(a[184] & b[162])^(a[183] & b[163])^(a[182] & b[164])^(a[181] & b[165])^(a[180] & b[166])^(a[179] & b[167])^(a[178] & b[168])^(a[177] & b[169])^(a[176] & b[170])^(a[175] & b[171])^(a[174] & b[172])^(a[173] & b[173])^(a[172] & b[174])^(a[171] & b[175])^(a[170] & b[176])^(a[169] & b[177])^(a[168] & b[178])^(a[167] & b[179])^(a[166] & b[180])^(a[165] & b[181])^(a[164] & b[182])^(a[163] & b[183])^(a[162] & b[184])^(a[161] & b[185])^(a[160] & b[186])^(a[159] & b[187])^(a[158] & b[188])^(a[157] & b[189])^(a[156] & b[190])^(a[155] & b[191])^(a[154] & b[192])^(a[153] & b[193])^(a[152] & b[194])^(a[151] & b[195])^(a[150] & b[196])^(a[149] & b[197])^(a[148] & b[198])^(a[147] & b[199])^(a[146] & b[200])^(a[145] & b[201])^(a[144] & b[202])^(a[143] & b[203])^(a[142] & b[204])^(a[141] & b[205])^(a[140] & b[206])^(a[139] & b[207])^(a[138] & b[208])^(a[137] & b[209])^(a[136] & b[210])^(a[135] & b[211])^(a[134] & b[212])^(a[133] & b[213])^(a[132] & b[214])^(a[131] & b[215])^(a[130] & b[216])^(a[129] & b[217])^(a[128] & b[218])^(a[127] & b[219])^(a[126] & b[220])^(a[125] & b[221])^(a[124] & b[222])^(a[123] & b[223])^(a[122] & b[224])^(a[121] & b[225])^(a[120] & b[226])^(a[119] & b[227])^(a[118] & b[228])^(a[117] & b[229])^(a[116] & b[230])^(a[115] & b[231])^(a[114] & b[232])^(a[113] & b[233])^(a[112] & b[234])^(a[111] & b[235])^(a[110] & b[236])^(a[109] & b[237])^(a[108] & b[238])^(a[107] & b[239])^(a[106] & b[240])^(a[105] & b[241])^(a[104] & b[242])^(a[103] & b[243])^(a[102] & b[244])^(a[101] & b[245])^(a[100] & b[246])^(a[99] & b[247])^(a[98] & b[248])^(a[97] & b[249])^(a[96] & b[250])^(a[95] & b[251])^(a[94] & b[252])^(a[93] & b[253])^(a[92] & b[254])^(a[91] & b[255])^(a[90] & b[256])^(a[89] & b[257])^(a[88] & b[258])^(a[87] & b[259])^(a[86] & b[260])^(a[85] & b[261])^(a[84] & b[262])^(a[83] & b[263])^(a[82] & b[264])^(a[81] & b[265])^(a[80] & b[266])^(a[79] & b[267])^(a[78] & b[268])^(a[77] & b[269])^(a[76] & b[270])^(a[75] & b[271])^(a[74] & b[272])^(a[73] & b[273])^(a[72] & b[274])^(a[71] & b[275])^(a[70] & b[276])^(a[69] & b[277])^(a[68] & b[278])^(a[67] & b[279])^(a[66] & b[280])^(a[65] & b[281])^(a[64] & b[282])^(a[63] & b[283])^(a[62] & b[284])^(a[61] & b[285])^(a[60] & b[286])^(a[59] & b[287])^(a[58] & b[288])^(a[57] & b[289])^(a[56] & b[290])^(a[55] & b[291])^(a[54] & b[292])^(a[53] & b[293])^(a[52] & b[294])^(a[51] & b[295])^(a[50] & b[296])^(a[49] & b[297])^(a[48] & b[298])^(a[47] & b[299])^(a[46] & b[300])^(a[45] & b[301])^(a[44] & b[302])^(a[43] & b[303])^(a[42] & b[304])^(a[41] & b[305])^(a[40] & b[306])^(a[39] & b[307])^(a[38] & b[308])^(a[37] & b[309])^(a[36] & b[310])^(a[35] & b[311])^(a[34] & b[312])^(a[33] & b[313])^(a[32] & b[314])^(a[31] & b[315])^(a[30] & b[316])^(a[29] & b[317])^(a[28] & b[318])^(a[27] & b[319])^(a[26] & b[320])^(a[25] & b[321])^(a[24] & b[322])^(a[23] & b[323])^(a[22] & b[324])^(a[21] & b[325])^(a[20] & b[326])^(a[19] & b[327])^(a[18] & b[328])^(a[17] & b[329])^(a[16] & b[330])^(a[15] & b[331])^(a[14] & b[332])^(a[13] & b[333])^(a[12] & b[334])^(a[11] & b[335])^(a[10] & b[336])^(a[9] & b[337])^(a[8] & b[338])^(a[7] & b[339])^(a[6] & b[340])^(a[5] & b[341])^(a[4] & b[342])^(a[3] & b[343])^(a[2] & b[344])^(a[1] & b[345])^(a[0] & b[346]);
assign y[347] = (a[347] & b[0])^(a[346] & b[1])^(a[345] & b[2])^(a[344] & b[3])^(a[343] & b[4])^(a[342] & b[5])^(a[341] & b[6])^(a[340] & b[7])^(a[339] & b[8])^(a[338] & b[9])^(a[337] & b[10])^(a[336] & b[11])^(a[335] & b[12])^(a[334] & b[13])^(a[333] & b[14])^(a[332] & b[15])^(a[331] & b[16])^(a[330] & b[17])^(a[329] & b[18])^(a[328] & b[19])^(a[327] & b[20])^(a[326] & b[21])^(a[325] & b[22])^(a[324] & b[23])^(a[323] & b[24])^(a[322] & b[25])^(a[321] & b[26])^(a[320] & b[27])^(a[319] & b[28])^(a[318] & b[29])^(a[317] & b[30])^(a[316] & b[31])^(a[315] & b[32])^(a[314] & b[33])^(a[313] & b[34])^(a[312] & b[35])^(a[311] & b[36])^(a[310] & b[37])^(a[309] & b[38])^(a[308] & b[39])^(a[307] & b[40])^(a[306] & b[41])^(a[305] & b[42])^(a[304] & b[43])^(a[303] & b[44])^(a[302] & b[45])^(a[301] & b[46])^(a[300] & b[47])^(a[299] & b[48])^(a[298] & b[49])^(a[297] & b[50])^(a[296] & b[51])^(a[295] & b[52])^(a[294] & b[53])^(a[293] & b[54])^(a[292] & b[55])^(a[291] & b[56])^(a[290] & b[57])^(a[289] & b[58])^(a[288] & b[59])^(a[287] & b[60])^(a[286] & b[61])^(a[285] & b[62])^(a[284] & b[63])^(a[283] & b[64])^(a[282] & b[65])^(a[281] & b[66])^(a[280] & b[67])^(a[279] & b[68])^(a[278] & b[69])^(a[277] & b[70])^(a[276] & b[71])^(a[275] & b[72])^(a[274] & b[73])^(a[273] & b[74])^(a[272] & b[75])^(a[271] & b[76])^(a[270] & b[77])^(a[269] & b[78])^(a[268] & b[79])^(a[267] & b[80])^(a[266] & b[81])^(a[265] & b[82])^(a[264] & b[83])^(a[263] & b[84])^(a[262] & b[85])^(a[261] & b[86])^(a[260] & b[87])^(a[259] & b[88])^(a[258] & b[89])^(a[257] & b[90])^(a[256] & b[91])^(a[255] & b[92])^(a[254] & b[93])^(a[253] & b[94])^(a[252] & b[95])^(a[251] & b[96])^(a[250] & b[97])^(a[249] & b[98])^(a[248] & b[99])^(a[247] & b[100])^(a[246] & b[101])^(a[245] & b[102])^(a[244] & b[103])^(a[243] & b[104])^(a[242] & b[105])^(a[241] & b[106])^(a[240] & b[107])^(a[239] & b[108])^(a[238] & b[109])^(a[237] & b[110])^(a[236] & b[111])^(a[235] & b[112])^(a[234] & b[113])^(a[233] & b[114])^(a[232] & b[115])^(a[231] & b[116])^(a[230] & b[117])^(a[229] & b[118])^(a[228] & b[119])^(a[227] & b[120])^(a[226] & b[121])^(a[225] & b[122])^(a[224] & b[123])^(a[223] & b[124])^(a[222] & b[125])^(a[221] & b[126])^(a[220] & b[127])^(a[219] & b[128])^(a[218] & b[129])^(a[217] & b[130])^(a[216] & b[131])^(a[215] & b[132])^(a[214] & b[133])^(a[213] & b[134])^(a[212] & b[135])^(a[211] & b[136])^(a[210] & b[137])^(a[209] & b[138])^(a[208] & b[139])^(a[207] & b[140])^(a[206] & b[141])^(a[205] & b[142])^(a[204] & b[143])^(a[203] & b[144])^(a[202] & b[145])^(a[201] & b[146])^(a[200] & b[147])^(a[199] & b[148])^(a[198] & b[149])^(a[197] & b[150])^(a[196] & b[151])^(a[195] & b[152])^(a[194] & b[153])^(a[193] & b[154])^(a[192] & b[155])^(a[191] & b[156])^(a[190] & b[157])^(a[189] & b[158])^(a[188] & b[159])^(a[187] & b[160])^(a[186] & b[161])^(a[185] & b[162])^(a[184] & b[163])^(a[183] & b[164])^(a[182] & b[165])^(a[181] & b[166])^(a[180] & b[167])^(a[179] & b[168])^(a[178] & b[169])^(a[177] & b[170])^(a[176] & b[171])^(a[175] & b[172])^(a[174] & b[173])^(a[173] & b[174])^(a[172] & b[175])^(a[171] & b[176])^(a[170] & b[177])^(a[169] & b[178])^(a[168] & b[179])^(a[167] & b[180])^(a[166] & b[181])^(a[165] & b[182])^(a[164] & b[183])^(a[163] & b[184])^(a[162] & b[185])^(a[161] & b[186])^(a[160] & b[187])^(a[159] & b[188])^(a[158] & b[189])^(a[157] & b[190])^(a[156] & b[191])^(a[155] & b[192])^(a[154] & b[193])^(a[153] & b[194])^(a[152] & b[195])^(a[151] & b[196])^(a[150] & b[197])^(a[149] & b[198])^(a[148] & b[199])^(a[147] & b[200])^(a[146] & b[201])^(a[145] & b[202])^(a[144] & b[203])^(a[143] & b[204])^(a[142] & b[205])^(a[141] & b[206])^(a[140] & b[207])^(a[139] & b[208])^(a[138] & b[209])^(a[137] & b[210])^(a[136] & b[211])^(a[135] & b[212])^(a[134] & b[213])^(a[133] & b[214])^(a[132] & b[215])^(a[131] & b[216])^(a[130] & b[217])^(a[129] & b[218])^(a[128] & b[219])^(a[127] & b[220])^(a[126] & b[221])^(a[125] & b[222])^(a[124] & b[223])^(a[123] & b[224])^(a[122] & b[225])^(a[121] & b[226])^(a[120] & b[227])^(a[119] & b[228])^(a[118] & b[229])^(a[117] & b[230])^(a[116] & b[231])^(a[115] & b[232])^(a[114] & b[233])^(a[113] & b[234])^(a[112] & b[235])^(a[111] & b[236])^(a[110] & b[237])^(a[109] & b[238])^(a[108] & b[239])^(a[107] & b[240])^(a[106] & b[241])^(a[105] & b[242])^(a[104] & b[243])^(a[103] & b[244])^(a[102] & b[245])^(a[101] & b[246])^(a[100] & b[247])^(a[99] & b[248])^(a[98] & b[249])^(a[97] & b[250])^(a[96] & b[251])^(a[95] & b[252])^(a[94] & b[253])^(a[93] & b[254])^(a[92] & b[255])^(a[91] & b[256])^(a[90] & b[257])^(a[89] & b[258])^(a[88] & b[259])^(a[87] & b[260])^(a[86] & b[261])^(a[85] & b[262])^(a[84] & b[263])^(a[83] & b[264])^(a[82] & b[265])^(a[81] & b[266])^(a[80] & b[267])^(a[79] & b[268])^(a[78] & b[269])^(a[77] & b[270])^(a[76] & b[271])^(a[75] & b[272])^(a[74] & b[273])^(a[73] & b[274])^(a[72] & b[275])^(a[71] & b[276])^(a[70] & b[277])^(a[69] & b[278])^(a[68] & b[279])^(a[67] & b[280])^(a[66] & b[281])^(a[65] & b[282])^(a[64] & b[283])^(a[63] & b[284])^(a[62] & b[285])^(a[61] & b[286])^(a[60] & b[287])^(a[59] & b[288])^(a[58] & b[289])^(a[57] & b[290])^(a[56] & b[291])^(a[55] & b[292])^(a[54] & b[293])^(a[53] & b[294])^(a[52] & b[295])^(a[51] & b[296])^(a[50] & b[297])^(a[49] & b[298])^(a[48] & b[299])^(a[47] & b[300])^(a[46] & b[301])^(a[45] & b[302])^(a[44] & b[303])^(a[43] & b[304])^(a[42] & b[305])^(a[41] & b[306])^(a[40] & b[307])^(a[39] & b[308])^(a[38] & b[309])^(a[37] & b[310])^(a[36] & b[311])^(a[35] & b[312])^(a[34] & b[313])^(a[33] & b[314])^(a[32] & b[315])^(a[31] & b[316])^(a[30] & b[317])^(a[29] & b[318])^(a[28] & b[319])^(a[27] & b[320])^(a[26] & b[321])^(a[25] & b[322])^(a[24] & b[323])^(a[23] & b[324])^(a[22] & b[325])^(a[21] & b[326])^(a[20] & b[327])^(a[19] & b[328])^(a[18] & b[329])^(a[17] & b[330])^(a[16] & b[331])^(a[15] & b[332])^(a[14] & b[333])^(a[13] & b[334])^(a[12] & b[335])^(a[11] & b[336])^(a[10] & b[337])^(a[9] & b[338])^(a[8] & b[339])^(a[7] & b[340])^(a[6] & b[341])^(a[5] & b[342])^(a[4] & b[343])^(a[3] & b[344])^(a[2] & b[345])^(a[1] & b[346])^(a[0] & b[347]);
assign y[348] = (a[348] & b[0])^(a[347] & b[1])^(a[346] & b[2])^(a[345] & b[3])^(a[344] & b[4])^(a[343] & b[5])^(a[342] & b[6])^(a[341] & b[7])^(a[340] & b[8])^(a[339] & b[9])^(a[338] & b[10])^(a[337] & b[11])^(a[336] & b[12])^(a[335] & b[13])^(a[334] & b[14])^(a[333] & b[15])^(a[332] & b[16])^(a[331] & b[17])^(a[330] & b[18])^(a[329] & b[19])^(a[328] & b[20])^(a[327] & b[21])^(a[326] & b[22])^(a[325] & b[23])^(a[324] & b[24])^(a[323] & b[25])^(a[322] & b[26])^(a[321] & b[27])^(a[320] & b[28])^(a[319] & b[29])^(a[318] & b[30])^(a[317] & b[31])^(a[316] & b[32])^(a[315] & b[33])^(a[314] & b[34])^(a[313] & b[35])^(a[312] & b[36])^(a[311] & b[37])^(a[310] & b[38])^(a[309] & b[39])^(a[308] & b[40])^(a[307] & b[41])^(a[306] & b[42])^(a[305] & b[43])^(a[304] & b[44])^(a[303] & b[45])^(a[302] & b[46])^(a[301] & b[47])^(a[300] & b[48])^(a[299] & b[49])^(a[298] & b[50])^(a[297] & b[51])^(a[296] & b[52])^(a[295] & b[53])^(a[294] & b[54])^(a[293] & b[55])^(a[292] & b[56])^(a[291] & b[57])^(a[290] & b[58])^(a[289] & b[59])^(a[288] & b[60])^(a[287] & b[61])^(a[286] & b[62])^(a[285] & b[63])^(a[284] & b[64])^(a[283] & b[65])^(a[282] & b[66])^(a[281] & b[67])^(a[280] & b[68])^(a[279] & b[69])^(a[278] & b[70])^(a[277] & b[71])^(a[276] & b[72])^(a[275] & b[73])^(a[274] & b[74])^(a[273] & b[75])^(a[272] & b[76])^(a[271] & b[77])^(a[270] & b[78])^(a[269] & b[79])^(a[268] & b[80])^(a[267] & b[81])^(a[266] & b[82])^(a[265] & b[83])^(a[264] & b[84])^(a[263] & b[85])^(a[262] & b[86])^(a[261] & b[87])^(a[260] & b[88])^(a[259] & b[89])^(a[258] & b[90])^(a[257] & b[91])^(a[256] & b[92])^(a[255] & b[93])^(a[254] & b[94])^(a[253] & b[95])^(a[252] & b[96])^(a[251] & b[97])^(a[250] & b[98])^(a[249] & b[99])^(a[248] & b[100])^(a[247] & b[101])^(a[246] & b[102])^(a[245] & b[103])^(a[244] & b[104])^(a[243] & b[105])^(a[242] & b[106])^(a[241] & b[107])^(a[240] & b[108])^(a[239] & b[109])^(a[238] & b[110])^(a[237] & b[111])^(a[236] & b[112])^(a[235] & b[113])^(a[234] & b[114])^(a[233] & b[115])^(a[232] & b[116])^(a[231] & b[117])^(a[230] & b[118])^(a[229] & b[119])^(a[228] & b[120])^(a[227] & b[121])^(a[226] & b[122])^(a[225] & b[123])^(a[224] & b[124])^(a[223] & b[125])^(a[222] & b[126])^(a[221] & b[127])^(a[220] & b[128])^(a[219] & b[129])^(a[218] & b[130])^(a[217] & b[131])^(a[216] & b[132])^(a[215] & b[133])^(a[214] & b[134])^(a[213] & b[135])^(a[212] & b[136])^(a[211] & b[137])^(a[210] & b[138])^(a[209] & b[139])^(a[208] & b[140])^(a[207] & b[141])^(a[206] & b[142])^(a[205] & b[143])^(a[204] & b[144])^(a[203] & b[145])^(a[202] & b[146])^(a[201] & b[147])^(a[200] & b[148])^(a[199] & b[149])^(a[198] & b[150])^(a[197] & b[151])^(a[196] & b[152])^(a[195] & b[153])^(a[194] & b[154])^(a[193] & b[155])^(a[192] & b[156])^(a[191] & b[157])^(a[190] & b[158])^(a[189] & b[159])^(a[188] & b[160])^(a[187] & b[161])^(a[186] & b[162])^(a[185] & b[163])^(a[184] & b[164])^(a[183] & b[165])^(a[182] & b[166])^(a[181] & b[167])^(a[180] & b[168])^(a[179] & b[169])^(a[178] & b[170])^(a[177] & b[171])^(a[176] & b[172])^(a[175] & b[173])^(a[174] & b[174])^(a[173] & b[175])^(a[172] & b[176])^(a[171] & b[177])^(a[170] & b[178])^(a[169] & b[179])^(a[168] & b[180])^(a[167] & b[181])^(a[166] & b[182])^(a[165] & b[183])^(a[164] & b[184])^(a[163] & b[185])^(a[162] & b[186])^(a[161] & b[187])^(a[160] & b[188])^(a[159] & b[189])^(a[158] & b[190])^(a[157] & b[191])^(a[156] & b[192])^(a[155] & b[193])^(a[154] & b[194])^(a[153] & b[195])^(a[152] & b[196])^(a[151] & b[197])^(a[150] & b[198])^(a[149] & b[199])^(a[148] & b[200])^(a[147] & b[201])^(a[146] & b[202])^(a[145] & b[203])^(a[144] & b[204])^(a[143] & b[205])^(a[142] & b[206])^(a[141] & b[207])^(a[140] & b[208])^(a[139] & b[209])^(a[138] & b[210])^(a[137] & b[211])^(a[136] & b[212])^(a[135] & b[213])^(a[134] & b[214])^(a[133] & b[215])^(a[132] & b[216])^(a[131] & b[217])^(a[130] & b[218])^(a[129] & b[219])^(a[128] & b[220])^(a[127] & b[221])^(a[126] & b[222])^(a[125] & b[223])^(a[124] & b[224])^(a[123] & b[225])^(a[122] & b[226])^(a[121] & b[227])^(a[120] & b[228])^(a[119] & b[229])^(a[118] & b[230])^(a[117] & b[231])^(a[116] & b[232])^(a[115] & b[233])^(a[114] & b[234])^(a[113] & b[235])^(a[112] & b[236])^(a[111] & b[237])^(a[110] & b[238])^(a[109] & b[239])^(a[108] & b[240])^(a[107] & b[241])^(a[106] & b[242])^(a[105] & b[243])^(a[104] & b[244])^(a[103] & b[245])^(a[102] & b[246])^(a[101] & b[247])^(a[100] & b[248])^(a[99] & b[249])^(a[98] & b[250])^(a[97] & b[251])^(a[96] & b[252])^(a[95] & b[253])^(a[94] & b[254])^(a[93] & b[255])^(a[92] & b[256])^(a[91] & b[257])^(a[90] & b[258])^(a[89] & b[259])^(a[88] & b[260])^(a[87] & b[261])^(a[86] & b[262])^(a[85] & b[263])^(a[84] & b[264])^(a[83] & b[265])^(a[82] & b[266])^(a[81] & b[267])^(a[80] & b[268])^(a[79] & b[269])^(a[78] & b[270])^(a[77] & b[271])^(a[76] & b[272])^(a[75] & b[273])^(a[74] & b[274])^(a[73] & b[275])^(a[72] & b[276])^(a[71] & b[277])^(a[70] & b[278])^(a[69] & b[279])^(a[68] & b[280])^(a[67] & b[281])^(a[66] & b[282])^(a[65] & b[283])^(a[64] & b[284])^(a[63] & b[285])^(a[62] & b[286])^(a[61] & b[287])^(a[60] & b[288])^(a[59] & b[289])^(a[58] & b[290])^(a[57] & b[291])^(a[56] & b[292])^(a[55] & b[293])^(a[54] & b[294])^(a[53] & b[295])^(a[52] & b[296])^(a[51] & b[297])^(a[50] & b[298])^(a[49] & b[299])^(a[48] & b[300])^(a[47] & b[301])^(a[46] & b[302])^(a[45] & b[303])^(a[44] & b[304])^(a[43] & b[305])^(a[42] & b[306])^(a[41] & b[307])^(a[40] & b[308])^(a[39] & b[309])^(a[38] & b[310])^(a[37] & b[311])^(a[36] & b[312])^(a[35] & b[313])^(a[34] & b[314])^(a[33] & b[315])^(a[32] & b[316])^(a[31] & b[317])^(a[30] & b[318])^(a[29] & b[319])^(a[28] & b[320])^(a[27] & b[321])^(a[26] & b[322])^(a[25] & b[323])^(a[24] & b[324])^(a[23] & b[325])^(a[22] & b[326])^(a[21] & b[327])^(a[20] & b[328])^(a[19] & b[329])^(a[18] & b[330])^(a[17] & b[331])^(a[16] & b[332])^(a[15] & b[333])^(a[14] & b[334])^(a[13] & b[335])^(a[12] & b[336])^(a[11] & b[337])^(a[10] & b[338])^(a[9] & b[339])^(a[8] & b[340])^(a[7] & b[341])^(a[6] & b[342])^(a[5] & b[343])^(a[4] & b[344])^(a[3] & b[345])^(a[2] & b[346])^(a[1] & b[347])^(a[0] & b[348]);
assign y[349] = (a[349] & b[0])^(a[348] & b[1])^(a[347] & b[2])^(a[346] & b[3])^(a[345] & b[4])^(a[344] & b[5])^(a[343] & b[6])^(a[342] & b[7])^(a[341] & b[8])^(a[340] & b[9])^(a[339] & b[10])^(a[338] & b[11])^(a[337] & b[12])^(a[336] & b[13])^(a[335] & b[14])^(a[334] & b[15])^(a[333] & b[16])^(a[332] & b[17])^(a[331] & b[18])^(a[330] & b[19])^(a[329] & b[20])^(a[328] & b[21])^(a[327] & b[22])^(a[326] & b[23])^(a[325] & b[24])^(a[324] & b[25])^(a[323] & b[26])^(a[322] & b[27])^(a[321] & b[28])^(a[320] & b[29])^(a[319] & b[30])^(a[318] & b[31])^(a[317] & b[32])^(a[316] & b[33])^(a[315] & b[34])^(a[314] & b[35])^(a[313] & b[36])^(a[312] & b[37])^(a[311] & b[38])^(a[310] & b[39])^(a[309] & b[40])^(a[308] & b[41])^(a[307] & b[42])^(a[306] & b[43])^(a[305] & b[44])^(a[304] & b[45])^(a[303] & b[46])^(a[302] & b[47])^(a[301] & b[48])^(a[300] & b[49])^(a[299] & b[50])^(a[298] & b[51])^(a[297] & b[52])^(a[296] & b[53])^(a[295] & b[54])^(a[294] & b[55])^(a[293] & b[56])^(a[292] & b[57])^(a[291] & b[58])^(a[290] & b[59])^(a[289] & b[60])^(a[288] & b[61])^(a[287] & b[62])^(a[286] & b[63])^(a[285] & b[64])^(a[284] & b[65])^(a[283] & b[66])^(a[282] & b[67])^(a[281] & b[68])^(a[280] & b[69])^(a[279] & b[70])^(a[278] & b[71])^(a[277] & b[72])^(a[276] & b[73])^(a[275] & b[74])^(a[274] & b[75])^(a[273] & b[76])^(a[272] & b[77])^(a[271] & b[78])^(a[270] & b[79])^(a[269] & b[80])^(a[268] & b[81])^(a[267] & b[82])^(a[266] & b[83])^(a[265] & b[84])^(a[264] & b[85])^(a[263] & b[86])^(a[262] & b[87])^(a[261] & b[88])^(a[260] & b[89])^(a[259] & b[90])^(a[258] & b[91])^(a[257] & b[92])^(a[256] & b[93])^(a[255] & b[94])^(a[254] & b[95])^(a[253] & b[96])^(a[252] & b[97])^(a[251] & b[98])^(a[250] & b[99])^(a[249] & b[100])^(a[248] & b[101])^(a[247] & b[102])^(a[246] & b[103])^(a[245] & b[104])^(a[244] & b[105])^(a[243] & b[106])^(a[242] & b[107])^(a[241] & b[108])^(a[240] & b[109])^(a[239] & b[110])^(a[238] & b[111])^(a[237] & b[112])^(a[236] & b[113])^(a[235] & b[114])^(a[234] & b[115])^(a[233] & b[116])^(a[232] & b[117])^(a[231] & b[118])^(a[230] & b[119])^(a[229] & b[120])^(a[228] & b[121])^(a[227] & b[122])^(a[226] & b[123])^(a[225] & b[124])^(a[224] & b[125])^(a[223] & b[126])^(a[222] & b[127])^(a[221] & b[128])^(a[220] & b[129])^(a[219] & b[130])^(a[218] & b[131])^(a[217] & b[132])^(a[216] & b[133])^(a[215] & b[134])^(a[214] & b[135])^(a[213] & b[136])^(a[212] & b[137])^(a[211] & b[138])^(a[210] & b[139])^(a[209] & b[140])^(a[208] & b[141])^(a[207] & b[142])^(a[206] & b[143])^(a[205] & b[144])^(a[204] & b[145])^(a[203] & b[146])^(a[202] & b[147])^(a[201] & b[148])^(a[200] & b[149])^(a[199] & b[150])^(a[198] & b[151])^(a[197] & b[152])^(a[196] & b[153])^(a[195] & b[154])^(a[194] & b[155])^(a[193] & b[156])^(a[192] & b[157])^(a[191] & b[158])^(a[190] & b[159])^(a[189] & b[160])^(a[188] & b[161])^(a[187] & b[162])^(a[186] & b[163])^(a[185] & b[164])^(a[184] & b[165])^(a[183] & b[166])^(a[182] & b[167])^(a[181] & b[168])^(a[180] & b[169])^(a[179] & b[170])^(a[178] & b[171])^(a[177] & b[172])^(a[176] & b[173])^(a[175] & b[174])^(a[174] & b[175])^(a[173] & b[176])^(a[172] & b[177])^(a[171] & b[178])^(a[170] & b[179])^(a[169] & b[180])^(a[168] & b[181])^(a[167] & b[182])^(a[166] & b[183])^(a[165] & b[184])^(a[164] & b[185])^(a[163] & b[186])^(a[162] & b[187])^(a[161] & b[188])^(a[160] & b[189])^(a[159] & b[190])^(a[158] & b[191])^(a[157] & b[192])^(a[156] & b[193])^(a[155] & b[194])^(a[154] & b[195])^(a[153] & b[196])^(a[152] & b[197])^(a[151] & b[198])^(a[150] & b[199])^(a[149] & b[200])^(a[148] & b[201])^(a[147] & b[202])^(a[146] & b[203])^(a[145] & b[204])^(a[144] & b[205])^(a[143] & b[206])^(a[142] & b[207])^(a[141] & b[208])^(a[140] & b[209])^(a[139] & b[210])^(a[138] & b[211])^(a[137] & b[212])^(a[136] & b[213])^(a[135] & b[214])^(a[134] & b[215])^(a[133] & b[216])^(a[132] & b[217])^(a[131] & b[218])^(a[130] & b[219])^(a[129] & b[220])^(a[128] & b[221])^(a[127] & b[222])^(a[126] & b[223])^(a[125] & b[224])^(a[124] & b[225])^(a[123] & b[226])^(a[122] & b[227])^(a[121] & b[228])^(a[120] & b[229])^(a[119] & b[230])^(a[118] & b[231])^(a[117] & b[232])^(a[116] & b[233])^(a[115] & b[234])^(a[114] & b[235])^(a[113] & b[236])^(a[112] & b[237])^(a[111] & b[238])^(a[110] & b[239])^(a[109] & b[240])^(a[108] & b[241])^(a[107] & b[242])^(a[106] & b[243])^(a[105] & b[244])^(a[104] & b[245])^(a[103] & b[246])^(a[102] & b[247])^(a[101] & b[248])^(a[100] & b[249])^(a[99] & b[250])^(a[98] & b[251])^(a[97] & b[252])^(a[96] & b[253])^(a[95] & b[254])^(a[94] & b[255])^(a[93] & b[256])^(a[92] & b[257])^(a[91] & b[258])^(a[90] & b[259])^(a[89] & b[260])^(a[88] & b[261])^(a[87] & b[262])^(a[86] & b[263])^(a[85] & b[264])^(a[84] & b[265])^(a[83] & b[266])^(a[82] & b[267])^(a[81] & b[268])^(a[80] & b[269])^(a[79] & b[270])^(a[78] & b[271])^(a[77] & b[272])^(a[76] & b[273])^(a[75] & b[274])^(a[74] & b[275])^(a[73] & b[276])^(a[72] & b[277])^(a[71] & b[278])^(a[70] & b[279])^(a[69] & b[280])^(a[68] & b[281])^(a[67] & b[282])^(a[66] & b[283])^(a[65] & b[284])^(a[64] & b[285])^(a[63] & b[286])^(a[62] & b[287])^(a[61] & b[288])^(a[60] & b[289])^(a[59] & b[290])^(a[58] & b[291])^(a[57] & b[292])^(a[56] & b[293])^(a[55] & b[294])^(a[54] & b[295])^(a[53] & b[296])^(a[52] & b[297])^(a[51] & b[298])^(a[50] & b[299])^(a[49] & b[300])^(a[48] & b[301])^(a[47] & b[302])^(a[46] & b[303])^(a[45] & b[304])^(a[44] & b[305])^(a[43] & b[306])^(a[42] & b[307])^(a[41] & b[308])^(a[40] & b[309])^(a[39] & b[310])^(a[38] & b[311])^(a[37] & b[312])^(a[36] & b[313])^(a[35] & b[314])^(a[34] & b[315])^(a[33] & b[316])^(a[32] & b[317])^(a[31] & b[318])^(a[30] & b[319])^(a[29] & b[320])^(a[28] & b[321])^(a[27] & b[322])^(a[26] & b[323])^(a[25] & b[324])^(a[24] & b[325])^(a[23] & b[326])^(a[22] & b[327])^(a[21] & b[328])^(a[20] & b[329])^(a[19] & b[330])^(a[18] & b[331])^(a[17] & b[332])^(a[16] & b[333])^(a[15] & b[334])^(a[14] & b[335])^(a[13] & b[336])^(a[12] & b[337])^(a[11] & b[338])^(a[10] & b[339])^(a[9] & b[340])^(a[8] & b[341])^(a[7] & b[342])^(a[6] & b[343])^(a[5] & b[344])^(a[4] & b[345])^(a[3] & b[346])^(a[2] & b[347])^(a[1] & b[348])^(a[0] & b[349]);
assign y[350] = (a[350] & b[0])^(a[349] & b[1])^(a[348] & b[2])^(a[347] & b[3])^(a[346] & b[4])^(a[345] & b[5])^(a[344] & b[6])^(a[343] & b[7])^(a[342] & b[8])^(a[341] & b[9])^(a[340] & b[10])^(a[339] & b[11])^(a[338] & b[12])^(a[337] & b[13])^(a[336] & b[14])^(a[335] & b[15])^(a[334] & b[16])^(a[333] & b[17])^(a[332] & b[18])^(a[331] & b[19])^(a[330] & b[20])^(a[329] & b[21])^(a[328] & b[22])^(a[327] & b[23])^(a[326] & b[24])^(a[325] & b[25])^(a[324] & b[26])^(a[323] & b[27])^(a[322] & b[28])^(a[321] & b[29])^(a[320] & b[30])^(a[319] & b[31])^(a[318] & b[32])^(a[317] & b[33])^(a[316] & b[34])^(a[315] & b[35])^(a[314] & b[36])^(a[313] & b[37])^(a[312] & b[38])^(a[311] & b[39])^(a[310] & b[40])^(a[309] & b[41])^(a[308] & b[42])^(a[307] & b[43])^(a[306] & b[44])^(a[305] & b[45])^(a[304] & b[46])^(a[303] & b[47])^(a[302] & b[48])^(a[301] & b[49])^(a[300] & b[50])^(a[299] & b[51])^(a[298] & b[52])^(a[297] & b[53])^(a[296] & b[54])^(a[295] & b[55])^(a[294] & b[56])^(a[293] & b[57])^(a[292] & b[58])^(a[291] & b[59])^(a[290] & b[60])^(a[289] & b[61])^(a[288] & b[62])^(a[287] & b[63])^(a[286] & b[64])^(a[285] & b[65])^(a[284] & b[66])^(a[283] & b[67])^(a[282] & b[68])^(a[281] & b[69])^(a[280] & b[70])^(a[279] & b[71])^(a[278] & b[72])^(a[277] & b[73])^(a[276] & b[74])^(a[275] & b[75])^(a[274] & b[76])^(a[273] & b[77])^(a[272] & b[78])^(a[271] & b[79])^(a[270] & b[80])^(a[269] & b[81])^(a[268] & b[82])^(a[267] & b[83])^(a[266] & b[84])^(a[265] & b[85])^(a[264] & b[86])^(a[263] & b[87])^(a[262] & b[88])^(a[261] & b[89])^(a[260] & b[90])^(a[259] & b[91])^(a[258] & b[92])^(a[257] & b[93])^(a[256] & b[94])^(a[255] & b[95])^(a[254] & b[96])^(a[253] & b[97])^(a[252] & b[98])^(a[251] & b[99])^(a[250] & b[100])^(a[249] & b[101])^(a[248] & b[102])^(a[247] & b[103])^(a[246] & b[104])^(a[245] & b[105])^(a[244] & b[106])^(a[243] & b[107])^(a[242] & b[108])^(a[241] & b[109])^(a[240] & b[110])^(a[239] & b[111])^(a[238] & b[112])^(a[237] & b[113])^(a[236] & b[114])^(a[235] & b[115])^(a[234] & b[116])^(a[233] & b[117])^(a[232] & b[118])^(a[231] & b[119])^(a[230] & b[120])^(a[229] & b[121])^(a[228] & b[122])^(a[227] & b[123])^(a[226] & b[124])^(a[225] & b[125])^(a[224] & b[126])^(a[223] & b[127])^(a[222] & b[128])^(a[221] & b[129])^(a[220] & b[130])^(a[219] & b[131])^(a[218] & b[132])^(a[217] & b[133])^(a[216] & b[134])^(a[215] & b[135])^(a[214] & b[136])^(a[213] & b[137])^(a[212] & b[138])^(a[211] & b[139])^(a[210] & b[140])^(a[209] & b[141])^(a[208] & b[142])^(a[207] & b[143])^(a[206] & b[144])^(a[205] & b[145])^(a[204] & b[146])^(a[203] & b[147])^(a[202] & b[148])^(a[201] & b[149])^(a[200] & b[150])^(a[199] & b[151])^(a[198] & b[152])^(a[197] & b[153])^(a[196] & b[154])^(a[195] & b[155])^(a[194] & b[156])^(a[193] & b[157])^(a[192] & b[158])^(a[191] & b[159])^(a[190] & b[160])^(a[189] & b[161])^(a[188] & b[162])^(a[187] & b[163])^(a[186] & b[164])^(a[185] & b[165])^(a[184] & b[166])^(a[183] & b[167])^(a[182] & b[168])^(a[181] & b[169])^(a[180] & b[170])^(a[179] & b[171])^(a[178] & b[172])^(a[177] & b[173])^(a[176] & b[174])^(a[175] & b[175])^(a[174] & b[176])^(a[173] & b[177])^(a[172] & b[178])^(a[171] & b[179])^(a[170] & b[180])^(a[169] & b[181])^(a[168] & b[182])^(a[167] & b[183])^(a[166] & b[184])^(a[165] & b[185])^(a[164] & b[186])^(a[163] & b[187])^(a[162] & b[188])^(a[161] & b[189])^(a[160] & b[190])^(a[159] & b[191])^(a[158] & b[192])^(a[157] & b[193])^(a[156] & b[194])^(a[155] & b[195])^(a[154] & b[196])^(a[153] & b[197])^(a[152] & b[198])^(a[151] & b[199])^(a[150] & b[200])^(a[149] & b[201])^(a[148] & b[202])^(a[147] & b[203])^(a[146] & b[204])^(a[145] & b[205])^(a[144] & b[206])^(a[143] & b[207])^(a[142] & b[208])^(a[141] & b[209])^(a[140] & b[210])^(a[139] & b[211])^(a[138] & b[212])^(a[137] & b[213])^(a[136] & b[214])^(a[135] & b[215])^(a[134] & b[216])^(a[133] & b[217])^(a[132] & b[218])^(a[131] & b[219])^(a[130] & b[220])^(a[129] & b[221])^(a[128] & b[222])^(a[127] & b[223])^(a[126] & b[224])^(a[125] & b[225])^(a[124] & b[226])^(a[123] & b[227])^(a[122] & b[228])^(a[121] & b[229])^(a[120] & b[230])^(a[119] & b[231])^(a[118] & b[232])^(a[117] & b[233])^(a[116] & b[234])^(a[115] & b[235])^(a[114] & b[236])^(a[113] & b[237])^(a[112] & b[238])^(a[111] & b[239])^(a[110] & b[240])^(a[109] & b[241])^(a[108] & b[242])^(a[107] & b[243])^(a[106] & b[244])^(a[105] & b[245])^(a[104] & b[246])^(a[103] & b[247])^(a[102] & b[248])^(a[101] & b[249])^(a[100] & b[250])^(a[99] & b[251])^(a[98] & b[252])^(a[97] & b[253])^(a[96] & b[254])^(a[95] & b[255])^(a[94] & b[256])^(a[93] & b[257])^(a[92] & b[258])^(a[91] & b[259])^(a[90] & b[260])^(a[89] & b[261])^(a[88] & b[262])^(a[87] & b[263])^(a[86] & b[264])^(a[85] & b[265])^(a[84] & b[266])^(a[83] & b[267])^(a[82] & b[268])^(a[81] & b[269])^(a[80] & b[270])^(a[79] & b[271])^(a[78] & b[272])^(a[77] & b[273])^(a[76] & b[274])^(a[75] & b[275])^(a[74] & b[276])^(a[73] & b[277])^(a[72] & b[278])^(a[71] & b[279])^(a[70] & b[280])^(a[69] & b[281])^(a[68] & b[282])^(a[67] & b[283])^(a[66] & b[284])^(a[65] & b[285])^(a[64] & b[286])^(a[63] & b[287])^(a[62] & b[288])^(a[61] & b[289])^(a[60] & b[290])^(a[59] & b[291])^(a[58] & b[292])^(a[57] & b[293])^(a[56] & b[294])^(a[55] & b[295])^(a[54] & b[296])^(a[53] & b[297])^(a[52] & b[298])^(a[51] & b[299])^(a[50] & b[300])^(a[49] & b[301])^(a[48] & b[302])^(a[47] & b[303])^(a[46] & b[304])^(a[45] & b[305])^(a[44] & b[306])^(a[43] & b[307])^(a[42] & b[308])^(a[41] & b[309])^(a[40] & b[310])^(a[39] & b[311])^(a[38] & b[312])^(a[37] & b[313])^(a[36] & b[314])^(a[35] & b[315])^(a[34] & b[316])^(a[33] & b[317])^(a[32] & b[318])^(a[31] & b[319])^(a[30] & b[320])^(a[29] & b[321])^(a[28] & b[322])^(a[27] & b[323])^(a[26] & b[324])^(a[25] & b[325])^(a[24] & b[326])^(a[23] & b[327])^(a[22] & b[328])^(a[21] & b[329])^(a[20] & b[330])^(a[19] & b[331])^(a[18] & b[332])^(a[17] & b[333])^(a[16] & b[334])^(a[15] & b[335])^(a[14] & b[336])^(a[13] & b[337])^(a[12] & b[338])^(a[11] & b[339])^(a[10] & b[340])^(a[9] & b[341])^(a[8] & b[342])^(a[7] & b[343])^(a[6] & b[344])^(a[5] & b[345])^(a[4] & b[346])^(a[3] & b[347])^(a[2] & b[348])^(a[1] & b[349])^(a[0] & b[350]);
assign y[351] = (a[351] & b[0])^(a[350] & b[1])^(a[349] & b[2])^(a[348] & b[3])^(a[347] & b[4])^(a[346] & b[5])^(a[345] & b[6])^(a[344] & b[7])^(a[343] & b[8])^(a[342] & b[9])^(a[341] & b[10])^(a[340] & b[11])^(a[339] & b[12])^(a[338] & b[13])^(a[337] & b[14])^(a[336] & b[15])^(a[335] & b[16])^(a[334] & b[17])^(a[333] & b[18])^(a[332] & b[19])^(a[331] & b[20])^(a[330] & b[21])^(a[329] & b[22])^(a[328] & b[23])^(a[327] & b[24])^(a[326] & b[25])^(a[325] & b[26])^(a[324] & b[27])^(a[323] & b[28])^(a[322] & b[29])^(a[321] & b[30])^(a[320] & b[31])^(a[319] & b[32])^(a[318] & b[33])^(a[317] & b[34])^(a[316] & b[35])^(a[315] & b[36])^(a[314] & b[37])^(a[313] & b[38])^(a[312] & b[39])^(a[311] & b[40])^(a[310] & b[41])^(a[309] & b[42])^(a[308] & b[43])^(a[307] & b[44])^(a[306] & b[45])^(a[305] & b[46])^(a[304] & b[47])^(a[303] & b[48])^(a[302] & b[49])^(a[301] & b[50])^(a[300] & b[51])^(a[299] & b[52])^(a[298] & b[53])^(a[297] & b[54])^(a[296] & b[55])^(a[295] & b[56])^(a[294] & b[57])^(a[293] & b[58])^(a[292] & b[59])^(a[291] & b[60])^(a[290] & b[61])^(a[289] & b[62])^(a[288] & b[63])^(a[287] & b[64])^(a[286] & b[65])^(a[285] & b[66])^(a[284] & b[67])^(a[283] & b[68])^(a[282] & b[69])^(a[281] & b[70])^(a[280] & b[71])^(a[279] & b[72])^(a[278] & b[73])^(a[277] & b[74])^(a[276] & b[75])^(a[275] & b[76])^(a[274] & b[77])^(a[273] & b[78])^(a[272] & b[79])^(a[271] & b[80])^(a[270] & b[81])^(a[269] & b[82])^(a[268] & b[83])^(a[267] & b[84])^(a[266] & b[85])^(a[265] & b[86])^(a[264] & b[87])^(a[263] & b[88])^(a[262] & b[89])^(a[261] & b[90])^(a[260] & b[91])^(a[259] & b[92])^(a[258] & b[93])^(a[257] & b[94])^(a[256] & b[95])^(a[255] & b[96])^(a[254] & b[97])^(a[253] & b[98])^(a[252] & b[99])^(a[251] & b[100])^(a[250] & b[101])^(a[249] & b[102])^(a[248] & b[103])^(a[247] & b[104])^(a[246] & b[105])^(a[245] & b[106])^(a[244] & b[107])^(a[243] & b[108])^(a[242] & b[109])^(a[241] & b[110])^(a[240] & b[111])^(a[239] & b[112])^(a[238] & b[113])^(a[237] & b[114])^(a[236] & b[115])^(a[235] & b[116])^(a[234] & b[117])^(a[233] & b[118])^(a[232] & b[119])^(a[231] & b[120])^(a[230] & b[121])^(a[229] & b[122])^(a[228] & b[123])^(a[227] & b[124])^(a[226] & b[125])^(a[225] & b[126])^(a[224] & b[127])^(a[223] & b[128])^(a[222] & b[129])^(a[221] & b[130])^(a[220] & b[131])^(a[219] & b[132])^(a[218] & b[133])^(a[217] & b[134])^(a[216] & b[135])^(a[215] & b[136])^(a[214] & b[137])^(a[213] & b[138])^(a[212] & b[139])^(a[211] & b[140])^(a[210] & b[141])^(a[209] & b[142])^(a[208] & b[143])^(a[207] & b[144])^(a[206] & b[145])^(a[205] & b[146])^(a[204] & b[147])^(a[203] & b[148])^(a[202] & b[149])^(a[201] & b[150])^(a[200] & b[151])^(a[199] & b[152])^(a[198] & b[153])^(a[197] & b[154])^(a[196] & b[155])^(a[195] & b[156])^(a[194] & b[157])^(a[193] & b[158])^(a[192] & b[159])^(a[191] & b[160])^(a[190] & b[161])^(a[189] & b[162])^(a[188] & b[163])^(a[187] & b[164])^(a[186] & b[165])^(a[185] & b[166])^(a[184] & b[167])^(a[183] & b[168])^(a[182] & b[169])^(a[181] & b[170])^(a[180] & b[171])^(a[179] & b[172])^(a[178] & b[173])^(a[177] & b[174])^(a[176] & b[175])^(a[175] & b[176])^(a[174] & b[177])^(a[173] & b[178])^(a[172] & b[179])^(a[171] & b[180])^(a[170] & b[181])^(a[169] & b[182])^(a[168] & b[183])^(a[167] & b[184])^(a[166] & b[185])^(a[165] & b[186])^(a[164] & b[187])^(a[163] & b[188])^(a[162] & b[189])^(a[161] & b[190])^(a[160] & b[191])^(a[159] & b[192])^(a[158] & b[193])^(a[157] & b[194])^(a[156] & b[195])^(a[155] & b[196])^(a[154] & b[197])^(a[153] & b[198])^(a[152] & b[199])^(a[151] & b[200])^(a[150] & b[201])^(a[149] & b[202])^(a[148] & b[203])^(a[147] & b[204])^(a[146] & b[205])^(a[145] & b[206])^(a[144] & b[207])^(a[143] & b[208])^(a[142] & b[209])^(a[141] & b[210])^(a[140] & b[211])^(a[139] & b[212])^(a[138] & b[213])^(a[137] & b[214])^(a[136] & b[215])^(a[135] & b[216])^(a[134] & b[217])^(a[133] & b[218])^(a[132] & b[219])^(a[131] & b[220])^(a[130] & b[221])^(a[129] & b[222])^(a[128] & b[223])^(a[127] & b[224])^(a[126] & b[225])^(a[125] & b[226])^(a[124] & b[227])^(a[123] & b[228])^(a[122] & b[229])^(a[121] & b[230])^(a[120] & b[231])^(a[119] & b[232])^(a[118] & b[233])^(a[117] & b[234])^(a[116] & b[235])^(a[115] & b[236])^(a[114] & b[237])^(a[113] & b[238])^(a[112] & b[239])^(a[111] & b[240])^(a[110] & b[241])^(a[109] & b[242])^(a[108] & b[243])^(a[107] & b[244])^(a[106] & b[245])^(a[105] & b[246])^(a[104] & b[247])^(a[103] & b[248])^(a[102] & b[249])^(a[101] & b[250])^(a[100] & b[251])^(a[99] & b[252])^(a[98] & b[253])^(a[97] & b[254])^(a[96] & b[255])^(a[95] & b[256])^(a[94] & b[257])^(a[93] & b[258])^(a[92] & b[259])^(a[91] & b[260])^(a[90] & b[261])^(a[89] & b[262])^(a[88] & b[263])^(a[87] & b[264])^(a[86] & b[265])^(a[85] & b[266])^(a[84] & b[267])^(a[83] & b[268])^(a[82] & b[269])^(a[81] & b[270])^(a[80] & b[271])^(a[79] & b[272])^(a[78] & b[273])^(a[77] & b[274])^(a[76] & b[275])^(a[75] & b[276])^(a[74] & b[277])^(a[73] & b[278])^(a[72] & b[279])^(a[71] & b[280])^(a[70] & b[281])^(a[69] & b[282])^(a[68] & b[283])^(a[67] & b[284])^(a[66] & b[285])^(a[65] & b[286])^(a[64] & b[287])^(a[63] & b[288])^(a[62] & b[289])^(a[61] & b[290])^(a[60] & b[291])^(a[59] & b[292])^(a[58] & b[293])^(a[57] & b[294])^(a[56] & b[295])^(a[55] & b[296])^(a[54] & b[297])^(a[53] & b[298])^(a[52] & b[299])^(a[51] & b[300])^(a[50] & b[301])^(a[49] & b[302])^(a[48] & b[303])^(a[47] & b[304])^(a[46] & b[305])^(a[45] & b[306])^(a[44] & b[307])^(a[43] & b[308])^(a[42] & b[309])^(a[41] & b[310])^(a[40] & b[311])^(a[39] & b[312])^(a[38] & b[313])^(a[37] & b[314])^(a[36] & b[315])^(a[35] & b[316])^(a[34] & b[317])^(a[33] & b[318])^(a[32] & b[319])^(a[31] & b[320])^(a[30] & b[321])^(a[29] & b[322])^(a[28] & b[323])^(a[27] & b[324])^(a[26] & b[325])^(a[25] & b[326])^(a[24] & b[327])^(a[23] & b[328])^(a[22] & b[329])^(a[21] & b[330])^(a[20] & b[331])^(a[19] & b[332])^(a[18] & b[333])^(a[17] & b[334])^(a[16] & b[335])^(a[15] & b[336])^(a[14] & b[337])^(a[13] & b[338])^(a[12] & b[339])^(a[11] & b[340])^(a[10] & b[341])^(a[9] & b[342])^(a[8] & b[343])^(a[7] & b[344])^(a[6] & b[345])^(a[5] & b[346])^(a[4] & b[347])^(a[3] & b[348])^(a[2] & b[349])^(a[1] & b[350])^(a[0] & b[351]);
assign y[352] = (a[352] & b[0])^(a[351] & b[1])^(a[350] & b[2])^(a[349] & b[3])^(a[348] & b[4])^(a[347] & b[5])^(a[346] & b[6])^(a[345] & b[7])^(a[344] & b[8])^(a[343] & b[9])^(a[342] & b[10])^(a[341] & b[11])^(a[340] & b[12])^(a[339] & b[13])^(a[338] & b[14])^(a[337] & b[15])^(a[336] & b[16])^(a[335] & b[17])^(a[334] & b[18])^(a[333] & b[19])^(a[332] & b[20])^(a[331] & b[21])^(a[330] & b[22])^(a[329] & b[23])^(a[328] & b[24])^(a[327] & b[25])^(a[326] & b[26])^(a[325] & b[27])^(a[324] & b[28])^(a[323] & b[29])^(a[322] & b[30])^(a[321] & b[31])^(a[320] & b[32])^(a[319] & b[33])^(a[318] & b[34])^(a[317] & b[35])^(a[316] & b[36])^(a[315] & b[37])^(a[314] & b[38])^(a[313] & b[39])^(a[312] & b[40])^(a[311] & b[41])^(a[310] & b[42])^(a[309] & b[43])^(a[308] & b[44])^(a[307] & b[45])^(a[306] & b[46])^(a[305] & b[47])^(a[304] & b[48])^(a[303] & b[49])^(a[302] & b[50])^(a[301] & b[51])^(a[300] & b[52])^(a[299] & b[53])^(a[298] & b[54])^(a[297] & b[55])^(a[296] & b[56])^(a[295] & b[57])^(a[294] & b[58])^(a[293] & b[59])^(a[292] & b[60])^(a[291] & b[61])^(a[290] & b[62])^(a[289] & b[63])^(a[288] & b[64])^(a[287] & b[65])^(a[286] & b[66])^(a[285] & b[67])^(a[284] & b[68])^(a[283] & b[69])^(a[282] & b[70])^(a[281] & b[71])^(a[280] & b[72])^(a[279] & b[73])^(a[278] & b[74])^(a[277] & b[75])^(a[276] & b[76])^(a[275] & b[77])^(a[274] & b[78])^(a[273] & b[79])^(a[272] & b[80])^(a[271] & b[81])^(a[270] & b[82])^(a[269] & b[83])^(a[268] & b[84])^(a[267] & b[85])^(a[266] & b[86])^(a[265] & b[87])^(a[264] & b[88])^(a[263] & b[89])^(a[262] & b[90])^(a[261] & b[91])^(a[260] & b[92])^(a[259] & b[93])^(a[258] & b[94])^(a[257] & b[95])^(a[256] & b[96])^(a[255] & b[97])^(a[254] & b[98])^(a[253] & b[99])^(a[252] & b[100])^(a[251] & b[101])^(a[250] & b[102])^(a[249] & b[103])^(a[248] & b[104])^(a[247] & b[105])^(a[246] & b[106])^(a[245] & b[107])^(a[244] & b[108])^(a[243] & b[109])^(a[242] & b[110])^(a[241] & b[111])^(a[240] & b[112])^(a[239] & b[113])^(a[238] & b[114])^(a[237] & b[115])^(a[236] & b[116])^(a[235] & b[117])^(a[234] & b[118])^(a[233] & b[119])^(a[232] & b[120])^(a[231] & b[121])^(a[230] & b[122])^(a[229] & b[123])^(a[228] & b[124])^(a[227] & b[125])^(a[226] & b[126])^(a[225] & b[127])^(a[224] & b[128])^(a[223] & b[129])^(a[222] & b[130])^(a[221] & b[131])^(a[220] & b[132])^(a[219] & b[133])^(a[218] & b[134])^(a[217] & b[135])^(a[216] & b[136])^(a[215] & b[137])^(a[214] & b[138])^(a[213] & b[139])^(a[212] & b[140])^(a[211] & b[141])^(a[210] & b[142])^(a[209] & b[143])^(a[208] & b[144])^(a[207] & b[145])^(a[206] & b[146])^(a[205] & b[147])^(a[204] & b[148])^(a[203] & b[149])^(a[202] & b[150])^(a[201] & b[151])^(a[200] & b[152])^(a[199] & b[153])^(a[198] & b[154])^(a[197] & b[155])^(a[196] & b[156])^(a[195] & b[157])^(a[194] & b[158])^(a[193] & b[159])^(a[192] & b[160])^(a[191] & b[161])^(a[190] & b[162])^(a[189] & b[163])^(a[188] & b[164])^(a[187] & b[165])^(a[186] & b[166])^(a[185] & b[167])^(a[184] & b[168])^(a[183] & b[169])^(a[182] & b[170])^(a[181] & b[171])^(a[180] & b[172])^(a[179] & b[173])^(a[178] & b[174])^(a[177] & b[175])^(a[176] & b[176])^(a[175] & b[177])^(a[174] & b[178])^(a[173] & b[179])^(a[172] & b[180])^(a[171] & b[181])^(a[170] & b[182])^(a[169] & b[183])^(a[168] & b[184])^(a[167] & b[185])^(a[166] & b[186])^(a[165] & b[187])^(a[164] & b[188])^(a[163] & b[189])^(a[162] & b[190])^(a[161] & b[191])^(a[160] & b[192])^(a[159] & b[193])^(a[158] & b[194])^(a[157] & b[195])^(a[156] & b[196])^(a[155] & b[197])^(a[154] & b[198])^(a[153] & b[199])^(a[152] & b[200])^(a[151] & b[201])^(a[150] & b[202])^(a[149] & b[203])^(a[148] & b[204])^(a[147] & b[205])^(a[146] & b[206])^(a[145] & b[207])^(a[144] & b[208])^(a[143] & b[209])^(a[142] & b[210])^(a[141] & b[211])^(a[140] & b[212])^(a[139] & b[213])^(a[138] & b[214])^(a[137] & b[215])^(a[136] & b[216])^(a[135] & b[217])^(a[134] & b[218])^(a[133] & b[219])^(a[132] & b[220])^(a[131] & b[221])^(a[130] & b[222])^(a[129] & b[223])^(a[128] & b[224])^(a[127] & b[225])^(a[126] & b[226])^(a[125] & b[227])^(a[124] & b[228])^(a[123] & b[229])^(a[122] & b[230])^(a[121] & b[231])^(a[120] & b[232])^(a[119] & b[233])^(a[118] & b[234])^(a[117] & b[235])^(a[116] & b[236])^(a[115] & b[237])^(a[114] & b[238])^(a[113] & b[239])^(a[112] & b[240])^(a[111] & b[241])^(a[110] & b[242])^(a[109] & b[243])^(a[108] & b[244])^(a[107] & b[245])^(a[106] & b[246])^(a[105] & b[247])^(a[104] & b[248])^(a[103] & b[249])^(a[102] & b[250])^(a[101] & b[251])^(a[100] & b[252])^(a[99] & b[253])^(a[98] & b[254])^(a[97] & b[255])^(a[96] & b[256])^(a[95] & b[257])^(a[94] & b[258])^(a[93] & b[259])^(a[92] & b[260])^(a[91] & b[261])^(a[90] & b[262])^(a[89] & b[263])^(a[88] & b[264])^(a[87] & b[265])^(a[86] & b[266])^(a[85] & b[267])^(a[84] & b[268])^(a[83] & b[269])^(a[82] & b[270])^(a[81] & b[271])^(a[80] & b[272])^(a[79] & b[273])^(a[78] & b[274])^(a[77] & b[275])^(a[76] & b[276])^(a[75] & b[277])^(a[74] & b[278])^(a[73] & b[279])^(a[72] & b[280])^(a[71] & b[281])^(a[70] & b[282])^(a[69] & b[283])^(a[68] & b[284])^(a[67] & b[285])^(a[66] & b[286])^(a[65] & b[287])^(a[64] & b[288])^(a[63] & b[289])^(a[62] & b[290])^(a[61] & b[291])^(a[60] & b[292])^(a[59] & b[293])^(a[58] & b[294])^(a[57] & b[295])^(a[56] & b[296])^(a[55] & b[297])^(a[54] & b[298])^(a[53] & b[299])^(a[52] & b[300])^(a[51] & b[301])^(a[50] & b[302])^(a[49] & b[303])^(a[48] & b[304])^(a[47] & b[305])^(a[46] & b[306])^(a[45] & b[307])^(a[44] & b[308])^(a[43] & b[309])^(a[42] & b[310])^(a[41] & b[311])^(a[40] & b[312])^(a[39] & b[313])^(a[38] & b[314])^(a[37] & b[315])^(a[36] & b[316])^(a[35] & b[317])^(a[34] & b[318])^(a[33] & b[319])^(a[32] & b[320])^(a[31] & b[321])^(a[30] & b[322])^(a[29] & b[323])^(a[28] & b[324])^(a[27] & b[325])^(a[26] & b[326])^(a[25] & b[327])^(a[24] & b[328])^(a[23] & b[329])^(a[22] & b[330])^(a[21] & b[331])^(a[20] & b[332])^(a[19] & b[333])^(a[18] & b[334])^(a[17] & b[335])^(a[16] & b[336])^(a[15] & b[337])^(a[14] & b[338])^(a[13] & b[339])^(a[12] & b[340])^(a[11] & b[341])^(a[10] & b[342])^(a[9] & b[343])^(a[8] & b[344])^(a[7] & b[345])^(a[6] & b[346])^(a[5] & b[347])^(a[4] & b[348])^(a[3] & b[349])^(a[2] & b[350])^(a[1] & b[351])^(a[0] & b[352]);
assign y[353] = (a[353] & b[0])^(a[352] & b[1])^(a[351] & b[2])^(a[350] & b[3])^(a[349] & b[4])^(a[348] & b[5])^(a[347] & b[6])^(a[346] & b[7])^(a[345] & b[8])^(a[344] & b[9])^(a[343] & b[10])^(a[342] & b[11])^(a[341] & b[12])^(a[340] & b[13])^(a[339] & b[14])^(a[338] & b[15])^(a[337] & b[16])^(a[336] & b[17])^(a[335] & b[18])^(a[334] & b[19])^(a[333] & b[20])^(a[332] & b[21])^(a[331] & b[22])^(a[330] & b[23])^(a[329] & b[24])^(a[328] & b[25])^(a[327] & b[26])^(a[326] & b[27])^(a[325] & b[28])^(a[324] & b[29])^(a[323] & b[30])^(a[322] & b[31])^(a[321] & b[32])^(a[320] & b[33])^(a[319] & b[34])^(a[318] & b[35])^(a[317] & b[36])^(a[316] & b[37])^(a[315] & b[38])^(a[314] & b[39])^(a[313] & b[40])^(a[312] & b[41])^(a[311] & b[42])^(a[310] & b[43])^(a[309] & b[44])^(a[308] & b[45])^(a[307] & b[46])^(a[306] & b[47])^(a[305] & b[48])^(a[304] & b[49])^(a[303] & b[50])^(a[302] & b[51])^(a[301] & b[52])^(a[300] & b[53])^(a[299] & b[54])^(a[298] & b[55])^(a[297] & b[56])^(a[296] & b[57])^(a[295] & b[58])^(a[294] & b[59])^(a[293] & b[60])^(a[292] & b[61])^(a[291] & b[62])^(a[290] & b[63])^(a[289] & b[64])^(a[288] & b[65])^(a[287] & b[66])^(a[286] & b[67])^(a[285] & b[68])^(a[284] & b[69])^(a[283] & b[70])^(a[282] & b[71])^(a[281] & b[72])^(a[280] & b[73])^(a[279] & b[74])^(a[278] & b[75])^(a[277] & b[76])^(a[276] & b[77])^(a[275] & b[78])^(a[274] & b[79])^(a[273] & b[80])^(a[272] & b[81])^(a[271] & b[82])^(a[270] & b[83])^(a[269] & b[84])^(a[268] & b[85])^(a[267] & b[86])^(a[266] & b[87])^(a[265] & b[88])^(a[264] & b[89])^(a[263] & b[90])^(a[262] & b[91])^(a[261] & b[92])^(a[260] & b[93])^(a[259] & b[94])^(a[258] & b[95])^(a[257] & b[96])^(a[256] & b[97])^(a[255] & b[98])^(a[254] & b[99])^(a[253] & b[100])^(a[252] & b[101])^(a[251] & b[102])^(a[250] & b[103])^(a[249] & b[104])^(a[248] & b[105])^(a[247] & b[106])^(a[246] & b[107])^(a[245] & b[108])^(a[244] & b[109])^(a[243] & b[110])^(a[242] & b[111])^(a[241] & b[112])^(a[240] & b[113])^(a[239] & b[114])^(a[238] & b[115])^(a[237] & b[116])^(a[236] & b[117])^(a[235] & b[118])^(a[234] & b[119])^(a[233] & b[120])^(a[232] & b[121])^(a[231] & b[122])^(a[230] & b[123])^(a[229] & b[124])^(a[228] & b[125])^(a[227] & b[126])^(a[226] & b[127])^(a[225] & b[128])^(a[224] & b[129])^(a[223] & b[130])^(a[222] & b[131])^(a[221] & b[132])^(a[220] & b[133])^(a[219] & b[134])^(a[218] & b[135])^(a[217] & b[136])^(a[216] & b[137])^(a[215] & b[138])^(a[214] & b[139])^(a[213] & b[140])^(a[212] & b[141])^(a[211] & b[142])^(a[210] & b[143])^(a[209] & b[144])^(a[208] & b[145])^(a[207] & b[146])^(a[206] & b[147])^(a[205] & b[148])^(a[204] & b[149])^(a[203] & b[150])^(a[202] & b[151])^(a[201] & b[152])^(a[200] & b[153])^(a[199] & b[154])^(a[198] & b[155])^(a[197] & b[156])^(a[196] & b[157])^(a[195] & b[158])^(a[194] & b[159])^(a[193] & b[160])^(a[192] & b[161])^(a[191] & b[162])^(a[190] & b[163])^(a[189] & b[164])^(a[188] & b[165])^(a[187] & b[166])^(a[186] & b[167])^(a[185] & b[168])^(a[184] & b[169])^(a[183] & b[170])^(a[182] & b[171])^(a[181] & b[172])^(a[180] & b[173])^(a[179] & b[174])^(a[178] & b[175])^(a[177] & b[176])^(a[176] & b[177])^(a[175] & b[178])^(a[174] & b[179])^(a[173] & b[180])^(a[172] & b[181])^(a[171] & b[182])^(a[170] & b[183])^(a[169] & b[184])^(a[168] & b[185])^(a[167] & b[186])^(a[166] & b[187])^(a[165] & b[188])^(a[164] & b[189])^(a[163] & b[190])^(a[162] & b[191])^(a[161] & b[192])^(a[160] & b[193])^(a[159] & b[194])^(a[158] & b[195])^(a[157] & b[196])^(a[156] & b[197])^(a[155] & b[198])^(a[154] & b[199])^(a[153] & b[200])^(a[152] & b[201])^(a[151] & b[202])^(a[150] & b[203])^(a[149] & b[204])^(a[148] & b[205])^(a[147] & b[206])^(a[146] & b[207])^(a[145] & b[208])^(a[144] & b[209])^(a[143] & b[210])^(a[142] & b[211])^(a[141] & b[212])^(a[140] & b[213])^(a[139] & b[214])^(a[138] & b[215])^(a[137] & b[216])^(a[136] & b[217])^(a[135] & b[218])^(a[134] & b[219])^(a[133] & b[220])^(a[132] & b[221])^(a[131] & b[222])^(a[130] & b[223])^(a[129] & b[224])^(a[128] & b[225])^(a[127] & b[226])^(a[126] & b[227])^(a[125] & b[228])^(a[124] & b[229])^(a[123] & b[230])^(a[122] & b[231])^(a[121] & b[232])^(a[120] & b[233])^(a[119] & b[234])^(a[118] & b[235])^(a[117] & b[236])^(a[116] & b[237])^(a[115] & b[238])^(a[114] & b[239])^(a[113] & b[240])^(a[112] & b[241])^(a[111] & b[242])^(a[110] & b[243])^(a[109] & b[244])^(a[108] & b[245])^(a[107] & b[246])^(a[106] & b[247])^(a[105] & b[248])^(a[104] & b[249])^(a[103] & b[250])^(a[102] & b[251])^(a[101] & b[252])^(a[100] & b[253])^(a[99] & b[254])^(a[98] & b[255])^(a[97] & b[256])^(a[96] & b[257])^(a[95] & b[258])^(a[94] & b[259])^(a[93] & b[260])^(a[92] & b[261])^(a[91] & b[262])^(a[90] & b[263])^(a[89] & b[264])^(a[88] & b[265])^(a[87] & b[266])^(a[86] & b[267])^(a[85] & b[268])^(a[84] & b[269])^(a[83] & b[270])^(a[82] & b[271])^(a[81] & b[272])^(a[80] & b[273])^(a[79] & b[274])^(a[78] & b[275])^(a[77] & b[276])^(a[76] & b[277])^(a[75] & b[278])^(a[74] & b[279])^(a[73] & b[280])^(a[72] & b[281])^(a[71] & b[282])^(a[70] & b[283])^(a[69] & b[284])^(a[68] & b[285])^(a[67] & b[286])^(a[66] & b[287])^(a[65] & b[288])^(a[64] & b[289])^(a[63] & b[290])^(a[62] & b[291])^(a[61] & b[292])^(a[60] & b[293])^(a[59] & b[294])^(a[58] & b[295])^(a[57] & b[296])^(a[56] & b[297])^(a[55] & b[298])^(a[54] & b[299])^(a[53] & b[300])^(a[52] & b[301])^(a[51] & b[302])^(a[50] & b[303])^(a[49] & b[304])^(a[48] & b[305])^(a[47] & b[306])^(a[46] & b[307])^(a[45] & b[308])^(a[44] & b[309])^(a[43] & b[310])^(a[42] & b[311])^(a[41] & b[312])^(a[40] & b[313])^(a[39] & b[314])^(a[38] & b[315])^(a[37] & b[316])^(a[36] & b[317])^(a[35] & b[318])^(a[34] & b[319])^(a[33] & b[320])^(a[32] & b[321])^(a[31] & b[322])^(a[30] & b[323])^(a[29] & b[324])^(a[28] & b[325])^(a[27] & b[326])^(a[26] & b[327])^(a[25] & b[328])^(a[24] & b[329])^(a[23] & b[330])^(a[22] & b[331])^(a[21] & b[332])^(a[20] & b[333])^(a[19] & b[334])^(a[18] & b[335])^(a[17] & b[336])^(a[16] & b[337])^(a[15] & b[338])^(a[14] & b[339])^(a[13] & b[340])^(a[12] & b[341])^(a[11] & b[342])^(a[10] & b[343])^(a[9] & b[344])^(a[8] & b[345])^(a[7] & b[346])^(a[6] & b[347])^(a[5] & b[348])^(a[4] & b[349])^(a[3] & b[350])^(a[2] & b[351])^(a[1] & b[352])^(a[0] & b[353]);
assign y[354] = (a[354] & b[0])^(a[353] & b[1])^(a[352] & b[2])^(a[351] & b[3])^(a[350] & b[4])^(a[349] & b[5])^(a[348] & b[6])^(a[347] & b[7])^(a[346] & b[8])^(a[345] & b[9])^(a[344] & b[10])^(a[343] & b[11])^(a[342] & b[12])^(a[341] & b[13])^(a[340] & b[14])^(a[339] & b[15])^(a[338] & b[16])^(a[337] & b[17])^(a[336] & b[18])^(a[335] & b[19])^(a[334] & b[20])^(a[333] & b[21])^(a[332] & b[22])^(a[331] & b[23])^(a[330] & b[24])^(a[329] & b[25])^(a[328] & b[26])^(a[327] & b[27])^(a[326] & b[28])^(a[325] & b[29])^(a[324] & b[30])^(a[323] & b[31])^(a[322] & b[32])^(a[321] & b[33])^(a[320] & b[34])^(a[319] & b[35])^(a[318] & b[36])^(a[317] & b[37])^(a[316] & b[38])^(a[315] & b[39])^(a[314] & b[40])^(a[313] & b[41])^(a[312] & b[42])^(a[311] & b[43])^(a[310] & b[44])^(a[309] & b[45])^(a[308] & b[46])^(a[307] & b[47])^(a[306] & b[48])^(a[305] & b[49])^(a[304] & b[50])^(a[303] & b[51])^(a[302] & b[52])^(a[301] & b[53])^(a[300] & b[54])^(a[299] & b[55])^(a[298] & b[56])^(a[297] & b[57])^(a[296] & b[58])^(a[295] & b[59])^(a[294] & b[60])^(a[293] & b[61])^(a[292] & b[62])^(a[291] & b[63])^(a[290] & b[64])^(a[289] & b[65])^(a[288] & b[66])^(a[287] & b[67])^(a[286] & b[68])^(a[285] & b[69])^(a[284] & b[70])^(a[283] & b[71])^(a[282] & b[72])^(a[281] & b[73])^(a[280] & b[74])^(a[279] & b[75])^(a[278] & b[76])^(a[277] & b[77])^(a[276] & b[78])^(a[275] & b[79])^(a[274] & b[80])^(a[273] & b[81])^(a[272] & b[82])^(a[271] & b[83])^(a[270] & b[84])^(a[269] & b[85])^(a[268] & b[86])^(a[267] & b[87])^(a[266] & b[88])^(a[265] & b[89])^(a[264] & b[90])^(a[263] & b[91])^(a[262] & b[92])^(a[261] & b[93])^(a[260] & b[94])^(a[259] & b[95])^(a[258] & b[96])^(a[257] & b[97])^(a[256] & b[98])^(a[255] & b[99])^(a[254] & b[100])^(a[253] & b[101])^(a[252] & b[102])^(a[251] & b[103])^(a[250] & b[104])^(a[249] & b[105])^(a[248] & b[106])^(a[247] & b[107])^(a[246] & b[108])^(a[245] & b[109])^(a[244] & b[110])^(a[243] & b[111])^(a[242] & b[112])^(a[241] & b[113])^(a[240] & b[114])^(a[239] & b[115])^(a[238] & b[116])^(a[237] & b[117])^(a[236] & b[118])^(a[235] & b[119])^(a[234] & b[120])^(a[233] & b[121])^(a[232] & b[122])^(a[231] & b[123])^(a[230] & b[124])^(a[229] & b[125])^(a[228] & b[126])^(a[227] & b[127])^(a[226] & b[128])^(a[225] & b[129])^(a[224] & b[130])^(a[223] & b[131])^(a[222] & b[132])^(a[221] & b[133])^(a[220] & b[134])^(a[219] & b[135])^(a[218] & b[136])^(a[217] & b[137])^(a[216] & b[138])^(a[215] & b[139])^(a[214] & b[140])^(a[213] & b[141])^(a[212] & b[142])^(a[211] & b[143])^(a[210] & b[144])^(a[209] & b[145])^(a[208] & b[146])^(a[207] & b[147])^(a[206] & b[148])^(a[205] & b[149])^(a[204] & b[150])^(a[203] & b[151])^(a[202] & b[152])^(a[201] & b[153])^(a[200] & b[154])^(a[199] & b[155])^(a[198] & b[156])^(a[197] & b[157])^(a[196] & b[158])^(a[195] & b[159])^(a[194] & b[160])^(a[193] & b[161])^(a[192] & b[162])^(a[191] & b[163])^(a[190] & b[164])^(a[189] & b[165])^(a[188] & b[166])^(a[187] & b[167])^(a[186] & b[168])^(a[185] & b[169])^(a[184] & b[170])^(a[183] & b[171])^(a[182] & b[172])^(a[181] & b[173])^(a[180] & b[174])^(a[179] & b[175])^(a[178] & b[176])^(a[177] & b[177])^(a[176] & b[178])^(a[175] & b[179])^(a[174] & b[180])^(a[173] & b[181])^(a[172] & b[182])^(a[171] & b[183])^(a[170] & b[184])^(a[169] & b[185])^(a[168] & b[186])^(a[167] & b[187])^(a[166] & b[188])^(a[165] & b[189])^(a[164] & b[190])^(a[163] & b[191])^(a[162] & b[192])^(a[161] & b[193])^(a[160] & b[194])^(a[159] & b[195])^(a[158] & b[196])^(a[157] & b[197])^(a[156] & b[198])^(a[155] & b[199])^(a[154] & b[200])^(a[153] & b[201])^(a[152] & b[202])^(a[151] & b[203])^(a[150] & b[204])^(a[149] & b[205])^(a[148] & b[206])^(a[147] & b[207])^(a[146] & b[208])^(a[145] & b[209])^(a[144] & b[210])^(a[143] & b[211])^(a[142] & b[212])^(a[141] & b[213])^(a[140] & b[214])^(a[139] & b[215])^(a[138] & b[216])^(a[137] & b[217])^(a[136] & b[218])^(a[135] & b[219])^(a[134] & b[220])^(a[133] & b[221])^(a[132] & b[222])^(a[131] & b[223])^(a[130] & b[224])^(a[129] & b[225])^(a[128] & b[226])^(a[127] & b[227])^(a[126] & b[228])^(a[125] & b[229])^(a[124] & b[230])^(a[123] & b[231])^(a[122] & b[232])^(a[121] & b[233])^(a[120] & b[234])^(a[119] & b[235])^(a[118] & b[236])^(a[117] & b[237])^(a[116] & b[238])^(a[115] & b[239])^(a[114] & b[240])^(a[113] & b[241])^(a[112] & b[242])^(a[111] & b[243])^(a[110] & b[244])^(a[109] & b[245])^(a[108] & b[246])^(a[107] & b[247])^(a[106] & b[248])^(a[105] & b[249])^(a[104] & b[250])^(a[103] & b[251])^(a[102] & b[252])^(a[101] & b[253])^(a[100] & b[254])^(a[99] & b[255])^(a[98] & b[256])^(a[97] & b[257])^(a[96] & b[258])^(a[95] & b[259])^(a[94] & b[260])^(a[93] & b[261])^(a[92] & b[262])^(a[91] & b[263])^(a[90] & b[264])^(a[89] & b[265])^(a[88] & b[266])^(a[87] & b[267])^(a[86] & b[268])^(a[85] & b[269])^(a[84] & b[270])^(a[83] & b[271])^(a[82] & b[272])^(a[81] & b[273])^(a[80] & b[274])^(a[79] & b[275])^(a[78] & b[276])^(a[77] & b[277])^(a[76] & b[278])^(a[75] & b[279])^(a[74] & b[280])^(a[73] & b[281])^(a[72] & b[282])^(a[71] & b[283])^(a[70] & b[284])^(a[69] & b[285])^(a[68] & b[286])^(a[67] & b[287])^(a[66] & b[288])^(a[65] & b[289])^(a[64] & b[290])^(a[63] & b[291])^(a[62] & b[292])^(a[61] & b[293])^(a[60] & b[294])^(a[59] & b[295])^(a[58] & b[296])^(a[57] & b[297])^(a[56] & b[298])^(a[55] & b[299])^(a[54] & b[300])^(a[53] & b[301])^(a[52] & b[302])^(a[51] & b[303])^(a[50] & b[304])^(a[49] & b[305])^(a[48] & b[306])^(a[47] & b[307])^(a[46] & b[308])^(a[45] & b[309])^(a[44] & b[310])^(a[43] & b[311])^(a[42] & b[312])^(a[41] & b[313])^(a[40] & b[314])^(a[39] & b[315])^(a[38] & b[316])^(a[37] & b[317])^(a[36] & b[318])^(a[35] & b[319])^(a[34] & b[320])^(a[33] & b[321])^(a[32] & b[322])^(a[31] & b[323])^(a[30] & b[324])^(a[29] & b[325])^(a[28] & b[326])^(a[27] & b[327])^(a[26] & b[328])^(a[25] & b[329])^(a[24] & b[330])^(a[23] & b[331])^(a[22] & b[332])^(a[21] & b[333])^(a[20] & b[334])^(a[19] & b[335])^(a[18] & b[336])^(a[17] & b[337])^(a[16] & b[338])^(a[15] & b[339])^(a[14] & b[340])^(a[13] & b[341])^(a[12] & b[342])^(a[11] & b[343])^(a[10] & b[344])^(a[9] & b[345])^(a[8] & b[346])^(a[7] & b[347])^(a[6] & b[348])^(a[5] & b[349])^(a[4] & b[350])^(a[3] & b[351])^(a[2] & b[352])^(a[1] & b[353])^(a[0] & b[354]);
assign y[355] = (a[355] & b[0])^(a[354] & b[1])^(a[353] & b[2])^(a[352] & b[3])^(a[351] & b[4])^(a[350] & b[5])^(a[349] & b[6])^(a[348] & b[7])^(a[347] & b[8])^(a[346] & b[9])^(a[345] & b[10])^(a[344] & b[11])^(a[343] & b[12])^(a[342] & b[13])^(a[341] & b[14])^(a[340] & b[15])^(a[339] & b[16])^(a[338] & b[17])^(a[337] & b[18])^(a[336] & b[19])^(a[335] & b[20])^(a[334] & b[21])^(a[333] & b[22])^(a[332] & b[23])^(a[331] & b[24])^(a[330] & b[25])^(a[329] & b[26])^(a[328] & b[27])^(a[327] & b[28])^(a[326] & b[29])^(a[325] & b[30])^(a[324] & b[31])^(a[323] & b[32])^(a[322] & b[33])^(a[321] & b[34])^(a[320] & b[35])^(a[319] & b[36])^(a[318] & b[37])^(a[317] & b[38])^(a[316] & b[39])^(a[315] & b[40])^(a[314] & b[41])^(a[313] & b[42])^(a[312] & b[43])^(a[311] & b[44])^(a[310] & b[45])^(a[309] & b[46])^(a[308] & b[47])^(a[307] & b[48])^(a[306] & b[49])^(a[305] & b[50])^(a[304] & b[51])^(a[303] & b[52])^(a[302] & b[53])^(a[301] & b[54])^(a[300] & b[55])^(a[299] & b[56])^(a[298] & b[57])^(a[297] & b[58])^(a[296] & b[59])^(a[295] & b[60])^(a[294] & b[61])^(a[293] & b[62])^(a[292] & b[63])^(a[291] & b[64])^(a[290] & b[65])^(a[289] & b[66])^(a[288] & b[67])^(a[287] & b[68])^(a[286] & b[69])^(a[285] & b[70])^(a[284] & b[71])^(a[283] & b[72])^(a[282] & b[73])^(a[281] & b[74])^(a[280] & b[75])^(a[279] & b[76])^(a[278] & b[77])^(a[277] & b[78])^(a[276] & b[79])^(a[275] & b[80])^(a[274] & b[81])^(a[273] & b[82])^(a[272] & b[83])^(a[271] & b[84])^(a[270] & b[85])^(a[269] & b[86])^(a[268] & b[87])^(a[267] & b[88])^(a[266] & b[89])^(a[265] & b[90])^(a[264] & b[91])^(a[263] & b[92])^(a[262] & b[93])^(a[261] & b[94])^(a[260] & b[95])^(a[259] & b[96])^(a[258] & b[97])^(a[257] & b[98])^(a[256] & b[99])^(a[255] & b[100])^(a[254] & b[101])^(a[253] & b[102])^(a[252] & b[103])^(a[251] & b[104])^(a[250] & b[105])^(a[249] & b[106])^(a[248] & b[107])^(a[247] & b[108])^(a[246] & b[109])^(a[245] & b[110])^(a[244] & b[111])^(a[243] & b[112])^(a[242] & b[113])^(a[241] & b[114])^(a[240] & b[115])^(a[239] & b[116])^(a[238] & b[117])^(a[237] & b[118])^(a[236] & b[119])^(a[235] & b[120])^(a[234] & b[121])^(a[233] & b[122])^(a[232] & b[123])^(a[231] & b[124])^(a[230] & b[125])^(a[229] & b[126])^(a[228] & b[127])^(a[227] & b[128])^(a[226] & b[129])^(a[225] & b[130])^(a[224] & b[131])^(a[223] & b[132])^(a[222] & b[133])^(a[221] & b[134])^(a[220] & b[135])^(a[219] & b[136])^(a[218] & b[137])^(a[217] & b[138])^(a[216] & b[139])^(a[215] & b[140])^(a[214] & b[141])^(a[213] & b[142])^(a[212] & b[143])^(a[211] & b[144])^(a[210] & b[145])^(a[209] & b[146])^(a[208] & b[147])^(a[207] & b[148])^(a[206] & b[149])^(a[205] & b[150])^(a[204] & b[151])^(a[203] & b[152])^(a[202] & b[153])^(a[201] & b[154])^(a[200] & b[155])^(a[199] & b[156])^(a[198] & b[157])^(a[197] & b[158])^(a[196] & b[159])^(a[195] & b[160])^(a[194] & b[161])^(a[193] & b[162])^(a[192] & b[163])^(a[191] & b[164])^(a[190] & b[165])^(a[189] & b[166])^(a[188] & b[167])^(a[187] & b[168])^(a[186] & b[169])^(a[185] & b[170])^(a[184] & b[171])^(a[183] & b[172])^(a[182] & b[173])^(a[181] & b[174])^(a[180] & b[175])^(a[179] & b[176])^(a[178] & b[177])^(a[177] & b[178])^(a[176] & b[179])^(a[175] & b[180])^(a[174] & b[181])^(a[173] & b[182])^(a[172] & b[183])^(a[171] & b[184])^(a[170] & b[185])^(a[169] & b[186])^(a[168] & b[187])^(a[167] & b[188])^(a[166] & b[189])^(a[165] & b[190])^(a[164] & b[191])^(a[163] & b[192])^(a[162] & b[193])^(a[161] & b[194])^(a[160] & b[195])^(a[159] & b[196])^(a[158] & b[197])^(a[157] & b[198])^(a[156] & b[199])^(a[155] & b[200])^(a[154] & b[201])^(a[153] & b[202])^(a[152] & b[203])^(a[151] & b[204])^(a[150] & b[205])^(a[149] & b[206])^(a[148] & b[207])^(a[147] & b[208])^(a[146] & b[209])^(a[145] & b[210])^(a[144] & b[211])^(a[143] & b[212])^(a[142] & b[213])^(a[141] & b[214])^(a[140] & b[215])^(a[139] & b[216])^(a[138] & b[217])^(a[137] & b[218])^(a[136] & b[219])^(a[135] & b[220])^(a[134] & b[221])^(a[133] & b[222])^(a[132] & b[223])^(a[131] & b[224])^(a[130] & b[225])^(a[129] & b[226])^(a[128] & b[227])^(a[127] & b[228])^(a[126] & b[229])^(a[125] & b[230])^(a[124] & b[231])^(a[123] & b[232])^(a[122] & b[233])^(a[121] & b[234])^(a[120] & b[235])^(a[119] & b[236])^(a[118] & b[237])^(a[117] & b[238])^(a[116] & b[239])^(a[115] & b[240])^(a[114] & b[241])^(a[113] & b[242])^(a[112] & b[243])^(a[111] & b[244])^(a[110] & b[245])^(a[109] & b[246])^(a[108] & b[247])^(a[107] & b[248])^(a[106] & b[249])^(a[105] & b[250])^(a[104] & b[251])^(a[103] & b[252])^(a[102] & b[253])^(a[101] & b[254])^(a[100] & b[255])^(a[99] & b[256])^(a[98] & b[257])^(a[97] & b[258])^(a[96] & b[259])^(a[95] & b[260])^(a[94] & b[261])^(a[93] & b[262])^(a[92] & b[263])^(a[91] & b[264])^(a[90] & b[265])^(a[89] & b[266])^(a[88] & b[267])^(a[87] & b[268])^(a[86] & b[269])^(a[85] & b[270])^(a[84] & b[271])^(a[83] & b[272])^(a[82] & b[273])^(a[81] & b[274])^(a[80] & b[275])^(a[79] & b[276])^(a[78] & b[277])^(a[77] & b[278])^(a[76] & b[279])^(a[75] & b[280])^(a[74] & b[281])^(a[73] & b[282])^(a[72] & b[283])^(a[71] & b[284])^(a[70] & b[285])^(a[69] & b[286])^(a[68] & b[287])^(a[67] & b[288])^(a[66] & b[289])^(a[65] & b[290])^(a[64] & b[291])^(a[63] & b[292])^(a[62] & b[293])^(a[61] & b[294])^(a[60] & b[295])^(a[59] & b[296])^(a[58] & b[297])^(a[57] & b[298])^(a[56] & b[299])^(a[55] & b[300])^(a[54] & b[301])^(a[53] & b[302])^(a[52] & b[303])^(a[51] & b[304])^(a[50] & b[305])^(a[49] & b[306])^(a[48] & b[307])^(a[47] & b[308])^(a[46] & b[309])^(a[45] & b[310])^(a[44] & b[311])^(a[43] & b[312])^(a[42] & b[313])^(a[41] & b[314])^(a[40] & b[315])^(a[39] & b[316])^(a[38] & b[317])^(a[37] & b[318])^(a[36] & b[319])^(a[35] & b[320])^(a[34] & b[321])^(a[33] & b[322])^(a[32] & b[323])^(a[31] & b[324])^(a[30] & b[325])^(a[29] & b[326])^(a[28] & b[327])^(a[27] & b[328])^(a[26] & b[329])^(a[25] & b[330])^(a[24] & b[331])^(a[23] & b[332])^(a[22] & b[333])^(a[21] & b[334])^(a[20] & b[335])^(a[19] & b[336])^(a[18] & b[337])^(a[17] & b[338])^(a[16] & b[339])^(a[15] & b[340])^(a[14] & b[341])^(a[13] & b[342])^(a[12] & b[343])^(a[11] & b[344])^(a[10] & b[345])^(a[9] & b[346])^(a[8] & b[347])^(a[7] & b[348])^(a[6] & b[349])^(a[5] & b[350])^(a[4] & b[351])^(a[3] & b[352])^(a[2] & b[353])^(a[1] & b[354])^(a[0] & b[355]);
assign y[356] = (a[356] & b[0])^(a[355] & b[1])^(a[354] & b[2])^(a[353] & b[3])^(a[352] & b[4])^(a[351] & b[5])^(a[350] & b[6])^(a[349] & b[7])^(a[348] & b[8])^(a[347] & b[9])^(a[346] & b[10])^(a[345] & b[11])^(a[344] & b[12])^(a[343] & b[13])^(a[342] & b[14])^(a[341] & b[15])^(a[340] & b[16])^(a[339] & b[17])^(a[338] & b[18])^(a[337] & b[19])^(a[336] & b[20])^(a[335] & b[21])^(a[334] & b[22])^(a[333] & b[23])^(a[332] & b[24])^(a[331] & b[25])^(a[330] & b[26])^(a[329] & b[27])^(a[328] & b[28])^(a[327] & b[29])^(a[326] & b[30])^(a[325] & b[31])^(a[324] & b[32])^(a[323] & b[33])^(a[322] & b[34])^(a[321] & b[35])^(a[320] & b[36])^(a[319] & b[37])^(a[318] & b[38])^(a[317] & b[39])^(a[316] & b[40])^(a[315] & b[41])^(a[314] & b[42])^(a[313] & b[43])^(a[312] & b[44])^(a[311] & b[45])^(a[310] & b[46])^(a[309] & b[47])^(a[308] & b[48])^(a[307] & b[49])^(a[306] & b[50])^(a[305] & b[51])^(a[304] & b[52])^(a[303] & b[53])^(a[302] & b[54])^(a[301] & b[55])^(a[300] & b[56])^(a[299] & b[57])^(a[298] & b[58])^(a[297] & b[59])^(a[296] & b[60])^(a[295] & b[61])^(a[294] & b[62])^(a[293] & b[63])^(a[292] & b[64])^(a[291] & b[65])^(a[290] & b[66])^(a[289] & b[67])^(a[288] & b[68])^(a[287] & b[69])^(a[286] & b[70])^(a[285] & b[71])^(a[284] & b[72])^(a[283] & b[73])^(a[282] & b[74])^(a[281] & b[75])^(a[280] & b[76])^(a[279] & b[77])^(a[278] & b[78])^(a[277] & b[79])^(a[276] & b[80])^(a[275] & b[81])^(a[274] & b[82])^(a[273] & b[83])^(a[272] & b[84])^(a[271] & b[85])^(a[270] & b[86])^(a[269] & b[87])^(a[268] & b[88])^(a[267] & b[89])^(a[266] & b[90])^(a[265] & b[91])^(a[264] & b[92])^(a[263] & b[93])^(a[262] & b[94])^(a[261] & b[95])^(a[260] & b[96])^(a[259] & b[97])^(a[258] & b[98])^(a[257] & b[99])^(a[256] & b[100])^(a[255] & b[101])^(a[254] & b[102])^(a[253] & b[103])^(a[252] & b[104])^(a[251] & b[105])^(a[250] & b[106])^(a[249] & b[107])^(a[248] & b[108])^(a[247] & b[109])^(a[246] & b[110])^(a[245] & b[111])^(a[244] & b[112])^(a[243] & b[113])^(a[242] & b[114])^(a[241] & b[115])^(a[240] & b[116])^(a[239] & b[117])^(a[238] & b[118])^(a[237] & b[119])^(a[236] & b[120])^(a[235] & b[121])^(a[234] & b[122])^(a[233] & b[123])^(a[232] & b[124])^(a[231] & b[125])^(a[230] & b[126])^(a[229] & b[127])^(a[228] & b[128])^(a[227] & b[129])^(a[226] & b[130])^(a[225] & b[131])^(a[224] & b[132])^(a[223] & b[133])^(a[222] & b[134])^(a[221] & b[135])^(a[220] & b[136])^(a[219] & b[137])^(a[218] & b[138])^(a[217] & b[139])^(a[216] & b[140])^(a[215] & b[141])^(a[214] & b[142])^(a[213] & b[143])^(a[212] & b[144])^(a[211] & b[145])^(a[210] & b[146])^(a[209] & b[147])^(a[208] & b[148])^(a[207] & b[149])^(a[206] & b[150])^(a[205] & b[151])^(a[204] & b[152])^(a[203] & b[153])^(a[202] & b[154])^(a[201] & b[155])^(a[200] & b[156])^(a[199] & b[157])^(a[198] & b[158])^(a[197] & b[159])^(a[196] & b[160])^(a[195] & b[161])^(a[194] & b[162])^(a[193] & b[163])^(a[192] & b[164])^(a[191] & b[165])^(a[190] & b[166])^(a[189] & b[167])^(a[188] & b[168])^(a[187] & b[169])^(a[186] & b[170])^(a[185] & b[171])^(a[184] & b[172])^(a[183] & b[173])^(a[182] & b[174])^(a[181] & b[175])^(a[180] & b[176])^(a[179] & b[177])^(a[178] & b[178])^(a[177] & b[179])^(a[176] & b[180])^(a[175] & b[181])^(a[174] & b[182])^(a[173] & b[183])^(a[172] & b[184])^(a[171] & b[185])^(a[170] & b[186])^(a[169] & b[187])^(a[168] & b[188])^(a[167] & b[189])^(a[166] & b[190])^(a[165] & b[191])^(a[164] & b[192])^(a[163] & b[193])^(a[162] & b[194])^(a[161] & b[195])^(a[160] & b[196])^(a[159] & b[197])^(a[158] & b[198])^(a[157] & b[199])^(a[156] & b[200])^(a[155] & b[201])^(a[154] & b[202])^(a[153] & b[203])^(a[152] & b[204])^(a[151] & b[205])^(a[150] & b[206])^(a[149] & b[207])^(a[148] & b[208])^(a[147] & b[209])^(a[146] & b[210])^(a[145] & b[211])^(a[144] & b[212])^(a[143] & b[213])^(a[142] & b[214])^(a[141] & b[215])^(a[140] & b[216])^(a[139] & b[217])^(a[138] & b[218])^(a[137] & b[219])^(a[136] & b[220])^(a[135] & b[221])^(a[134] & b[222])^(a[133] & b[223])^(a[132] & b[224])^(a[131] & b[225])^(a[130] & b[226])^(a[129] & b[227])^(a[128] & b[228])^(a[127] & b[229])^(a[126] & b[230])^(a[125] & b[231])^(a[124] & b[232])^(a[123] & b[233])^(a[122] & b[234])^(a[121] & b[235])^(a[120] & b[236])^(a[119] & b[237])^(a[118] & b[238])^(a[117] & b[239])^(a[116] & b[240])^(a[115] & b[241])^(a[114] & b[242])^(a[113] & b[243])^(a[112] & b[244])^(a[111] & b[245])^(a[110] & b[246])^(a[109] & b[247])^(a[108] & b[248])^(a[107] & b[249])^(a[106] & b[250])^(a[105] & b[251])^(a[104] & b[252])^(a[103] & b[253])^(a[102] & b[254])^(a[101] & b[255])^(a[100] & b[256])^(a[99] & b[257])^(a[98] & b[258])^(a[97] & b[259])^(a[96] & b[260])^(a[95] & b[261])^(a[94] & b[262])^(a[93] & b[263])^(a[92] & b[264])^(a[91] & b[265])^(a[90] & b[266])^(a[89] & b[267])^(a[88] & b[268])^(a[87] & b[269])^(a[86] & b[270])^(a[85] & b[271])^(a[84] & b[272])^(a[83] & b[273])^(a[82] & b[274])^(a[81] & b[275])^(a[80] & b[276])^(a[79] & b[277])^(a[78] & b[278])^(a[77] & b[279])^(a[76] & b[280])^(a[75] & b[281])^(a[74] & b[282])^(a[73] & b[283])^(a[72] & b[284])^(a[71] & b[285])^(a[70] & b[286])^(a[69] & b[287])^(a[68] & b[288])^(a[67] & b[289])^(a[66] & b[290])^(a[65] & b[291])^(a[64] & b[292])^(a[63] & b[293])^(a[62] & b[294])^(a[61] & b[295])^(a[60] & b[296])^(a[59] & b[297])^(a[58] & b[298])^(a[57] & b[299])^(a[56] & b[300])^(a[55] & b[301])^(a[54] & b[302])^(a[53] & b[303])^(a[52] & b[304])^(a[51] & b[305])^(a[50] & b[306])^(a[49] & b[307])^(a[48] & b[308])^(a[47] & b[309])^(a[46] & b[310])^(a[45] & b[311])^(a[44] & b[312])^(a[43] & b[313])^(a[42] & b[314])^(a[41] & b[315])^(a[40] & b[316])^(a[39] & b[317])^(a[38] & b[318])^(a[37] & b[319])^(a[36] & b[320])^(a[35] & b[321])^(a[34] & b[322])^(a[33] & b[323])^(a[32] & b[324])^(a[31] & b[325])^(a[30] & b[326])^(a[29] & b[327])^(a[28] & b[328])^(a[27] & b[329])^(a[26] & b[330])^(a[25] & b[331])^(a[24] & b[332])^(a[23] & b[333])^(a[22] & b[334])^(a[21] & b[335])^(a[20] & b[336])^(a[19] & b[337])^(a[18] & b[338])^(a[17] & b[339])^(a[16] & b[340])^(a[15] & b[341])^(a[14] & b[342])^(a[13] & b[343])^(a[12] & b[344])^(a[11] & b[345])^(a[10] & b[346])^(a[9] & b[347])^(a[8] & b[348])^(a[7] & b[349])^(a[6] & b[350])^(a[5] & b[351])^(a[4] & b[352])^(a[3] & b[353])^(a[2] & b[354])^(a[1] & b[355])^(a[0] & b[356]);
assign y[357] = (a[357] & b[0])^(a[356] & b[1])^(a[355] & b[2])^(a[354] & b[3])^(a[353] & b[4])^(a[352] & b[5])^(a[351] & b[6])^(a[350] & b[7])^(a[349] & b[8])^(a[348] & b[9])^(a[347] & b[10])^(a[346] & b[11])^(a[345] & b[12])^(a[344] & b[13])^(a[343] & b[14])^(a[342] & b[15])^(a[341] & b[16])^(a[340] & b[17])^(a[339] & b[18])^(a[338] & b[19])^(a[337] & b[20])^(a[336] & b[21])^(a[335] & b[22])^(a[334] & b[23])^(a[333] & b[24])^(a[332] & b[25])^(a[331] & b[26])^(a[330] & b[27])^(a[329] & b[28])^(a[328] & b[29])^(a[327] & b[30])^(a[326] & b[31])^(a[325] & b[32])^(a[324] & b[33])^(a[323] & b[34])^(a[322] & b[35])^(a[321] & b[36])^(a[320] & b[37])^(a[319] & b[38])^(a[318] & b[39])^(a[317] & b[40])^(a[316] & b[41])^(a[315] & b[42])^(a[314] & b[43])^(a[313] & b[44])^(a[312] & b[45])^(a[311] & b[46])^(a[310] & b[47])^(a[309] & b[48])^(a[308] & b[49])^(a[307] & b[50])^(a[306] & b[51])^(a[305] & b[52])^(a[304] & b[53])^(a[303] & b[54])^(a[302] & b[55])^(a[301] & b[56])^(a[300] & b[57])^(a[299] & b[58])^(a[298] & b[59])^(a[297] & b[60])^(a[296] & b[61])^(a[295] & b[62])^(a[294] & b[63])^(a[293] & b[64])^(a[292] & b[65])^(a[291] & b[66])^(a[290] & b[67])^(a[289] & b[68])^(a[288] & b[69])^(a[287] & b[70])^(a[286] & b[71])^(a[285] & b[72])^(a[284] & b[73])^(a[283] & b[74])^(a[282] & b[75])^(a[281] & b[76])^(a[280] & b[77])^(a[279] & b[78])^(a[278] & b[79])^(a[277] & b[80])^(a[276] & b[81])^(a[275] & b[82])^(a[274] & b[83])^(a[273] & b[84])^(a[272] & b[85])^(a[271] & b[86])^(a[270] & b[87])^(a[269] & b[88])^(a[268] & b[89])^(a[267] & b[90])^(a[266] & b[91])^(a[265] & b[92])^(a[264] & b[93])^(a[263] & b[94])^(a[262] & b[95])^(a[261] & b[96])^(a[260] & b[97])^(a[259] & b[98])^(a[258] & b[99])^(a[257] & b[100])^(a[256] & b[101])^(a[255] & b[102])^(a[254] & b[103])^(a[253] & b[104])^(a[252] & b[105])^(a[251] & b[106])^(a[250] & b[107])^(a[249] & b[108])^(a[248] & b[109])^(a[247] & b[110])^(a[246] & b[111])^(a[245] & b[112])^(a[244] & b[113])^(a[243] & b[114])^(a[242] & b[115])^(a[241] & b[116])^(a[240] & b[117])^(a[239] & b[118])^(a[238] & b[119])^(a[237] & b[120])^(a[236] & b[121])^(a[235] & b[122])^(a[234] & b[123])^(a[233] & b[124])^(a[232] & b[125])^(a[231] & b[126])^(a[230] & b[127])^(a[229] & b[128])^(a[228] & b[129])^(a[227] & b[130])^(a[226] & b[131])^(a[225] & b[132])^(a[224] & b[133])^(a[223] & b[134])^(a[222] & b[135])^(a[221] & b[136])^(a[220] & b[137])^(a[219] & b[138])^(a[218] & b[139])^(a[217] & b[140])^(a[216] & b[141])^(a[215] & b[142])^(a[214] & b[143])^(a[213] & b[144])^(a[212] & b[145])^(a[211] & b[146])^(a[210] & b[147])^(a[209] & b[148])^(a[208] & b[149])^(a[207] & b[150])^(a[206] & b[151])^(a[205] & b[152])^(a[204] & b[153])^(a[203] & b[154])^(a[202] & b[155])^(a[201] & b[156])^(a[200] & b[157])^(a[199] & b[158])^(a[198] & b[159])^(a[197] & b[160])^(a[196] & b[161])^(a[195] & b[162])^(a[194] & b[163])^(a[193] & b[164])^(a[192] & b[165])^(a[191] & b[166])^(a[190] & b[167])^(a[189] & b[168])^(a[188] & b[169])^(a[187] & b[170])^(a[186] & b[171])^(a[185] & b[172])^(a[184] & b[173])^(a[183] & b[174])^(a[182] & b[175])^(a[181] & b[176])^(a[180] & b[177])^(a[179] & b[178])^(a[178] & b[179])^(a[177] & b[180])^(a[176] & b[181])^(a[175] & b[182])^(a[174] & b[183])^(a[173] & b[184])^(a[172] & b[185])^(a[171] & b[186])^(a[170] & b[187])^(a[169] & b[188])^(a[168] & b[189])^(a[167] & b[190])^(a[166] & b[191])^(a[165] & b[192])^(a[164] & b[193])^(a[163] & b[194])^(a[162] & b[195])^(a[161] & b[196])^(a[160] & b[197])^(a[159] & b[198])^(a[158] & b[199])^(a[157] & b[200])^(a[156] & b[201])^(a[155] & b[202])^(a[154] & b[203])^(a[153] & b[204])^(a[152] & b[205])^(a[151] & b[206])^(a[150] & b[207])^(a[149] & b[208])^(a[148] & b[209])^(a[147] & b[210])^(a[146] & b[211])^(a[145] & b[212])^(a[144] & b[213])^(a[143] & b[214])^(a[142] & b[215])^(a[141] & b[216])^(a[140] & b[217])^(a[139] & b[218])^(a[138] & b[219])^(a[137] & b[220])^(a[136] & b[221])^(a[135] & b[222])^(a[134] & b[223])^(a[133] & b[224])^(a[132] & b[225])^(a[131] & b[226])^(a[130] & b[227])^(a[129] & b[228])^(a[128] & b[229])^(a[127] & b[230])^(a[126] & b[231])^(a[125] & b[232])^(a[124] & b[233])^(a[123] & b[234])^(a[122] & b[235])^(a[121] & b[236])^(a[120] & b[237])^(a[119] & b[238])^(a[118] & b[239])^(a[117] & b[240])^(a[116] & b[241])^(a[115] & b[242])^(a[114] & b[243])^(a[113] & b[244])^(a[112] & b[245])^(a[111] & b[246])^(a[110] & b[247])^(a[109] & b[248])^(a[108] & b[249])^(a[107] & b[250])^(a[106] & b[251])^(a[105] & b[252])^(a[104] & b[253])^(a[103] & b[254])^(a[102] & b[255])^(a[101] & b[256])^(a[100] & b[257])^(a[99] & b[258])^(a[98] & b[259])^(a[97] & b[260])^(a[96] & b[261])^(a[95] & b[262])^(a[94] & b[263])^(a[93] & b[264])^(a[92] & b[265])^(a[91] & b[266])^(a[90] & b[267])^(a[89] & b[268])^(a[88] & b[269])^(a[87] & b[270])^(a[86] & b[271])^(a[85] & b[272])^(a[84] & b[273])^(a[83] & b[274])^(a[82] & b[275])^(a[81] & b[276])^(a[80] & b[277])^(a[79] & b[278])^(a[78] & b[279])^(a[77] & b[280])^(a[76] & b[281])^(a[75] & b[282])^(a[74] & b[283])^(a[73] & b[284])^(a[72] & b[285])^(a[71] & b[286])^(a[70] & b[287])^(a[69] & b[288])^(a[68] & b[289])^(a[67] & b[290])^(a[66] & b[291])^(a[65] & b[292])^(a[64] & b[293])^(a[63] & b[294])^(a[62] & b[295])^(a[61] & b[296])^(a[60] & b[297])^(a[59] & b[298])^(a[58] & b[299])^(a[57] & b[300])^(a[56] & b[301])^(a[55] & b[302])^(a[54] & b[303])^(a[53] & b[304])^(a[52] & b[305])^(a[51] & b[306])^(a[50] & b[307])^(a[49] & b[308])^(a[48] & b[309])^(a[47] & b[310])^(a[46] & b[311])^(a[45] & b[312])^(a[44] & b[313])^(a[43] & b[314])^(a[42] & b[315])^(a[41] & b[316])^(a[40] & b[317])^(a[39] & b[318])^(a[38] & b[319])^(a[37] & b[320])^(a[36] & b[321])^(a[35] & b[322])^(a[34] & b[323])^(a[33] & b[324])^(a[32] & b[325])^(a[31] & b[326])^(a[30] & b[327])^(a[29] & b[328])^(a[28] & b[329])^(a[27] & b[330])^(a[26] & b[331])^(a[25] & b[332])^(a[24] & b[333])^(a[23] & b[334])^(a[22] & b[335])^(a[21] & b[336])^(a[20] & b[337])^(a[19] & b[338])^(a[18] & b[339])^(a[17] & b[340])^(a[16] & b[341])^(a[15] & b[342])^(a[14] & b[343])^(a[13] & b[344])^(a[12] & b[345])^(a[11] & b[346])^(a[10] & b[347])^(a[9] & b[348])^(a[8] & b[349])^(a[7] & b[350])^(a[6] & b[351])^(a[5] & b[352])^(a[4] & b[353])^(a[3] & b[354])^(a[2] & b[355])^(a[1] & b[356])^(a[0] & b[357]);
assign y[358] = (a[358] & b[0])^(a[357] & b[1])^(a[356] & b[2])^(a[355] & b[3])^(a[354] & b[4])^(a[353] & b[5])^(a[352] & b[6])^(a[351] & b[7])^(a[350] & b[8])^(a[349] & b[9])^(a[348] & b[10])^(a[347] & b[11])^(a[346] & b[12])^(a[345] & b[13])^(a[344] & b[14])^(a[343] & b[15])^(a[342] & b[16])^(a[341] & b[17])^(a[340] & b[18])^(a[339] & b[19])^(a[338] & b[20])^(a[337] & b[21])^(a[336] & b[22])^(a[335] & b[23])^(a[334] & b[24])^(a[333] & b[25])^(a[332] & b[26])^(a[331] & b[27])^(a[330] & b[28])^(a[329] & b[29])^(a[328] & b[30])^(a[327] & b[31])^(a[326] & b[32])^(a[325] & b[33])^(a[324] & b[34])^(a[323] & b[35])^(a[322] & b[36])^(a[321] & b[37])^(a[320] & b[38])^(a[319] & b[39])^(a[318] & b[40])^(a[317] & b[41])^(a[316] & b[42])^(a[315] & b[43])^(a[314] & b[44])^(a[313] & b[45])^(a[312] & b[46])^(a[311] & b[47])^(a[310] & b[48])^(a[309] & b[49])^(a[308] & b[50])^(a[307] & b[51])^(a[306] & b[52])^(a[305] & b[53])^(a[304] & b[54])^(a[303] & b[55])^(a[302] & b[56])^(a[301] & b[57])^(a[300] & b[58])^(a[299] & b[59])^(a[298] & b[60])^(a[297] & b[61])^(a[296] & b[62])^(a[295] & b[63])^(a[294] & b[64])^(a[293] & b[65])^(a[292] & b[66])^(a[291] & b[67])^(a[290] & b[68])^(a[289] & b[69])^(a[288] & b[70])^(a[287] & b[71])^(a[286] & b[72])^(a[285] & b[73])^(a[284] & b[74])^(a[283] & b[75])^(a[282] & b[76])^(a[281] & b[77])^(a[280] & b[78])^(a[279] & b[79])^(a[278] & b[80])^(a[277] & b[81])^(a[276] & b[82])^(a[275] & b[83])^(a[274] & b[84])^(a[273] & b[85])^(a[272] & b[86])^(a[271] & b[87])^(a[270] & b[88])^(a[269] & b[89])^(a[268] & b[90])^(a[267] & b[91])^(a[266] & b[92])^(a[265] & b[93])^(a[264] & b[94])^(a[263] & b[95])^(a[262] & b[96])^(a[261] & b[97])^(a[260] & b[98])^(a[259] & b[99])^(a[258] & b[100])^(a[257] & b[101])^(a[256] & b[102])^(a[255] & b[103])^(a[254] & b[104])^(a[253] & b[105])^(a[252] & b[106])^(a[251] & b[107])^(a[250] & b[108])^(a[249] & b[109])^(a[248] & b[110])^(a[247] & b[111])^(a[246] & b[112])^(a[245] & b[113])^(a[244] & b[114])^(a[243] & b[115])^(a[242] & b[116])^(a[241] & b[117])^(a[240] & b[118])^(a[239] & b[119])^(a[238] & b[120])^(a[237] & b[121])^(a[236] & b[122])^(a[235] & b[123])^(a[234] & b[124])^(a[233] & b[125])^(a[232] & b[126])^(a[231] & b[127])^(a[230] & b[128])^(a[229] & b[129])^(a[228] & b[130])^(a[227] & b[131])^(a[226] & b[132])^(a[225] & b[133])^(a[224] & b[134])^(a[223] & b[135])^(a[222] & b[136])^(a[221] & b[137])^(a[220] & b[138])^(a[219] & b[139])^(a[218] & b[140])^(a[217] & b[141])^(a[216] & b[142])^(a[215] & b[143])^(a[214] & b[144])^(a[213] & b[145])^(a[212] & b[146])^(a[211] & b[147])^(a[210] & b[148])^(a[209] & b[149])^(a[208] & b[150])^(a[207] & b[151])^(a[206] & b[152])^(a[205] & b[153])^(a[204] & b[154])^(a[203] & b[155])^(a[202] & b[156])^(a[201] & b[157])^(a[200] & b[158])^(a[199] & b[159])^(a[198] & b[160])^(a[197] & b[161])^(a[196] & b[162])^(a[195] & b[163])^(a[194] & b[164])^(a[193] & b[165])^(a[192] & b[166])^(a[191] & b[167])^(a[190] & b[168])^(a[189] & b[169])^(a[188] & b[170])^(a[187] & b[171])^(a[186] & b[172])^(a[185] & b[173])^(a[184] & b[174])^(a[183] & b[175])^(a[182] & b[176])^(a[181] & b[177])^(a[180] & b[178])^(a[179] & b[179])^(a[178] & b[180])^(a[177] & b[181])^(a[176] & b[182])^(a[175] & b[183])^(a[174] & b[184])^(a[173] & b[185])^(a[172] & b[186])^(a[171] & b[187])^(a[170] & b[188])^(a[169] & b[189])^(a[168] & b[190])^(a[167] & b[191])^(a[166] & b[192])^(a[165] & b[193])^(a[164] & b[194])^(a[163] & b[195])^(a[162] & b[196])^(a[161] & b[197])^(a[160] & b[198])^(a[159] & b[199])^(a[158] & b[200])^(a[157] & b[201])^(a[156] & b[202])^(a[155] & b[203])^(a[154] & b[204])^(a[153] & b[205])^(a[152] & b[206])^(a[151] & b[207])^(a[150] & b[208])^(a[149] & b[209])^(a[148] & b[210])^(a[147] & b[211])^(a[146] & b[212])^(a[145] & b[213])^(a[144] & b[214])^(a[143] & b[215])^(a[142] & b[216])^(a[141] & b[217])^(a[140] & b[218])^(a[139] & b[219])^(a[138] & b[220])^(a[137] & b[221])^(a[136] & b[222])^(a[135] & b[223])^(a[134] & b[224])^(a[133] & b[225])^(a[132] & b[226])^(a[131] & b[227])^(a[130] & b[228])^(a[129] & b[229])^(a[128] & b[230])^(a[127] & b[231])^(a[126] & b[232])^(a[125] & b[233])^(a[124] & b[234])^(a[123] & b[235])^(a[122] & b[236])^(a[121] & b[237])^(a[120] & b[238])^(a[119] & b[239])^(a[118] & b[240])^(a[117] & b[241])^(a[116] & b[242])^(a[115] & b[243])^(a[114] & b[244])^(a[113] & b[245])^(a[112] & b[246])^(a[111] & b[247])^(a[110] & b[248])^(a[109] & b[249])^(a[108] & b[250])^(a[107] & b[251])^(a[106] & b[252])^(a[105] & b[253])^(a[104] & b[254])^(a[103] & b[255])^(a[102] & b[256])^(a[101] & b[257])^(a[100] & b[258])^(a[99] & b[259])^(a[98] & b[260])^(a[97] & b[261])^(a[96] & b[262])^(a[95] & b[263])^(a[94] & b[264])^(a[93] & b[265])^(a[92] & b[266])^(a[91] & b[267])^(a[90] & b[268])^(a[89] & b[269])^(a[88] & b[270])^(a[87] & b[271])^(a[86] & b[272])^(a[85] & b[273])^(a[84] & b[274])^(a[83] & b[275])^(a[82] & b[276])^(a[81] & b[277])^(a[80] & b[278])^(a[79] & b[279])^(a[78] & b[280])^(a[77] & b[281])^(a[76] & b[282])^(a[75] & b[283])^(a[74] & b[284])^(a[73] & b[285])^(a[72] & b[286])^(a[71] & b[287])^(a[70] & b[288])^(a[69] & b[289])^(a[68] & b[290])^(a[67] & b[291])^(a[66] & b[292])^(a[65] & b[293])^(a[64] & b[294])^(a[63] & b[295])^(a[62] & b[296])^(a[61] & b[297])^(a[60] & b[298])^(a[59] & b[299])^(a[58] & b[300])^(a[57] & b[301])^(a[56] & b[302])^(a[55] & b[303])^(a[54] & b[304])^(a[53] & b[305])^(a[52] & b[306])^(a[51] & b[307])^(a[50] & b[308])^(a[49] & b[309])^(a[48] & b[310])^(a[47] & b[311])^(a[46] & b[312])^(a[45] & b[313])^(a[44] & b[314])^(a[43] & b[315])^(a[42] & b[316])^(a[41] & b[317])^(a[40] & b[318])^(a[39] & b[319])^(a[38] & b[320])^(a[37] & b[321])^(a[36] & b[322])^(a[35] & b[323])^(a[34] & b[324])^(a[33] & b[325])^(a[32] & b[326])^(a[31] & b[327])^(a[30] & b[328])^(a[29] & b[329])^(a[28] & b[330])^(a[27] & b[331])^(a[26] & b[332])^(a[25] & b[333])^(a[24] & b[334])^(a[23] & b[335])^(a[22] & b[336])^(a[21] & b[337])^(a[20] & b[338])^(a[19] & b[339])^(a[18] & b[340])^(a[17] & b[341])^(a[16] & b[342])^(a[15] & b[343])^(a[14] & b[344])^(a[13] & b[345])^(a[12] & b[346])^(a[11] & b[347])^(a[10] & b[348])^(a[9] & b[349])^(a[8] & b[350])^(a[7] & b[351])^(a[6] & b[352])^(a[5] & b[353])^(a[4] & b[354])^(a[3] & b[355])^(a[2] & b[356])^(a[1] & b[357])^(a[0] & b[358]);
assign y[359] = (a[359] & b[0])^(a[358] & b[1])^(a[357] & b[2])^(a[356] & b[3])^(a[355] & b[4])^(a[354] & b[5])^(a[353] & b[6])^(a[352] & b[7])^(a[351] & b[8])^(a[350] & b[9])^(a[349] & b[10])^(a[348] & b[11])^(a[347] & b[12])^(a[346] & b[13])^(a[345] & b[14])^(a[344] & b[15])^(a[343] & b[16])^(a[342] & b[17])^(a[341] & b[18])^(a[340] & b[19])^(a[339] & b[20])^(a[338] & b[21])^(a[337] & b[22])^(a[336] & b[23])^(a[335] & b[24])^(a[334] & b[25])^(a[333] & b[26])^(a[332] & b[27])^(a[331] & b[28])^(a[330] & b[29])^(a[329] & b[30])^(a[328] & b[31])^(a[327] & b[32])^(a[326] & b[33])^(a[325] & b[34])^(a[324] & b[35])^(a[323] & b[36])^(a[322] & b[37])^(a[321] & b[38])^(a[320] & b[39])^(a[319] & b[40])^(a[318] & b[41])^(a[317] & b[42])^(a[316] & b[43])^(a[315] & b[44])^(a[314] & b[45])^(a[313] & b[46])^(a[312] & b[47])^(a[311] & b[48])^(a[310] & b[49])^(a[309] & b[50])^(a[308] & b[51])^(a[307] & b[52])^(a[306] & b[53])^(a[305] & b[54])^(a[304] & b[55])^(a[303] & b[56])^(a[302] & b[57])^(a[301] & b[58])^(a[300] & b[59])^(a[299] & b[60])^(a[298] & b[61])^(a[297] & b[62])^(a[296] & b[63])^(a[295] & b[64])^(a[294] & b[65])^(a[293] & b[66])^(a[292] & b[67])^(a[291] & b[68])^(a[290] & b[69])^(a[289] & b[70])^(a[288] & b[71])^(a[287] & b[72])^(a[286] & b[73])^(a[285] & b[74])^(a[284] & b[75])^(a[283] & b[76])^(a[282] & b[77])^(a[281] & b[78])^(a[280] & b[79])^(a[279] & b[80])^(a[278] & b[81])^(a[277] & b[82])^(a[276] & b[83])^(a[275] & b[84])^(a[274] & b[85])^(a[273] & b[86])^(a[272] & b[87])^(a[271] & b[88])^(a[270] & b[89])^(a[269] & b[90])^(a[268] & b[91])^(a[267] & b[92])^(a[266] & b[93])^(a[265] & b[94])^(a[264] & b[95])^(a[263] & b[96])^(a[262] & b[97])^(a[261] & b[98])^(a[260] & b[99])^(a[259] & b[100])^(a[258] & b[101])^(a[257] & b[102])^(a[256] & b[103])^(a[255] & b[104])^(a[254] & b[105])^(a[253] & b[106])^(a[252] & b[107])^(a[251] & b[108])^(a[250] & b[109])^(a[249] & b[110])^(a[248] & b[111])^(a[247] & b[112])^(a[246] & b[113])^(a[245] & b[114])^(a[244] & b[115])^(a[243] & b[116])^(a[242] & b[117])^(a[241] & b[118])^(a[240] & b[119])^(a[239] & b[120])^(a[238] & b[121])^(a[237] & b[122])^(a[236] & b[123])^(a[235] & b[124])^(a[234] & b[125])^(a[233] & b[126])^(a[232] & b[127])^(a[231] & b[128])^(a[230] & b[129])^(a[229] & b[130])^(a[228] & b[131])^(a[227] & b[132])^(a[226] & b[133])^(a[225] & b[134])^(a[224] & b[135])^(a[223] & b[136])^(a[222] & b[137])^(a[221] & b[138])^(a[220] & b[139])^(a[219] & b[140])^(a[218] & b[141])^(a[217] & b[142])^(a[216] & b[143])^(a[215] & b[144])^(a[214] & b[145])^(a[213] & b[146])^(a[212] & b[147])^(a[211] & b[148])^(a[210] & b[149])^(a[209] & b[150])^(a[208] & b[151])^(a[207] & b[152])^(a[206] & b[153])^(a[205] & b[154])^(a[204] & b[155])^(a[203] & b[156])^(a[202] & b[157])^(a[201] & b[158])^(a[200] & b[159])^(a[199] & b[160])^(a[198] & b[161])^(a[197] & b[162])^(a[196] & b[163])^(a[195] & b[164])^(a[194] & b[165])^(a[193] & b[166])^(a[192] & b[167])^(a[191] & b[168])^(a[190] & b[169])^(a[189] & b[170])^(a[188] & b[171])^(a[187] & b[172])^(a[186] & b[173])^(a[185] & b[174])^(a[184] & b[175])^(a[183] & b[176])^(a[182] & b[177])^(a[181] & b[178])^(a[180] & b[179])^(a[179] & b[180])^(a[178] & b[181])^(a[177] & b[182])^(a[176] & b[183])^(a[175] & b[184])^(a[174] & b[185])^(a[173] & b[186])^(a[172] & b[187])^(a[171] & b[188])^(a[170] & b[189])^(a[169] & b[190])^(a[168] & b[191])^(a[167] & b[192])^(a[166] & b[193])^(a[165] & b[194])^(a[164] & b[195])^(a[163] & b[196])^(a[162] & b[197])^(a[161] & b[198])^(a[160] & b[199])^(a[159] & b[200])^(a[158] & b[201])^(a[157] & b[202])^(a[156] & b[203])^(a[155] & b[204])^(a[154] & b[205])^(a[153] & b[206])^(a[152] & b[207])^(a[151] & b[208])^(a[150] & b[209])^(a[149] & b[210])^(a[148] & b[211])^(a[147] & b[212])^(a[146] & b[213])^(a[145] & b[214])^(a[144] & b[215])^(a[143] & b[216])^(a[142] & b[217])^(a[141] & b[218])^(a[140] & b[219])^(a[139] & b[220])^(a[138] & b[221])^(a[137] & b[222])^(a[136] & b[223])^(a[135] & b[224])^(a[134] & b[225])^(a[133] & b[226])^(a[132] & b[227])^(a[131] & b[228])^(a[130] & b[229])^(a[129] & b[230])^(a[128] & b[231])^(a[127] & b[232])^(a[126] & b[233])^(a[125] & b[234])^(a[124] & b[235])^(a[123] & b[236])^(a[122] & b[237])^(a[121] & b[238])^(a[120] & b[239])^(a[119] & b[240])^(a[118] & b[241])^(a[117] & b[242])^(a[116] & b[243])^(a[115] & b[244])^(a[114] & b[245])^(a[113] & b[246])^(a[112] & b[247])^(a[111] & b[248])^(a[110] & b[249])^(a[109] & b[250])^(a[108] & b[251])^(a[107] & b[252])^(a[106] & b[253])^(a[105] & b[254])^(a[104] & b[255])^(a[103] & b[256])^(a[102] & b[257])^(a[101] & b[258])^(a[100] & b[259])^(a[99] & b[260])^(a[98] & b[261])^(a[97] & b[262])^(a[96] & b[263])^(a[95] & b[264])^(a[94] & b[265])^(a[93] & b[266])^(a[92] & b[267])^(a[91] & b[268])^(a[90] & b[269])^(a[89] & b[270])^(a[88] & b[271])^(a[87] & b[272])^(a[86] & b[273])^(a[85] & b[274])^(a[84] & b[275])^(a[83] & b[276])^(a[82] & b[277])^(a[81] & b[278])^(a[80] & b[279])^(a[79] & b[280])^(a[78] & b[281])^(a[77] & b[282])^(a[76] & b[283])^(a[75] & b[284])^(a[74] & b[285])^(a[73] & b[286])^(a[72] & b[287])^(a[71] & b[288])^(a[70] & b[289])^(a[69] & b[290])^(a[68] & b[291])^(a[67] & b[292])^(a[66] & b[293])^(a[65] & b[294])^(a[64] & b[295])^(a[63] & b[296])^(a[62] & b[297])^(a[61] & b[298])^(a[60] & b[299])^(a[59] & b[300])^(a[58] & b[301])^(a[57] & b[302])^(a[56] & b[303])^(a[55] & b[304])^(a[54] & b[305])^(a[53] & b[306])^(a[52] & b[307])^(a[51] & b[308])^(a[50] & b[309])^(a[49] & b[310])^(a[48] & b[311])^(a[47] & b[312])^(a[46] & b[313])^(a[45] & b[314])^(a[44] & b[315])^(a[43] & b[316])^(a[42] & b[317])^(a[41] & b[318])^(a[40] & b[319])^(a[39] & b[320])^(a[38] & b[321])^(a[37] & b[322])^(a[36] & b[323])^(a[35] & b[324])^(a[34] & b[325])^(a[33] & b[326])^(a[32] & b[327])^(a[31] & b[328])^(a[30] & b[329])^(a[29] & b[330])^(a[28] & b[331])^(a[27] & b[332])^(a[26] & b[333])^(a[25] & b[334])^(a[24] & b[335])^(a[23] & b[336])^(a[22] & b[337])^(a[21] & b[338])^(a[20] & b[339])^(a[19] & b[340])^(a[18] & b[341])^(a[17] & b[342])^(a[16] & b[343])^(a[15] & b[344])^(a[14] & b[345])^(a[13] & b[346])^(a[12] & b[347])^(a[11] & b[348])^(a[10] & b[349])^(a[9] & b[350])^(a[8] & b[351])^(a[7] & b[352])^(a[6] & b[353])^(a[5] & b[354])^(a[4] & b[355])^(a[3] & b[356])^(a[2] & b[357])^(a[1] & b[358])^(a[0] & b[359]);
assign y[360] = (a[360] & b[0])^(a[359] & b[1])^(a[358] & b[2])^(a[357] & b[3])^(a[356] & b[4])^(a[355] & b[5])^(a[354] & b[6])^(a[353] & b[7])^(a[352] & b[8])^(a[351] & b[9])^(a[350] & b[10])^(a[349] & b[11])^(a[348] & b[12])^(a[347] & b[13])^(a[346] & b[14])^(a[345] & b[15])^(a[344] & b[16])^(a[343] & b[17])^(a[342] & b[18])^(a[341] & b[19])^(a[340] & b[20])^(a[339] & b[21])^(a[338] & b[22])^(a[337] & b[23])^(a[336] & b[24])^(a[335] & b[25])^(a[334] & b[26])^(a[333] & b[27])^(a[332] & b[28])^(a[331] & b[29])^(a[330] & b[30])^(a[329] & b[31])^(a[328] & b[32])^(a[327] & b[33])^(a[326] & b[34])^(a[325] & b[35])^(a[324] & b[36])^(a[323] & b[37])^(a[322] & b[38])^(a[321] & b[39])^(a[320] & b[40])^(a[319] & b[41])^(a[318] & b[42])^(a[317] & b[43])^(a[316] & b[44])^(a[315] & b[45])^(a[314] & b[46])^(a[313] & b[47])^(a[312] & b[48])^(a[311] & b[49])^(a[310] & b[50])^(a[309] & b[51])^(a[308] & b[52])^(a[307] & b[53])^(a[306] & b[54])^(a[305] & b[55])^(a[304] & b[56])^(a[303] & b[57])^(a[302] & b[58])^(a[301] & b[59])^(a[300] & b[60])^(a[299] & b[61])^(a[298] & b[62])^(a[297] & b[63])^(a[296] & b[64])^(a[295] & b[65])^(a[294] & b[66])^(a[293] & b[67])^(a[292] & b[68])^(a[291] & b[69])^(a[290] & b[70])^(a[289] & b[71])^(a[288] & b[72])^(a[287] & b[73])^(a[286] & b[74])^(a[285] & b[75])^(a[284] & b[76])^(a[283] & b[77])^(a[282] & b[78])^(a[281] & b[79])^(a[280] & b[80])^(a[279] & b[81])^(a[278] & b[82])^(a[277] & b[83])^(a[276] & b[84])^(a[275] & b[85])^(a[274] & b[86])^(a[273] & b[87])^(a[272] & b[88])^(a[271] & b[89])^(a[270] & b[90])^(a[269] & b[91])^(a[268] & b[92])^(a[267] & b[93])^(a[266] & b[94])^(a[265] & b[95])^(a[264] & b[96])^(a[263] & b[97])^(a[262] & b[98])^(a[261] & b[99])^(a[260] & b[100])^(a[259] & b[101])^(a[258] & b[102])^(a[257] & b[103])^(a[256] & b[104])^(a[255] & b[105])^(a[254] & b[106])^(a[253] & b[107])^(a[252] & b[108])^(a[251] & b[109])^(a[250] & b[110])^(a[249] & b[111])^(a[248] & b[112])^(a[247] & b[113])^(a[246] & b[114])^(a[245] & b[115])^(a[244] & b[116])^(a[243] & b[117])^(a[242] & b[118])^(a[241] & b[119])^(a[240] & b[120])^(a[239] & b[121])^(a[238] & b[122])^(a[237] & b[123])^(a[236] & b[124])^(a[235] & b[125])^(a[234] & b[126])^(a[233] & b[127])^(a[232] & b[128])^(a[231] & b[129])^(a[230] & b[130])^(a[229] & b[131])^(a[228] & b[132])^(a[227] & b[133])^(a[226] & b[134])^(a[225] & b[135])^(a[224] & b[136])^(a[223] & b[137])^(a[222] & b[138])^(a[221] & b[139])^(a[220] & b[140])^(a[219] & b[141])^(a[218] & b[142])^(a[217] & b[143])^(a[216] & b[144])^(a[215] & b[145])^(a[214] & b[146])^(a[213] & b[147])^(a[212] & b[148])^(a[211] & b[149])^(a[210] & b[150])^(a[209] & b[151])^(a[208] & b[152])^(a[207] & b[153])^(a[206] & b[154])^(a[205] & b[155])^(a[204] & b[156])^(a[203] & b[157])^(a[202] & b[158])^(a[201] & b[159])^(a[200] & b[160])^(a[199] & b[161])^(a[198] & b[162])^(a[197] & b[163])^(a[196] & b[164])^(a[195] & b[165])^(a[194] & b[166])^(a[193] & b[167])^(a[192] & b[168])^(a[191] & b[169])^(a[190] & b[170])^(a[189] & b[171])^(a[188] & b[172])^(a[187] & b[173])^(a[186] & b[174])^(a[185] & b[175])^(a[184] & b[176])^(a[183] & b[177])^(a[182] & b[178])^(a[181] & b[179])^(a[180] & b[180])^(a[179] & b[181])^(a[178] & b[182])^(a[177] & b[183])^(a[176] & b[184])^(a[175] & b[185])^(a[174] & b[186])^(a[173] & b[187])^(a[172] & b[188])^(a[171] & b[189])^(a[170] & b[190])^(a[169] & b[191])^(a[168] & b[192])^(a[167] & b[193])^(a[166] & b[194])^(a[165] & b[195])^(a[164] & b[196])^(a[163] & b[197])^(a[162] & b[198])^(a[161] & b[199])^(a[160] & b[200])^(a[159] & b[201])^(a[158] & b[202])^(a[157] & b[203])^(a[156] & b[204])^(a[155] & b[205])^(a[154] & b[206])^(a[153] & b[207])^(a[152] & b[208])^(a[151] & b[209])^(a[150] & b[210])^(a[149] & b[211])^(a[148] & b[212])^(a[147] & b[213])^(a[146] & b[214])^(a[145] & b[215])^(a[144] & b[216])^(a[143] & b[217])^(a[142] & b[218])^(a[141] & b[219])^(a[140] & b[220])^(a[139] & b[221])^(a[138] & b[222])^(a[137] & b[223])^(a[136] & b[224])^(a[135] & b[225])^(a[134] & b[226])^(a[133] & b[227])^(a[132] & b[228])^(a[131] & b[229])^(a[130] & b[230])^(a[129] & b[231])^(a[128] & b[232])^(a[127] & b[233])^(a[126] & b[234])^(a[125] & b[235])^(a[124] & b[236])^(a[123] & b[237])^(a[122] & b[238])^(a[121] & b[239])^(a[120] & b[240])^(a[119] & b[241])^(a[118] & b[242])^(a[117] & b[243])^(a[116] & b[244])^(a[115] & b[245])^(a[114] & b[246])^(a[113] & b[247])^(a[112] & b[248])^(a[111] & b[249])^(a[110] & b[250])^(a[109] & b[251])^(a[108] & b[252])^(a[107] & b[253])^(a[106] & b[254])^(a[105] & b[255])^(a[104] & b[256])^(a[103] & b[257])^(a[102] & b[258])^(a[101] & b[259])^(a[100] & b[260])^(a[99] & b[261])^(a[98] & b[262])^(a[97] & b[263])^(a[96] & b[264])^(a[95] & b[265])^(a[94] & b[266])^(a[93] & b[267])^(a[92] & b[268])^(a[91] & b[269])^(a[90] & b[270])^(a[89] & b[271])^(a[88] & b[272])^(a[87] & b[273])^(a[86] & b[274])^(a[85] & b[275])^(a[84] & b[276])^(a[83] & b[277])^(a[82] & b[278])^(a[81] & b[279])^(a[80] & b[280])^(a[79] & b[281])^(a[78] & b[282])^(a[77] & b[283])^(a[76] & b[284])^(a[75] & b[285])^(a[74] & b[286])^(a[73] & b[287])^(a[72] & b[288])^(a[71] & b[289])^(a[70] & b[290])^(a[69] & b[291])^(a[68] & b[292])^(a[67] & b[293])^(a[66] & b[294])^(a[65] & b[295])^(a[64] & b[296])^(a[63] & b[297])^(a[62] & b[298])^(a[61] & b[299])^(a[60] & b[300])^(a[59] & b[301])^(a[58] & b[302])^(a[57] & b[303])^(a[56] & b[304])^(a[55] & b[305])^(a[54] & b[306])^(a[53] & b[307])^(a[52] & b[308])^(a[51] & b[309])^(a[50] & b[310])^(a[49] & b[311])^(a[48] & b[312])^(a[47] & b[313])^(a[46] & b[314])^(a[45] & b[315])^(a[44] & b[316])^(a[43] & b[317])^(a[42] & b[318])^(a[41] & b[319])^(a[40] & b[320])^(a[39] & b[321])^(a[38] & b[322])^(a[37] & b[323])^(a[36] & b[324])^(a[35] & b[325])^(a[34] & b[326])^(a[33] & b[327])^(a[32] & b[328])^(a[31] & b[329])^(a[30] & b[330])^(a[29] & b[331])^(a[28] & b[332])^(a[27] & b[333])^(a[26] & b[334])^(a[25] & b[335])^(a[24] & b[336])^(a[23] & b[337])^(a[22] & b[338])^(a[21] & b[339])^(a[20] & b[340])^(a[19] & b[341])^(a[18] & b[342])^(a[17] & b[343])^(a[16] & b[344])^(a[15] & b[345])^(a[14] & b[346])^(a[13] & b[347])^(a[12] & b[348])^(a[11] & b[349])^(a[10] & b[350])^(a[9] & b[351])^(a[8] & b[352])^(a[7] & b[353])^(a[6] & b[354])^(a[5] & b[355])^(a[4] & b[356])^(a[3] & b[357])^(a[2] & b[358])^(a[1] & b[359])^(a[0] & b[360]);
assign y[361] = (a[361] & b[0])^(a[360] & b[1])^(a[359] & b[2])^(a[358] & b[3])^(a[357] & b[4])^(a[356] & b[5])^(a[355] & b[6])^(a[354] & b[7])^(a[353] & b[8])^(a[352] & b[9])^(a[351] & b[10])^(a[350] & b[11])^(a[349] & b[12])^(a[348] & b[13])^(a[347] & b[14])^(a[346] & b[15])^(a[345] & b[16])^(a[344] & b[17])^(a[343] & b[18])^(a[342] & b[19])^(a[341] & b[20])^(a[340] & b[21])^(a[339] & b[22])^(a[338] & b[23])^(a[337] & b[24])^(a[336] & b[25])^(a[335] & b[26])^(a[334] & b[27])^(a[333] & b[28])^(a[332] & b[29])^(a[331] & b[30])^(a[330] & b[31])^(a[329] & b[32])^(a[328] & b[33])^(a[327] & b[34])^(a[326] & b[35])^(a[325] & b[36])^(a[324] & b[37])^(a[323] & b[38])^(a[322] & b[39])^(a[321] & b[40])^(a[320] & b[41])^(a[319] & b[42])^(a[318] & b[43])^(a[317] & b[44])^(a[316] & b[45])^(a[315] & b[46])^(a[314] & b[47])^(a[313] & b[48])^(a[312] & b[49])^(a[311] & b[50])^(a[310] & b[51])^(a[309] & b[52])^(a[308] & b[53])^(a[307] & b[54])^(a[306] & b[55])^(a[305] & b[56])^(a[304] & b[57])^(a[303] & b[58])^(a[302] & b[59])^(a[301] & b[60])^(a[300] & b[61])^(a[299] & b[62])^(a[298] & b[63])^(a[297] & b[64])^(a[296] & b[65])^(a[295] & b[66])^(a[294] & b[67])^(a[293] & b[68])^(a[292] & b[69])^(a[291] & b[70])^(a[290] & b[71])^(a[289] & b[72])^(a[288] & b[73])^(a[287] & b[74])^(a[286] & b[75])^(a[285] & b[76])^(a[284] & b[77])^(a[283] & b[78])^(a[282] & b[79])^(a[281] & b[80])^(a[280] & b[81])^(a[279] & b[82])^(a[278] & b[83])^(a[277] & b[84])^(a[276] & b[85])^(a[275] & b[86])^(a[274] & b[87])^(a[273] & b[88])^(a[272] & b[89])^(a[271] & b[90])^(a[270] & b[91])^(a[269] & b[92])^(a[268] & b[93])^(a[267] & b[94])^(a[266] & b[95])^(a[265] & b[96])^(a[264] & b[97])^(a[263] & b[98])^(a[262] & b[99])^(a[261] & b[100])^(a[260] & b[101])^(a[259] & b[102])^(a[258] & b[103])^(a[257] & b[104])^(a[256] & b[105])^(a[255] & b[106])^(a[254] & b[107])^(a[253] & b[108])^(a[252] & b[109])^(a[251] & b[110])^(a[250] & b[111])^(a[249] & b[112])^(a[248] & b[113])^(a[247] & b[114])^(a[246] & b[115])^(a[245] & b[116])^(a[244] & b[117])^(a[243] & b[118])^(a[242] & b[119])^(a[241] & b[120])^(a[240] & b[121])^(a[239] & b[122])^(a[238] & b[123])^(a[237] & b[124])^(a[236] & b[125])^(a[235] & b[126])^(a[234] & b[127])^(a[233] & b[128])^(a[232] & b[129])^(a[231] & b[130])^(a[230] & b[131])^(a[229] & b[132])^(a[228] & b[133])^(a[227] & b[134])^(a[226] & b[135])^(a[225] & b[136])^(a[224] & b[137])^(a[223] & b[138])^(a[222] & b[139])^(a[221] & b[140])^(a[220] & b[141])^(a[219] & b[142])^(a[218] & b[143])^(a[217] & b[144])^(a[216] & b[145])^(a[215] & b[146])^(a[214] & b[147])^(a[213] & b[148])^(a[212] & b[149])^(a[211] & b[150])^(a[210] & b[151])^(a[209] & b[152])^(a[208] & b[153])^(a[207] & b[154])^(a[206] & b[155])^(a[205] & b[156])^(a[204] & b[157])^(a[203] & b[158])^(a[202] & b[159])^(a[201] & b[160])^(a[200] & b[161])^(a[199] & b[162])^(a[198] & b[163])^(a[197] & b[164])^(a[196] & b[165])^(a[195] & b[166])^(a[194] & b[167])^(a[193] & b[168])^(a[192] & b[169])^(a[191] & b[170])^(a[190] & b[171])^(a[189] & b[172])^(a[188] & b[173])^(a[187] & b[174])^(a[186] & b[175])^(a[185] & b[176])^(a[184] & b[177])^(a[183] & b[178])^(a[182] & b[179])^(a[181] & b[180])^(a[180] & b[181])^(a[179] & b[182])^(a[178] & b[183])^(a[177] & b[184])^(a[176] & b[185])^(a[175] & b[186])^(a[174] & b[187])^(a[173] & b[188])^(a[172] & b[189])^(a[171] & b[190])^(a[170] & b[191])^(a[169] & b[192])^(a[168] & b[193])^(a[167] & b[194])^(a[166] & b[195])^(a[165] & b[196])^(a[164] & b[197])^(a[163] & b[198])^(a[162] & b[199])^(a[161] & b[200])^(a[160] & b[201])^(a[159] & b[202])^(a[158] & b[203])^(a[157] & b[204])^(a[156] & b[205])^(a[155] & b[206])^(a[154] & b[207])^(a[153] & b[208])^(a[152] & b[209])^(a[151] & b[210])^(a[150] & b[211])^(a[149] & b[212])^(a[148] & b[213])^(a[147] & b[214])^(a[146] & b[215])^(a[145] & b[216])^(a[144] & b[217])^(a[143] & b[218])^(a[142] & b[219])^(a[141] & b[220])^(a[140] & b[221])^(a[139] & b[222])^(a[138] & b[223])^(a[137] & b[224])^(a[136] & b[225])^(a[135] & b[226])^(a[134] & b[227])^(a[133] & b[228])^(a[132] & b[229])^(a[131] & b[230])^(a[130] & b[231])^(a[129] & b[232])^(a[128] & b[233])^(a[127] & b[234])^(a[126] & b[235])^(a[125] & b[236])^(a[124] & b[237])^(a[123] & b[238])^(a[122] & b[239])^(a[121] & b[240])^(a[120] & b[241])^(a[119] & b[242])^(a[118] & b[243])^(a[117] & b[244])^(a[116] & b[245])^(a[115] & b[246])^(a[114] & b[247])^(a[113] & b[248])^(a[112] & b[249])^(a[111] & b[250])^(a[110] & b[251])^(a[109] & b[252])^(a[108] & b[253])^(a[107] & b[254])^(a[106] & b[255])^(a[105] & b[256])^(a[104] & b[257])^(a[103] & b[258])^(a[102] & b[259])^(a[101] & b[260])^(a[100] & b[261])^(a[99] & b[262])^(a[98] & b[263])^(a[97] & b[264])^(a[96] & b[265])^(a[95] & b[266])^(a[94] & b[267])^(a[93] & b[268])^(a[92] & b[269])^(a[91] & b[270])^(a[90] & b[271])^(a[89] & b[272])^(a[88] & b[273])^(a[87] & b[274])^(a[86] & b[275])^(a[85] & b[276])^(a[84] & b[277])^(a[83] & b[278])^(a[82] & b[279])^(a[81] & b[280])^(a[80] & b[281])^(a[79] & b[282])^(a[78] & b[283])^(a[77] & b[284])^(a[76] & b[285])^(a[75] & b[286])^(a[74] & b[287])^(a[73] & b[288])^(a[72] & b[289])^(a[71] & b[290])^(a[70] & b[291])^(a[69] & b[292])^(a[68] & b[293])^(a[67] & b[294])^(a[66] & b[295])^(a[65] & b[296])^(a[64] & b[297])^(a[63] & b[298])^(a[62] & b[299])^(a[61] & b[300])^(a[60] & b[301])^(a[59] & b[302])^(a[58] & b[303])^(a[57] & b[304])^(a[56] & b[305])^(a[55] & b[306])^(a[54] & b[307])^(a[53] & b[308])^(a[52] & b[309])^(a[51] & b[310])^(a[50] & b[311])^(a[49] & b[312])^(a[48] & b[313])^(a[47] & b[314])^(a[46] & b[315])^(a[45] & b[316])^(a[44] & b[317])^(a[43] & b[318])^(a[42] & b[319])^(a[41] & b[320])^(a[40] & b[321])^(a[39] & b[322])^(a[38] & b[323])^(a[37] & b[324])^(a[36] & b[325])^(a[35] & b[326])^(a[34] & b[327])^(a[33] & b[328])^(a[32] & b[329])^(a[31] & b[330])^(a[30] & b[331])^(a[29] & b[332])^(a[28] & b[333])^(a[27] & b[334])^(a[26] & b[335])^(a[25] & b[336])^(a[24] & b[337])^(a[23] & b[338])^(a[22] & b[339])^(a[21] & b[340])^(a[20] & b[341])^(a[19] & b[342])^(a[18] & b[343])^(a[17] & b[344])^(a[16] & b[345])^(a[15] & b[346])^(a[14] & b[347])^(a[13] & b[348])^(a[12] & b[349])^(a[11] & b[350])^(a[10] & b[351])^(a[9] & b[352])^(a[8] & b[353])^(a[7] & b[354])^(a[6] & b[355])^(a[5] & b[356])^(a[4] & b[357])^(a[3] & b[358])^(a[2] & b[359])^(a[1] & b[360])^(a[0] & b[361]);
assign y[362] = (a[362] & b[0])^(a[361] & b[1])^(a[360] & b[2])^(a[359] & b[3])^(a[358] & b[4])^(a[357] & b[5])^(a[356] & b[6])^(a[355] & b[7])^(a[354] & b[8])^(a[353] & b[9])^(a[352] & b[10])^(a[351] & b[11])^(a[350] & b[12])^(a[349] & b[13])^(a[348] & b[14])^(a[347] & b[15])^(a[346] & b[16])^(a[345] & b[17])^(a[344] & b[18])^(a[343] & b[19])^(a[342] & b[20])^(a[341] & b[21])^(a[340] & b[22])^(a[339] & b[23])^(a[338] & b[24])^(a[337] & b[25])^(a[336] & b[26])^(a[335] & b[27])^(a[334] & b[28])^(a[333] & b[29])^(a[332] & b[30])^(a[331] & b[31])^(a[330] & b[32])^(a[329] & b[33])^(a[328] & b[34])^(a[327] & b[35])^(a[326] & b[36])^(a[325] & b[37])^(a[324] & b[38])^(a[323] & b[39])^(a[322] & b[40])^(a[321] & b[41])^(a[320] & b[42])^(a[319] & b[43])^(a[318] & b[44])^(a[317] & b[45])^(a[316] & b[46])^(a[315] & b[47])^(a[314] & b[48])^(a[313] & b[49])^(a[312] & b[50])^(a[311] & b[51])^(a[310] & b[52])^(a[309] & b[53])^(a[308] & b[54])^(a[307] & b[55])^(a[306] & b[56])^(a[305] & b[57])^(a[304] & b[58])^(a[303] & b[59])^(a[302] & b[60])^(a[301] & b[61])^(a[300] & b[62])^(a[299] & b[63])^(a[298] & b[64])^(a[297] & b[65])^(a[296] & b[66])^(a[295] & b[67])^(a[294] & b[68])^(a[293] & b[69])^(a[292] & b[70])^(a[291] & b[71])^(a[290] & b[72])^(a[289] & b[73])^(a[288] & b[74])^(a[287] & b[75])^(a[286] & b[76])^(a[285] & b[77])^(a[284] & b[78])^(a[283] & b[79])^(a[282] & b[80])^(a[281] & b[81])^(a[280] & b[82])^(a[279] & b[83])^(a[278] & b[84])^(a[277] & b[85])^(a[276] & b[86])^(a[275] & b[87])^(a[274] & b[88])^(a[273] & b[89])^(a[272] & b[90])^(a[271] & b[91])^(a[270] & b[92])^(a[269] & b[93])^(a[268] & b[94])^(a[267] & b[95])^(a[266] & b[96])^(a[265] & b[97])^(a[264] & b[98])^(a[263] & b[99])^(a[262] & b[100])^(a[261] & b[101])^(a[260] & b[102])^(a[259] & b[103])^(a[258] & b[104])^(a[257] & b[105])^(a[256] & b[106])^(a[255] & b[107])^(a[254] & b[108])^(a[253] & b[109])^(a[252] & b[110])^(a[251] & b[111])^(a[250] & b[112])^(a[249] & b[113])^(a[248] & b[114])^(a[247] & b[115])^(a[246] & b[116])^(a[245] & b[117])^(a[244] & b[118])^(a[243] & b[119])^(a[242] & b[120])^(a[241] & b[121])^(a[240] & b[122])^(a[239] & b[123])^(a[238] & b[124])^(a[237] & b[125])^(a[236] & b[126])^(a[235] & b[127])^(a[234] & b[128])^(a[233] & b[129])^(a[232] & b[130])^(a[231] & b[131])^(a[230] & b[132])^(a[229] & b[133])^(a[228] & b[134])^(a[227] & b[135])^(a[226] & b[136])^(a[225] & b[137])^(a[224] & b[138])^(a[223] & b[139])^(a[222] & b[140])^(a[221] & b[141])^(a[220] & b[142])^(a[219] & b[143])^(a[218] & b[144])^(a[217] & b[145])^(a[216] & b[146])^(a[215] & b[147])^(a[214] & b[148])^(a[213] & b[149])^(a[212] & b[150])^(a[211] & b[151])^(a[210] & b[152])^(a[209] & b[153])^(a[208] & b[154])^(a[207] & b[155])^(a[206] & b[156])^(a[205] & b[157])^(a[204] & b[158])^(a[203] & b[159])^(a[202] & b[160])^(a[201] & b[161])^(a[200] & b[162])^(a[199] & b[163])^(a[198] & b[164])^(a[197] & b[165])^(a[196] & b[166])^(a[195] & b[167])^(a[194] & b[168])^(a[193] & b[169])^(a[192] & b[170])^(a[191] & b[171])^(a[190] & b[172])^(a[189] & b[173])^(a[188] & b[174])^(a[187] & b[175])^(a[186] & b[176])^(a[185] & b[177])^(a[184] & b[178])^(a[183] & b[179])^(a[182] & b[180])^(a[181] & b[181])^(a[180] & b[182])^(a[179] & b[183])^(a[178] & b[184])^(a[177] & b[185])^(a[176] & b[186])^(a[175] & b[187])^(a[174] & b[188])^(a[173] & b[189])^(a[172] & b[190])^(a[171] & b[191])^(a[170] & b[192])^(a[169] & b[193])^(a[168] & b[194])^(a[167] & b[195])^(a[166] & b[196])^(a[165] & b[197])^(a[164] & b[198])^(a[163] & b[199])^(a[162] & b[200])^(a[161] & b[201])^(a[160] & b[202])^(a[159] & b[203])^(a[158] & b[204])^(a[157] & b[205])^(a[156] & b[206])^(a[155] & b[207])^(a[154] & b[208])^(a[153] & b[209])^(a[152] & b[210])^(a[151] & b[211])^(a[150] & b[212])^(a[149] & b[213])^(a[148] & b[214])^(a[147] & b[215])^(a[146] & b[216])^(a[145] & b[217])^(a[144] & b[218])^(a[143] & b[219])^(a[142] & b[220])^(a[141] & b[221])^(a[140] & b[222])^(a[139] & b[223])^(a[138] & b[224])^(a[137] & b[225])^(a[136] & b[226])^(a[135] & b[227])^(a[134] & b[228])^(a[133] & b[229])^(a[132] & b[230])^(a[131] & b[231])^(a[130] & b[232])^(a[129] & b[233])^(a[128] & b[234])^(a[127] & b[235])^(a[126] & b[236])^(a[125] & b[237])^(a[124] & b[238])^(a[123] & b[239])^(a[122] & b[240])^(a[121] & b[241])^(a[120] & b[242])^(a[119] & b[243])^(a[118] & b[244])^(a[117] & b[245])^(a[116] & b[246])^(a[115] & b[247])^(a[114] & b[248])^(a[113] & b[249])^(a[112] & b[250])^(a[111] & b[251])^(a[110] & b[252])^(a[109] & b[253])^(a[108] & b[254])^(a[107] & b[255])^(a[106] & b[256])^(a[105] & b[257])^(a[104] & b[258])^(a[103] & b[259])^(a[102] & b[260])^(a[101] & b[261])^(a[100] & b[262])^(a[99] & b[263])^(a[98] & b[264])^(a[97] & b[265])^(a[96] & b[266])^(a[95] & b[267])^(a[94] & b[268])^(a[93] & b[269])^(a[92] & b[270])^(a[91] & b[271])^(a[90] & b[272])^(a[89] & b[273])^(a[88] & b[274])^(a[87] & b[275])^(a[86] & b[276])^(a[85] & b[277])^(a[84] & b[278])^(a[83] & b[279])^(a[82] & b[280])^(a[81] & b[281])^(a[80] & b[282])^(a[79] & b[283])^(a[78] & b[284])^(a[77] & b[285])^(a[76] & b[286])^(a[75] & b[287])^(a[74] & b[288])^(a[73] & b[289])^(a[72] & b[290])^(a[71] & b[291])^(a[70] & b[292])^(a[69] & b[293])^(a[68] & b[294])^(a[67] & b[295])^(a[66] & b[296])^(a[65] & b[297])^(a[64] & b[298])^(a[63] & b[299])^(a[62] & b[300])^(a[61] & b[301])^(a[60] & b[302])^(a[59] & b[303])^(a[58] & b[304])^(a[57] & b[305])^(a[56] & b[306])^(a[55] & b[307])^(a[54] & b[308])^(a[53] & b[309])^(a[52] & b[310])^(a[51] & b[311])^(a[50] & b[312])^(a[49] & b[313])^(a[48] & b[314])^(a[47] & b[315])^(a[46] & b[316])^(a[45] & b[317])^(a[44] & b[318])^(a[43] & b[319])^(a[42] & b[320])^(a[41] & b[321])^(a[40] & b[322])^(a[39] & b[323])^(a[38] & b[324])^(a[37] & b[325])^(a[36] & b[326])^(a[35] & b[327])^(a[34] & b[328])^(a[33] & b[329])^(a[32] & b[330])^(a[31] & b[331])^(a[30] & b[332])^(a[29] & b[333])^(a[28] & b[334])^(a[27] & b[335])^(a[26] & b[336])^(a[25] & b[337])^(a[24] & b[338])^(a[23] & b[339])^(a[22] & b[340])^(a[21] & b[341])^(a[20] & b[342])^(a[19] & b[343])^(a[18] & b[344])^(a[17] & b[345])^(a[16] & b[346])^(a[15] & b[347])^(a[14] & b[348])^(a[13] & b[349])^(a[12] & b[350])^(a[11] & b[351])^(a[10] & b[352])^(a[9] & b[353])^(a[8] & b[354])^(a[7] & b[355])^(a[6] & b[356])^(a[5] & b[357])^(a[4] & b[358])^(a[3] & b[359])^(a[2] & b[360])^(a[1] & b[361])^(a[0] & b[362]);
assign y[363] = (a[363] & b[0])^(a[362] & b[1])^(a[361] & b[2])^(a[360] & b[3])^(a[359] & b[4])^(a[358] & b[5])^(a[357] & b[6])^(a[356] & b[7])^(a[355] & b[8])^(a[354] & b[9])^(a[353] & b[10])^(a[352] & b[11])^(a[351] & b[12])^(a[350] & b[13])^(a[349] & b[14])^(a[348] & b[15])^(a[347] & b[16])^(a[346] & b[17])^(a[345] & b[18])^(a[344] & b[19])^(a[343] & b[20])^(a[342] & b[21])^(a[341] & b[22])^(a[340] & b[23])^(a[339] & b[24])^(a[338] & b[25])^(a[337] & b[26])^(a[336] & b[27])^(a[335] & b[28])^(a[334] & b[29])^(a[333] & b[30])^(a[332] & b[31])^(a[331] & b[32])^(a[330] & b[33])^(a[329] & b[34])^(a[328] & b[35])^(a[327] & b[36])^(a[326] & b[37])^(a[325] & b[38])^(a[324] & b[39])^(a[323] & b[40])^(a[322] & b[41])^(a[321] & b[42])^(a[320] & b[43])^(a[319] & b[44])^(a[318] & b[45])^(a[317] & b[46])^(a[316] & b[47])^(a[315] & b[48])^(a[314] & b[49])^(a[313] & b[50])^(a[312] & b[51])^(a[311] & b[52])^(a[310] & b[53])^(a[309] & b[54])^(a[308] & b[55])^(a[307] & b[56])^(a[306] & b[57])^(a[305] & b[58])^(a[304] & b[59])^(a[303] & b[60])^(a[302] & b[61])^(a[301] & b[62])^(a[300] & b[63])^(a[299] & b[64])^(a[298] & b[65])^(a[297] & b[66])^(a[296] & b[67])^(a[295] & b[68])^(a[294] & b[69])^(a[293] & b[70])^(a[292] & b[71])^(a[291] & b[72])^(a[290] & b[73])^(a[289] & b[74])^(a[288] & b[75])^(a[287] & b[76])^(a[286] & b[77])^(a[285] & b[78])^(a[284] & b[79])^(a[283] & b[80])^(a[282] & b[81])^(a[281] & b[82])^(a[280] & b[83])^(a[279] & b[84])^(a[278] & b[85])^(a[277] & b[86])^(a[276] & b[87])^(a[275] & b[88])^(a[274] & b[89])^(a[273] & b[90])^(a[272] & b[91])^(a[271] & b[92])^(a[270] & b[93])^(a[269] & b[94])^(a[268] & b[95])^(a[267] & b[96])^(a[266] & b[97])^(a[265] & b[98])^(a[264] & b[99])^(a[263] & b[100])^(a[262] & b[101])^(a[261] & b[102])^(a[260] & b[103])^(a[259] & b[104])^(a[258] & b[105])^(a[257] & b[106])^(a[256] & b[107])^(a[255] & b[108])^(a[254] & b[109])^(a[253] & b[110])^(a[252] & b[111])^(a[251] & b[112])^(a[250] & b[113])^(a[249] & b[114])^(a[248] & b[115])^(a[247] & b[116])^(a[246] & b[117])^(a[245] & b[118])^(a[244] & b[119])^(a[243] & b[120])^(a[242] & b[121])^(a[241] & b[122])^(a[240] & b[123])^(a[239] & b[124])^(a[238] & b[125])^(a[237] & b[126])^(a[236] & b[127])^(a[235] & b[128])^(a[234] & b[129])^(a[233] & b[130])^(a[232] & b[131])^(a[231] & b[132])^(a[230] & b[133])^(a[229] & b[134])^(a[228] & b[135])^(a[227] & b[136])^(a[226] & b[137])^(a[225] & b[138])^(a[224] & b[139])^(a[223] & b[140])^(a[222] & b[141])^(a[221] & b[142])^(a[220] & b[143])^(a[219] & b[144])^(a[218] & b[145])^(a[217] & b[146])^(a[216] & b[147])^(a[215] & b[148])^(a[214] & b[149])^(a[213] & b[150])^(a[212] & b[151])^(a[211] & b[152])^(a[210] & b[153])^(a[209] & b[154])^(a[208] & b[155])^(a[207] & b[156])^(a[206] & b[157])^(a[205] & b[158])^(a[204] & b[159])^(a[203] & b[160])^(a[202] & b[161])^(a[201] & b[162])^(a[200] & b[163])^(a[199] & b[164])^(a[198] & b[165])^(a[197] & b[166])^(a[196] & b[167])^(a[195] & b[168])^(a[194] & b[169])^(a[193] & b[170])^(a[192] & b[171])^(a[191] & b[172])^(a[190] & b[173])^(a[189] & b[174])^(a[188] & b[175])^(a[187] & b[176])^(a[186] & b[177])^(a[185] & b[178])^(a[184] & b[179])^(a[183] & b[180])^(a[182] & b[181])^(a[181] & b[182])^(a[180] & b[183])^(a[179] & b[184])^(a[178] & b[185])^(a[177] & b[186])^(a[176] & b[187])^(a[175] & b[188])^(a[174] & b[189])^(a[173] & b[190])^(a[172] & b[191])^(a[171] & b[192])^(a[170] & b[193])^(a[169] & b[194])^(a[168] & b[195])^(a[167] & b[196])^(a[166] & b[197])^(a[165] & b[198])^(a[164] & b[199])^(a[163] & b[200])^(a[162] & b[201])^(a[161] & b[202])^(a[160] & b[203])^(a[159] & b[204])^(a[158] & b[205])^(a[157] & b[206])^(a[156] & b[207])^(a[155] & b[208])^(a[154] & b[209])^(a[153] & b[210])^(a[152] & b[211])^(a[151] & b[212])^(a[150] & b[213])^(a[149] & b[214])^(a[148] & b[215])^(a[147] & b[216])^(a[146] & b[217])^(a[145] & b[218])^(a[144] & b[219])^(a[143] & b[220])^(a[142] & b[221])^(a[141] & b[222])^(a[140] & b[223])^(a[139] & b[224])^(a[138] & b[225])^(a[137] & b[226])^(a[136] & b[227])^(a[135] & b[228])^(a[134] & b[229])^(a[133] & b[230])^(a[132] & b[231])^(a[131] & b[232])^(a[130] & b[233])^(a[129] & b[234])^(a[128] & b[235])^(a[127] & b[236])^(a[126] & b[237])^(a[125] & b[238])^(a[124] & b[239])^(a[123] & b[240])^(a[122] & b[241])^(a[121] & b[242])^(a[120] & b[243])^(a[119] & b[244])^(a[118] & b[245])^(a[117] & b[246])^(a[116] & b[247])^(a[115] & b[248])^(a[114] & b[249])^(a[113] & b[250])^(a[112] & b[251])^(a[111] & b[252])^(a[110] & b[253])^(a[109] & b[254])^(a[108] & b[255])^(a[107] & b[256])^(a[106] & b[257])^(a[105] & b[258])^(a[104] & b[259])^(a[103] & b[260])^(a[102] & b[261])^(a[101] & b[262])^(a[100] & b[263])^(a[99] & b[264])^(a[98] & b[265])^(a[97] & b[266])^(a[96] & b[267])^(a[95] & b[268])^(a[94] & b[269])^(a[93] & b[270])^(a[92] & b[271])^(a[91] & b[272])^(a[90] & b[273])^(a[89] & b[274])^(a[88] & b[275])^(a[87] & b[276])^(a[86] & b[277])^(a[85] & b[278])^(a[84] & b[279])^(a[83] & b[280])^(a[82] & b[281])^(a[81] & b[282])^(a[80] & b[283])^(a[79] & b[284])^(a[78] & b[285])^(a[77] & b[286])^(a[76] & b[287])^(a[75] & b[288])^(a[74] & b[289])^(a[73] & b[290])^(a[72] & b[291])^(a[71] & b[292])^(a[70] & b[293])^(a[69] & b[294])^(a[68] & b[295])^(a[67] & b[296])^(a[66] & b[297])^(a[65] & b[298])^(a[64] & b[299])^(a[63] & b[300])^(a[62] & b[301])^(a[61] & b[302])^(a[60] & b[303])^(a[59] & b[304])^(a[58] & b[305])^(a[57] & b[306])^(a[56] & b[307])^(a[55] & b[308])^(a[54] & b[309])^(a[53] & b[310])^(a[52] & b[311])^(a[51] & b[312])^(a[50] & b[313])^(a[49] & b[314])^(a[48] & b[315])^(a[47] & b[316])^(a[46] & b[317])^(a[45] & b[318])^(a[44] & b[319])^(a[43] & b[320])^(a[42] & b[321])^(a[41] & b[322])^(a[40] & b[323])^(a[39] & b[324])^(a[38] & b[325])^(a[37] & b[326])^(a[36] & b[327])^(a[35] & b[328])^(a[34] & b[329])^(a[33] & b[330])^(a[32] & b[331])^(a[31] & b[332])^(a[30] & b[333])^(a[29] & b[334])^(a[28] & b[335])^(a[27] & b[336])^(a[26] & b[337])^(a[25] & b[338])^(a[24] & b[339])^(a[23] & b[340])^(a[22] & b[341])^(a[21] & b[342])^(a[20] & b[343])^(a[19] & b[344])^(a[18] & b[345])^(a[17] & b[346])^(a[16] & b[347])^(a[15] & b[348])^(a[14] & b[349])^(a[13] & b[350])^(a[12] & b[351])^(a[11] & b[352])^(a[10] & b[353])^(a[9] & b[354])^(a[8] & b[355])^(a[7] & b[356])^(a[6] & b[357])^(a[5] & b[358])^(a[4] & b[359])^(a[3] & b[360])^(a[2] & b[361])^(a[1] & b[362])^(a[0] & b[363]);
assign y[364] = (a[364] & b[0])^(a[363] & b[1])^(a[362] & b[2])^(a[361] & b[3])^(a[360] & b[4])^(a[359] & b[5])^(a[358] & b[6])^(a[357] & b[7])^(a[356] & b[8])^(a[355] & b[9])^(a[354] & b[10])^(a[353] & b[11])^(a[352] & b[12])^(a[351] & b[13])^(a[350] & b[14])^(a[349] & b[15])^(a[348] & b[16])^(a[347] & b[17])^(a[346] & b[18])^(a[345] & b[19])^(a[344] & b[20])^(a[343] & b[21])^(a[342] & b[22])^(a[341] & b[23])^(a[340] & b[24])^(a[339] & b[25])^(a[338] & b[26])^(a[337] & b[27])^(a[336] & b[28])^(a[335] & b[29])^(a[334] & b[30])^(a[333] & b[31])^(a[332] & b[32])^(a[331] & b[33])^(a[330] & b[34])^(a[329] & b[35])^(a[328] & b[36])^(a[327] & b[37])^(a[326] & b[38])^(a[325] & b[39])^(a[324] & b[40])^(a[323] & b[41])^(a[322] & b[42])^(a[321] & b[43])^(a[320] & b[44])^(a[319] & b[45])^(a[318] & b[46])^(a[317] & b[47])^(a[316] & b[48])^(a[315] & b[49])^(a[314] & b[50])^(a[313] & b[51])^(a[312] & b[52])^(a[311] & b[53])^(a[310] & b[54])^(a[309] & b[55])^(a[308] & b[56])^(a[307] & b[57])^(a[306] & b[58])^(a[305] & b[59])^(a[304] & b[60])^(a[303] & b[61])^(a[302] & b[62])^(a[301] & b[63])^(a[300] & b[64])^(a[299] & b[65])^(a[298] & b[66])^(a[297] & b[67])^(a[296] & b[68])^(a[295] & b[69])^(a[294] & b[70])^(a[293] & b[71])^(a[292] & b[72])^(a[291] & b[73])^(a[290] & b[74])^(a[289] & b[75])^(a[288] & b[76])^(a[287] & b[77])^(a[286] & b[78])^(a[285] & b[79])^(a[284] & b[80])^(a[283] & b[81])^(a[282] & b[82])^(a[281] & b[83])^(a[280] & b[84])^(a[279] & b[85])^(a[278] & b[86])^(a[277] & b[87])^(a[276] & b[88])^(a[275] & b[89])^(a[274] & b[90])^(a[273] & b[91])^(a[272] & b[92])^(a[271] & b[93])^(a[270] & b[94])^(a[269] & b[95])^(a[268] & b[96])^(a[267] & b[97])^(a[266] & b[98])^(a[265] & b[99])^(a[264] & b[100])^(a[263] & b[101])^(a[262] & b[102])^(a[261] & b[103])^(a[260] & b[104])^(a[259] & b[105])^(a[258] & b[106])^(a[257] & b[107])^(a[256] & b[108])^(a[255] & b[109])^(a[254] & b[110])^(a[253] & b[111])^(a[252] & b[112])^(a[251] & b[113])^(a[250] & b[114])^(a[249] & b[115])^(a[248] & b[116])^(a[247] & b[117])^(a[246] & b[118])^(a[245] & b[119])^(a[244] & b[120])^(a[243] & b[121])^(a[242] & b[122])^(a[241] & b[123])^(a[240] & b[124])^(a[239] & b[125])^(a[238] & b[126])^(a[237] & b[127])^(a[236] & b[128])^(a[235] & b[129])^(a[234] & b[130])^(a[233] & b[131])^(a[232] & b[132])^(a[231] & b[133])^(a[230] & b[134])^(a[229] & b[135])^(a[228] & b[136])^(a[227] & b[137])^(a[226] & b[138])^(a[225] & b[139])^(a[224] & b[140])^(a[223] & b[141])^(a[222] & b[142])^(a[221] & b[143])^(a[220] & b[144])^(a[219] & b[145])^(a[218] & b[146])^(a[217] & b[147])^(a[216] & b[148])^(a[215] & b[149])^(a[214] & b[150])^(a[213] & b[151])^(a[212] & b[152])^(a[211] & b[153])^(a[210] & b[154])^(a[209] & b[155])^(a[208] & b[156])^(a[207] & b[157])^(a[206] & b[158])^(a[205] & b[159])^(a[204] & b[160])^(a[203] & b[161])^(a[202] & b[162])^(a[201] & b[163])^(a[200] & b[164])^(a[199] & b[165])^(a[198] & b[166])^(a[197] & b[167])^(a[196] & b[168])^(a[195] & b[169])^(a[194] & b[170])^(a[193] & b[171])^(a[192] & b[172])^(a[191] & b[173])^(a[190] & b[174])^(a[189] & b[175])^(a[188] & b[176])^(a[187] & b[177])^(a[186] & b[178])^(a[185] & b[179])^(a[184] & b[180])^(a[183] & b[181])^(a[182] & b[182])^(a[181] & b[183])^(a[180] & b[184])^(a[179] & b[185])^(a[178] & b[186])^(a[177] & b[187])^(a[176] & b[188])^(a[175] & b[189])^(a[174] & b[190])^(a[173] & b[191])^(a[172] & b[192])^(a[171] & b[193])^(a[170] & b[194])^(a[169] & b[195])^(a[168] & b[196])^(a[167] & b[197])^(a[166] & b[198])^(a[165] & b[199])^(a[164] & b[200])^(a[163] & b[201])^(a[162] & b[202])^(a[161] & b[203])^(a[160] & b[204])^(a[159] & b[205])^(a[158] & b[206])^(a[157] & b[207])^(a[156] & b[208])^(a[155] & b[209])^(a[154] & b[210])^(a[153] & b[211])^(a[152] & b[212])^(a[151] & b[213])^(a[150] & b[214])^(a[149] & b[215])^(a[148] & b[216])^(a[147] & b[217])^(a[146] & b[218])^(a[145] & b[219])^(a[144] & b[220])^(a[143] & b[221])^(a[142] & b[222])^(a[141] & b[223])^(a[140] & b[224])^(a[139] & b[225])^(a[138] & b[226])^(a[137] & b[227])^(a[136] & b[228])^(a[135] & b[229])^(a[134] & b[230])^(a[133] & b[231])^(a[132] & b[232])^(a[131] & b[233])^(a[130] & b[234])^(a[129] & b[235])^(a[128] & b[236])^(a[127] & b[237])^(a[126] & b[238])^(a[125] & b[239])^(a[124] & b[240])^(a[123] & b[241])^(a[122] & b[242])^(a[121] & b[243])^(a[120] & b[244])^(a[119] & b[245])^(a[118] & b[246])^(a[117] & b[247])^(a[116] & b[248])^(a[115] & b[249])^(a[114] & b[250])^(a[113] & b[251])^(a[112] & b[252])^(a[111] & b[253])^(a[110] & b[254])^(a[109] & b[255])^(a[108] & b[256])^(a[107] & b[257])^(a[106] & b[258])^(a[105] & b[259])^(a[104] & b[260])^(a[103] & b[261])^(a[102] & b[262])^(a[101] & b[263])^(a[100] & b[264])^(a[99] & b[265])^(a[98] & b[266])^(a[97] & b[267])^(a[96] & b[268])^(a[95] & b[269])^(a[94] & b[270])^(a[93] & b[271])^(a[92] & b[272])^(a[91] & b[273])^(a[90] & b[274])^(a[89] & b[275])^(a[88] & b[276])^(a[87] & b[277])^(a[86] & b[278])^(a[85] & b[279])^(a[84] & b[280])^(a[83] & b[281])^(a[82] & b[282])^(a[81] & b[283])^(a[80] & b[284])^(a[79] & b[285])^(a[78] & b[286])^(a[77] & b[287])^(a[76] & b[288])^(a[75] & b[289])^(a[74] & b[290])^(a[73] & b[291])^(a[72] & b[292])^(a[71] & b[293])^(a[70] & b[294])^(a[69] & b[295])^(a[68] & b[296])^(a[67] & b[297])^(a[66] & b[298])^(a[65] & b[299])^(a[64] & b[300])^(a[63] & b[301])^(a[62] & b[302])^(a[61] & b[303])^(a[60] & b[304])^(a[59] & b[305])^(a[58] & b[306])^(a[57] & b[307])^(a[56] & b[308])^(a[55] & b[309])^(a[54] & b[310])^(a[53] & b[311])^(a[52] & b[312])^(a[51] & b[313])^(a[50] & b[314])^(a[49] & b[315])^(a[48] & b[316])^(a[47] & b[317])^(a[46] & b[318])^(a[45] & b[319])^(a[44] & b[320])^(a[43] & b[321])^(a[42] & b[322])^(a[41] & b[323])^(a[40] & b[324])^(a[39] & b[325])^(a[38] & b[326])^(a[37] & b[327])^(a[36] & b[328])^(a[35] & b[329])^(a[34] & b[330])^(a[33] & b[331])^(a[32] & b[332])^(a[31] & b[333])^(a[30] & b[334])^(a[29] & b[335])^(a[28] & b[336])^(a[27] & b[337])^(a[26] & b[338])^(a[25] & b[339])^(a[24] & b[340])^(a[23] & b[341])^(a[22] & b[342])^(a[21] & b[343])^(a[20] & b[344])^(a[19] & b[345])^(a[18] & b[346])^(a[17] & b[347])^(a[16] & b[348])^(a[15] & b[349])^(a[14] & b[350])^(a[13] & b[351])^(a[12] & b[352])^(a[11] & b[353])^(a[10] & b[354])^(a[9] & b[355])^(a[8] & b[356])^(a[7] & b[357])^(a[6] & b[358])^(a[5] & b[359])^(a[4] & b[360])^(a[3] & b[361])^(a[2] & b[362])^(a[1] & b[363])^(a[0] & b[364]);
assign y[365] = (a[365] & b[0])^(a[364] & b[1])^(a[363] & b[2])^(a[362] & b[3])^(a[361] & b[4])^(a[360] & b[5])^(a[359] & b[6])^(a[358] & b[7])^(a[357] & b[8])^(a[356] & b[9])^(a[355] & b[10])^(a[354] & b[11])^(a[353] & b[12])^(a[352] & b[13])^(a[351] & b[14])^(a[350] & b[15])^(a[349] & b[16])^(a[348] & b[17])^(a[347] & b[18])^(a[346] & b[19])^(a[345] & b[20])^(a[344] & b[21])^(a[343] & b[22])^(a[342] & b[23])^(a[341] & b[24])^(a[340] & b[25])^(a[339] & b[26])^(a[338] & b[27])^(a[337] & b[28])^(a[336] & b[29])^(a[335] & b[30])^(a[334] & b[31])^(a[333] & b[32])^(a[332] & b[33])^(a[331] & b[34])^(a[330] & b[35])^(a[329] & b[36])^(a[328] & b[37])^(a[327] & b[38])^(a[326] & b[39])^(a[325] & b[40])^(a[324] & b[41])^(a[323] & b[42])^(a[322] & b[43])^(a[321] & b[44])^(a[320] & b[45])^(a[319] & b[46])^(a[318] & b[47])^(a[317] & b[48])^(a[316] & b[49])^(a[315] & b[50])^(a[314] & b[51])^(a[313] & b[52])^(a[312] & b[53])^(a[311] & b[54])^(a[310] & b[55])^(a[309] & b[56])^(a[308] & b[57])^(a[307] & b[58])^(a[306] & b[59])^(a[305] & b[60])^(a[304] & b[61])^(a[303] & b[62])^(a[302] & b[63])^(a[301] & b[64])^(a[300] & b[65])^(a[299] & b[66])^(a[298] & b[67])^(a[297] & b[68])^(a[296] & b[69])^(a[295] & b[70])^(a[294] & b[71])^(a[293] & b[72])^(a[292] & b[73])^(a[291] & b[74])^(a[290] & b[75])^(a[289] & b[76])^(a[288] & b[77])^(a[287] & b[78])^(a[286] & b[79])^(a[285] & b[80])^(a[284] & b[81])^(a[283] & b[82])^(a[282] & b[83])^(a[281] & b[84])^(a[280] & b[85])^(a[279] & b[86])^(a[278] & b[87])^(a[277] & b[88])^(a[276] & b[89])^(a[275] & b[90])^(a[274] & b[91])^(a[273] & b[92])^(a[272] & b[93])^(a[271] & b[94])^(a[270] & b[95])^(a[269] & b[96])^(a[268] & b[97])^(a[267] & b[98])^(a[266] & b[99])^(a[265] & b[100])^(a[264] & b[101])^(a[263] & b[102])^(a[262] & b[103])^(a[261] & b[104])^(a[260] & b[105])^(a[259] & b[106])^(a[258] & b[107])^(a[257] & b[108])^(a[256] & b[109])^(a[255] & b[110])^(a[254] & b[111])^(a[253] & b[112])^(a[252] & b[113])^(a[251] & b[114])^(a[250] & b[115])^(a[249] & b[116])^(a[248] & b[117])^(a[247] & b[118])^(a[246] & b[119])^(a[245] & b[120])^(a[244] & b[121])^(a[243] & b[122])^(a[242] & b[123])^(a[241] & b[124])^(a[240] & b[125])^(a[239] & b[126])^(a[238] & b[127])^(a[237] & b[128])^(a[236] & b[129])^(a[235] & b[130])^(a[234] & b[131])^(a[233] & b[132])^(a[232] & b[133])^(a[231] & b[134])^(a[230] & b[135])^(a[229] & b[136])^(a[228] & b[137])^(a[227] & b[138])^(a[226] & b[139])^(a[225] & b[140])^(a[224] & b[141])^(a[223] & b[142])^(a[222] & b[143])^(a[221] & b[144])^(a[220] & b[145])^(a[219] & b[146])^(a[218] & b[147])^(a[217] & b[148])^(a[216] & b[149])^(a[215] & b[150])^(a[214] & b[151])^(a[213] & b[152])^(a[212] & b[153])^(a[211] & b[154])^(a[210] & b[155])^(a[209] & b[156])^(a[208] & b[157])^(a[207] & b[158])^(a[206] & b[159])^(a[205] & b[160])^(a[204] & b[161])^(a[203] & b[162])^(a[202] & b[163])^(a[201] & b[164])^(a[200] & b[165])^(a[199] & b[166])^(a[198] & b[167])^(a[197] & b[168])^(a[196] & b[169])^(a[195] & b[170])^(a[194] & b[171])^(a[193] & b[172])^(a[192] & b[173])^(a[191] & b[174])^(a[190] & b[175])^(a[189] & b[176])^(a[188] & b[177])^(a[187] & b[178])^(a[186] & b[179])^(a[185] & b[180])^(a[184] & b[181])^(a[183] & b[182])^(a[182] & b[183])^(a[181] & b[184])^(a[180] & b[185])^(a[179] & b[186])^(a[178] & b[187])^(a[177] & b[188])^(a[176] & b[189])^(a[175] & b[190])^(a[174] & b[191])^(a[173] & b[192])^(a[172] & b[193])^(a[171] & b[194])^(a[170] & b[195])^(a[169] & b[196])^(a[168] & b[197])^(a[167] & b[198])^(a[166] & b[199])^(a[165] & b[200])^(a[164] & b[201])^(a[163] & b[202])^(a[162] & b[203])^(a[161] & b[204])^(a[160] & b[205])^(a[159] & b[206])^(a[158] & b[207])^(a[157] & b[208])^(a[156] & b[209])^(a[155] & b[210])^(a[154] & b[211])^(a[153] & b[212])^(a[152] & b[213])^(a[151] & b[214])^(a[150] & b[215])^(a[149] & b[216])^(a[148] & b[217])^(a[147] & b[218])^(a[146] & b[219])^(a[145] & b[220])^(a[144] & b[221])^(a[143] & b[222])^(a[142] & b[223])^(a[141] & b[224])^(a[140] & b[225])^(a[139] & b[226])^(a[138] & b[227])^(a[137] & b[228])^(a[136] & b[229])^(a[135] & b[230])^(a[134] & b[231])^(a[133] & b[232])^(a[132] & b[233])^(a[131] & b[234])^(a[130] & b[235])^(a[129] & b[236])^(a[128] & b[237])^(a[127] & b[238])^(a[126] & b[239])^(a[125] & b[240])^(a[124] & b[241])^(a[123] & b[242])^(a[122] & b[243])^(a[121] & b[244])^(a[120] & b[245])^(a[119] & b[246])^(a[118] & b[247])^(a[117] & b[248])^(a[116] & b[249])^(a[115] & b[250])^(a[114] & b[251])^(a[113] & b[252])^(a[112] & b[253])^(a[111] & b[254])^(a[110] & b[255])^(a[109] & b[256])^(a[108] & b[257])^(a[107] & b[258])^(a[106] & b[259])^(a[105] & b[260])^(a[104] & b[261])^(a[103] & b[262])^(a[102] & b[263])^(a[101] & b[264])^(a[100] & b[265])^(a[99] & b[266])^(a[98] & b[267])^(a[97] & b[268])^(a[96] & b[269])^(a[95] & b[270])^(a[94] & b[271])^(a[93] & b[272])^(a[92] & b[273])^(a[91] & b[274])^(a[90] & b[275])^(a[89] & b[276])^(a[88] & b[277])^(a[87] & b[278])^(a[86] & b[279])^(a[85] & b[280])^(a[84] & b[281])^(a[83] & b[282])^(a[82] & b[283])^(a[81] & b[284])^(a[80] & b[285])^(a[79] & b[286])^(a[78] & b[287])^(a[77] & b[288])^(a[76] & b[289])^(a[75] & b[290])^(a[74] & b[291])^(a[73] & b[292])^(a[72] & b[293])^(a[71] & b[294])^(a[70] & b[295])^(a[69] & b[296])^(a[68] & b[297])^(a[67] & b[298])^(a[66] & b[299])^(a[65] & b[300])^(a[64] & b[301])^(a[63] & b[302])^(a[62] & b[303])^(a[61] & b[304])^(a[60] & b[305])^(a[59] & b[306])^(a[58] & b[307])^(a[57] & b[308])^(a[56] & b[309])^(a[55] & b[310])^(a[54] & b[311])^(a[53] & b[312])^(a[52] & b[313])^(a[51] & b[314])^(a[50] & b[315])^(a[49] & b[316])^(a[48] & b[317])^(a[47] & b[318])^(a[46] & b[319])^(a[45] & b[320])^(a[44] & b[321])^(a[43] & b[322])^(a[42] & b[323])^(a[41] & b[324])^(a[40] & b[325])^(a[39] & b[326])^(a[38] & b[327])^(a[37] & b[328])^(a[36] & b[329])^(a[35] & b[330])^(a[34] & b[331])^(a[33] & b[332])^(a[32] & b[333])^(a[31] & b[334])^(a[30] & b[335])^(a[29] & b[336])^(a[28] & b[337])^(a[27] & b[338])^(a[26] & b[339])^(a[25] & b[340])^(a[24] & b[341])^(a[23] & b[342])^(a[22] & b[343])^(a[21] & b[344])^(a[20] & b[345])^(a[19] & b[346])^(a[18] & b[347])^(a[17] & b[348])^(a[16] & b[349])^(a[15] & b[350])^(a[14] & b[351])^(a[13] & b[352])^(a[12] & b[353])^(a[11] & b[354])^(a[10] & b[355])^(a[9] & b[356])^(a[8] & b[357])^(a[7] & b[358])^(a[6] & b[359])^(a[5] & b[360])^(a[4] & b[361])^(a[3] & b[362])^(a[2] & b[363])^(a[1] & b[364])^(a[0] & b[365]);
assign y[366] = (a[366] & b[0])^(a[365] & b[1])^(a[364] & b[2])^(a[363] & b[3])^(a[362] & b[4])^(a[361] & b[5])^(a[360] & b[6])^(a[359] & b[7])^(a[358] & b[8])^(a[357] & b[9])^(a[356] & b[10])^(a[355] & b[11])^(a[354] & b[12])^(a[353] & b[13])^(a[352] & b[14])^(a[351] & b[15])^(a[350] & b[16])^(a[349] & b[17])^(a[348] & b[18])^(a[347] & b[19])^(a[346] & b[20])^(a[345] & b[21])^(a[344] & b[22])^(a[343] & b[23])^(a[342] & b[24])^(a[341] & b[25])^(a[340] & b[26])^(a[339] & b[27])^(a[338] & b[28])^(a[337] & b[29])^(a[336] & b[30])^(a[335] & b[31])^(a[334] & b[32])^(a[333] & b[33])^(a[332] & b[34])^(a[331] & b[35])^(a[330] & b[36])^(a[329] & b[37])^(a[328] & b[38])^(a[327] & b[39])^(a[326] & b[40])^(a[325] & b[41])^(a[324] & b[42])^(a[323] & b[43])^(a[322] & b[44])^(a[321] & b[45])^(a[320] & b[46])^(a[319] & b[47])^(a[318] & b[48])^(a[317] & b[49])^(a[316] & b[50])^(a[315] & b[51])^(a[314] & b[52])^(a[313] & b[53])^(a[312] & b[54])^(a[311] & b[55])^(a[310] & b[56])^(a[309] & b[57])^(a[308] & b[58])^(a[307] & b[59])^(a[306] & b[60])^(a[305] & b[61])^(a[304] & b[62])^(a[303] & b[63])^(a[302] & b[64])^(a[301] & b[65])^(a[300] & b[66])^(a[299] & b[67])^(a[298] & b[68])^(a[297] & b[69])^(a[296] & b[70])^(a[295] & b[71])^(a[294] & b[72])^(a[293] & b[73])^(a[292] & b[74])^(a[291] & b[75])^(a[290] & b[76])^(a[289] & b[77])^(a[288] & b[78])^(a[287] & b[79])^(a[286] & b[80])^(a[285] & b[81])^(a[284] & b[82])^(a[283] & b[83])^(a[282] & b[84])^(a[281] & b[85])^(a[280] & b[86])^(a[279] & b[87])^(a[278] & b[88])^(a[277] & b[89])^(a[276] & b[90])^(a[275] & b[91])^(a[274] & b[92])^(a[273] & b[93])^(a[272] & b[94])^(a[271] & b[95])^(a[270] & b[96])^(a[269] & b[97])^(a[268] & b[98])^(a[267] & b[99])^(a[266] & b[100])^(a[265] & b[101])^(a[264] & b[102])^(a[263] & b[103])^(a[262] & b[104])^(a[261] & b[105])^(a[260] & b[106])^(a[259] & b[107])^(a[258] & b[108])^(a[257] & b[109])^(a[256] & b[110])^(a[255] & b[111])^(a[254] & b[112])^(a[253] & b[113])^(a[252] & b[114])^(a[251] & b[115])^(a[250] & b[116])^(a[249] & b[117])^(a[248] & b[118])^(a[247] & b[119])^(a[246] & b[120])^(a[245] & b[121])^(a[244] & b[122])^(a[243] & b[123])^(a[242] & b[124])^(a[241] & b[125])^(a[240] & b[126])^(a[239] & b[127])^(a[238] & b[128])^(a[237] & b[129])^(a[236] & b[130])^(a[235] & b[131])^(a[234] & b[132])^(a[233] & b[133])^(a[232] & b[134])^(a[231] & b[135])^(a[230] & b[136])^(a[229] & b[137])^(a[228] & b[138])^(a[227] & b[139])^(a[226] & b[140])^(a[225] & b[141])^(a[224] & b[142])^(a[223] & b[143])^(a[222] & b[144])^(a[221] & b[145])^(a[220] & b[146])^(a[219] & b[147])^(a[218] & b[148])^(a[217] & b[149])^(a[216] & b[150])^(a[215] & b[151])^(a[214] & b[152])^(a[213] & b[153])^(a[212] & b[154])^(a[211] & b[155])^(a[210] & b[156])^(a[209] & b[157])^(a[208] & b[158])^(a[207] & b[159])^(a[206] & b[160])^(a[205] & b[161])^(a[204] & b[162])^(a[203] & b[163])^(a[202] & b[164])^(a[201] & b[165])^(a[200] & b[166])^(a[199] & b[167])^(a[198] & b[168])^(a[197] & b[169])^(a[196] & b[170])^(a[195] & b[171])^(a[194] & b[172])^(a[193] & b[173])^(a[192] & b[174])^(a[191] & b[175])^(a[190] & b[176])^(a[189] & b[177])^(a[188] & b[178])^(a[187] & b[179])^(a[186] & b[180])^(a[185] & b[181])^(a[184] & b[182])^(a[183] & b[183])^(a[182] & b[184])^(a[181] & b[185])^(a[180] & b[186])^(a[179] & b[187])^(a[178] & b[188])^(a[177] & b[189])^(a[176] & b[190])^(a[175] & b[191])^(a[174] & b[192])^(a[173] & b[193])^(a[172] & b[194])^(a[171] & b[195])^(a[170] & b[196])^(a[169] & b[197])^(a[168] & b[198])^(a[167] & b[199])^(a[166] & b[200])^(a[165] & b[201])^(a[164] & b[202])^(a[163] & b[203])^(a[162] & b[204])^(a[161] & b[205])^(a[160] & b[206])^(a[159] & b[207])^(a[158] & b[208])^(a[157] & b[209])^(a[156] & b[210])^(a[155] & b[211])^(a[154] & b[212])^(a[153] & b[213])^(a[152] & b[214])^(a[151] & b[215])^(a[150] & b[216])^(a[149] & b[217])^(a[148] & b[218])^(a[147] & b[219])^(a[146] & b[220])^(a[145] & b[221])^(a[144] & b[222])^(a[143] & b[223])^(a[142] & b[224])^(a[141] & b[225])^(a[140] & b[226])^(a[139] & b[227])^(a[138] & b[228])^(a[137] & b[229])^(a[136] & b[230])^(a[135] & b[231])^(a[134] & b[232])^(a[133] & b[233])^(a[132] & b[234])^(a[131] & b[235])^(a[130] & b[236])^(a[129] & b[237])^(a[128] & b[238])^(a[127] & b[239])^(a[126] & b[240])^(a[125] & b[241])^(a[124] & b[242])^(a[123] & b[243])^(a[122] & b[244])^(a[121] & b[245])^(a[120] & b[246])^(a[119] & b[247])^(a[118] & b[248])^(a[117] & b[249])^(a[116] & b[250])^(a[115] & b[251])^(a[114] & b[252])^(a[113] & b[253])^(a[112] & b[254])^(a[111] & b[255])^(a[110] & b[256])^(a[109] & b[257])^(a[108] & b[258])^(a[107] & b[259])^(a[106] & b[260])^(a[105] & b[261])^(a[104] & b[262])^(a[103] & b[263])^(a[102] & b[264])^(a[101] & b[265])^(a[100] & b[266])^(a[99] & b[267])^(a[98] & b[268])^(a[97] & b[269])^(a[96] & b[270])^(a[95] & b[271])^(a[94] & b[272])^(a[93] & b[273])^(a[92] & b[274])^(a[91] & b[275])^(a[90] & b[276])^(a[89] & b[277])^(a[88] & b[278])^(a[87] & b[279])^(a[86] & b[280])^(a[85] & b[281])^(a[84] & b[282])^(a[83] & b[283])^(a[82] & b[284])^(a[81] & b[285])^(a[80] & b[286])^(a[79] & b[287])^(a[78] & b[288])^(a[77] & b[289])^(a[76] & b[290])^(a[75] & b[291])^(a[74] & b[292])^(a[73] & b[293])^(a[72] & b[294])^(a[71] & b[295])^(a[70] & b[296])^(a[69] & b[297])^(a[68] & b[298])^(a[67] & b[299])^(a[66] & b[300])^(a[65] & b[301])^(a[64] & b[302])^(a[63] & b[303])^(a[62] & b[304])^(a[61] & b[305])^(a[60] & b[306])^(a[59] & b[307])^(a[58] & b[308])^(a[57] & b[309])^(a[56] & b[310])^(a[55] & b[311])^(a[54] & b[312])^(a[53] & b[313])^(a[52] & b[314])^(a[51] & b[315])^(a[50] & b[316])^(a[49] & b[317])^(a[48] & b[318])^(a[47] & b[319])^(a[46] & b[320])^(a[45] & b[321])^(a[44] & b[322])^(a[43] & b[323])^(a[42] & b[324])^(a[41] & b[325])^(a[40] & b[326])^(a[39] & b[327])^(a[38] & b[328])^(a[37] & b[329])^(a[36] & b[330])^(a[35] & b[331])^(a[34] & b[332])^(a[33] & b[333])^(a[32] & b[334])^(a[31] & b[335])^(a[30] & b[336])^(a[29] & b[337])^(a[28] & b[338])^(a[27] & b[339])^(a[26] & b[340])^(a[25] & b[341])^(a[24] & b[342])^(a[23] & b[343])^(a[22] & b[344])^(a[21] & b[345])^(a[20] & b[346])^(a[19] & b[347])^(a[18] & b[348])^(a[17] & b[349])^(a[16] & b[350])^(a[15] & b[351])^(a[14] & b[352])^(a[13] & b[353])^(a[12] & b[354])^(a[11] & b[355])^(a[10] & b[356])^(a[9] & b[357])^(a[8] & b[358])^(a[7] & b[359])^(a[6] & b[360])^(a[5] & b[361])^(a[4] & b[362])^(a[3] & b[363])^(a[2] & b[364])^(a[1] & b[365])^(a[0] & b[366]);
assign y[367] = (a[367] & b[0])^(a[366] & b[1])^(a[365] & b[2])^(a[364] & b[3])^(a[363] & b[4])^(a[362] & b[5])^(a[361] & b[6])^(a[360] & b[7])^(a[359] & b[8])^(a[358] & b[9])^(a[357] & b[10])^(a[356] & b[11])^(a[355] & b[12])^(a[354] & b[13])^(a[353] & b[14])^(a[352] & b[15])^(a[351] & b[16])^(a[350] & b[17])^(a[349] & b[18])^(a[348] & b[19])^(a[347] & b[20])^(a[346] & b[21])^(a[345] & b[22])^(a[344] & b[23])^(a[343] & b[24])^(a[342] & b[25])^(a[341] & b[26])^(a[340] & b[27])^(a[339] & b[28])^(a[338] & b[29])^(a[337] & b[30])^(a[336] & b[31])^(a[335] & b[32])^(a[334] & b[33])^(a[333] & b[34])^(a[332] & b[35])^(a[331] & b[36])^(a[330] & b[37])^(a[329] & b[38])^(a[328] & b[39])^(a[327] & b[40])^(a[326] & b[41])^(a[325] & b[42])^(a[324] & b[43])^(a[323] & b[44])^(a[322] & b[45])^(a[321] & b[46])^(a[320] & b[47])^(a[319] & b[48])^(a[318] & b[49])^(a[317] & b[50])^(a[316] & b[51])^(a[315] & b[52])^(a[314] & b[53])^(a[313] & b[54])^(a[312] & b[55])^(a[311] & b[56])^(a[310] & b[57])^(a[309] & b[58])^(a[308] & b[59])^(a[307] & b[60])^(a[306] & b[61])^(a[305] & b[62])^(a[304] & b[63])^(a[303] & b[64])^(a[302] & b[65])^(a[301] & b[66])^(a[300] & b[67])^(a[299] & b[68])^(a[298] & b[69])^(a[297] & b[70])^(a[296] & b[71])^(a[295] & b[72])^(a[294] & b[73])^(a[293] & b[74])^(a[292] & b[75])^(a[291] & b[76])^(a[290] & b[77])^(a[289] & b[78])^(a[288] & b[79])^(a[287] & b[80])^(a[286] & b[81])^(a[285] & b[82])^(a[284] & b[83])^(a[283] & b[84])^(a[282] & b[85])^(a[281] & b[86])^(a[280] & b[87])^(a[279] & b[88])^(a[278] & b[89])^(a[277] & b[90])^(a[276] & b[91])^(a[275] & b[92])^(a[274] & b[93])^(a[273] & b[94])^(a[272] & b[95])^(a[271] & b[96])^(a[270] & b[97])^(a[269] & b[98])^(a[268] & b[99])^(a[267] & b[100])^(a[266] & b[101])^(a[265] & b[102])^(a[264] & b[103])^(a[263] & b[104])^(a[262] & b[105])^(a[261] & b[106])^(a[260] & b[107])^(a[259] & b[108])^(a[258] & b[109])^(a[257] & b[110])^(a[256] & b[111])^(a[255] & b[112])^(a[254] & b[113])^(a[253] & b[114])^(a[252] & b[115])^(a[251] & b[116])^(a[250] & b[117])^(a[249] & b[118])^(a[248] & b[119])^(a[247] & b[120])^(a[246] & b[121])^(a[245] & b[122])^(a[244] & b[123])^(a[243] & b[124])^(a[242] & b[125])^(a[241] & b[126])^(a[240] & b[127])^(a[239] & b[128])^(a[238] & b[129])^(a[237] & b[130])^(a[236] & b[131])^(a[235] & b[132])^(a[234] & b[133])^(a[233] & b[134])^(a[232] & b[135])^(a[231] & b[136])^(a[230] & b[137])^(a[229] & b[138])^(a[228] & b[139])^(a[227] & b[140])^(a[226] & b[141])^(a[225] & b[142])^(a[224] & b[143])^(a[223] & b[144])^(a[222] & b[145])^(a[221] & b[146])^(a[220] & b[147])^(a[219] & b[148])^(a[218] & b[149])^(a[217] & b[150])^(a[216] & b[151])^(a[215] & b[152])^(a[214] & b[153])^(a[213] & b[154])^(a[212] & b[155])^(a[211] & b[156])^(a[210] & b[157])^(a[209] & b[158])^(a[208] & b[159])^(a[207] & b[160])^(a[206] & b[161])^(a[205] & b[162])^(a[204] & b[163])^(a[203] & b[164])^(a[202] & b[165])^(a[201] & b[166])^(a[200] & b[167])^(a[199] & b[168])^(a[198] & b[169])^(a[197] & b[170])^(a[196] & b[171])^(a[195] & b[172])^(a[194] & b[173])^(a[193] & b[174])^(a[192] & b[175])^(a[191] & b[176])^(a[190] & b[177])^(a[189] & b[178])^(a[188] & b[179])^(a[187] & b[180])^(a[186] & b[181])^(a[185] & b[182])^(a[184] & b[183])^(a[183] & b[184])^(a[182] & b[185])^(a[181] & b[186])^(a[180] & b[187])^(a[179] & b[188])^(a[178] & b[189])^(a[177] & b[190])^(a[176] & b[191])^(a[175] & b[192])^(a[174] & b[193])^(a[173] & b[194])^(a[172] & b[195])^(a[171] & b[196])^(a[170] & b[197])^(a[169] & b[198])^(a[168] & b[199])^(a[167] & b[200])^(a[166] & b[201])^(a[165] & b[202])^(a[164] & b[203])^(a[163] & b[204])^(a[162] & b[205])^(a[161] & b[206])^(a[160] & b[207])^(a[159] & b[208])^(a[158] & b[209])^(a[157] & b[210])^(a[156] & b[211])^(a[155] & b[212])^(a[154] & b[213])^(a[153] & b[214])^(a[152] & b[215])^(a[151] & b[216])^(a[150] & b[217])^(a[149] & b[218])^(a[148] & b[219])^(a[147] & b[220])^(a[146] & b[221])^(a[145] & b[222])^(a[144] & b[223])^(a[143] & b[224])^(a[142] & b[225])^(a[141] & b[226])^(a[140] & b[227])^(a[139] & b[228])^(a[138] & b[229])^(a[137] & b[230])^(a[136] & b[231])^(a[135] & b[232])^(a[134] & b[233])^(a[133] & b[234])^(a[132] & b[235])^(a[131] & b[236])^(a[130] & b[237])^(a[129] & b[238])^(a[128] & b[239])^(a[127] & b[240])^(a[126] & b[241])^(a[125] & b[242])^(a[124] & b[243])^(a[123] & b[244])^(a[122] & b[245])^(a[121] & b[246])^(a[120] & b[247])^(a[119] & b[248])^(a[118] & b[249])^(a[117] & b[250])^(a[116] & b[251])^(a[115] & b[252])^(a[114] & b[253])^(a[113] & b[254])^(a[112] & b[255])^(a[111] & b[256])^(a[110] & b[257])^(a[109] & b[258])^(a[108] & b[259])^(a[107] & b[260])^(a[106] & b[261])^(a[105] & b[262])^(a[104] & b[263])^(a[103] & b[264])^(a[102] & b[265])^(a[101] & b[266])^(a[100] & b[267])^(a[99] & b[268])^(a[98] & b[269])^(a[97] & b[270])^(a[96] & b[271])^(a[95] & b[272])^(a[94] & b[273])^(a[93] & b[274])^(a[92] & b[275])^(a[91] & b[276])^(a[90] & b[277])^(a[89] & b[278])^(a[88] & b[279])^(a[87] & b[280])^(a[86] & b[281])^(a[85] & b[282])^(a[84] & b[283])^(a[83] & b[284])^(a[82] & b[285])^(a[81] & b[286])^(a[80] & b[287])^(a[79] & b[288])^(a[78] & b[289])^(a[77] & b[290])^(a[76] & b[291])^(a[75] & b[292])^(a[74] & b[293])^(a[73] & b[294])^(a[72] & b[295])^(a[71] & b[296])^(a[70] & b[297])^(a[69] & b[298])^(a[68] & b[299])^(a[67] & b[300])^(a[66] & b[301])^(a[65] & b[302])^(a[64] & b[303])^(a[63] & b[304])^(a[62] & b[305])^(a[61] & b[306])^(a[60] & b[307])^(a[59] & b[308])^(a[58] & b[309])^(a[57] & b[310])^(a[56] & b[311])^(a[55] & b[312])^(a[54] & b[313])^(a[53] & b[314])^(a[52] & b[315])^(a[51] & b[316])^(a[50] & b[317])^(a[49] & b[318])^(a[48] & b[319])^(a[47] & b[320])^(a[46] & b[321])^(a[45] & b[322])^(a[44] & b[323])^(a[43] & b[324])^(a[42] & b[325])^(a[41] & b[326])^(a[40] & b[327])^(a[39] & b[328])^(a[38] & b[329])^(a[37] & b[330])^(a[36] & b[331])^(a[35] & b[332])^(a[34] & b[333])^(a[33] & b[334])^(a[32] & b[335])^(a[31] & b[336])^(a[30] & b[337])^(a[29] & b[338])^(a[28] & b[339])^(a[27] & b[340])^(a[26] & b[341])^(a[25] & b[342])^(a[24] & b[343])^(a[23] & b[344])^(a[22] & b[345])^(a[21] & b[346])^(a[20] & b[347])^(a[19] & b[348])^(a[18] & b[349])^(a[17] & b[350])^(a[16] & b[351])^(a[15] & b[352])^(a[14] & b[353])^(a[13] & b[354])^(a[12] & b[355])^(a[11] & b[356])^(a[10] & b[357])^(a[9] & b[358])^(a[8] & b[359])^(a[7] & b[360])^(a[6] & b[361])^(a[5] & b[362])^(a[4] & b[363])^(a[3] & b[364])^(a[2] & b[365])^(a[1] & b[366])^(a[0] & b[367]);
assign y[368] = (a[368] & b[0])^(a[367] & b[1])^(a[366] & b[2])^(a[365] & b[3])^(a[364] & b[4])^(a[363] & b[5])^(a[362] & b[6])^(a[361] & b[7])^(a[360] & b[8])^(a[359] & b[9])^(a[358] & b[10])^(a[357] & b[11])^(a[356] & b[12])^(a[355] & b[13])^(a[354] & b[14])^(a[353] & b[15])^(a[352] & b[16])^(a[351] & b[17])^(a[350] & b[18])^(a[349] & b[19])^(a[348] & b[20])^(a[347] & b[21])^(a[346] & b[22])^(a[345] & b[23])^(a[344] & b[24])^(a[343] & b[25])^(a[342] & b[26])^(a[341] & b[27])^(a[340] & b[28])^(a[339] & b[29])^(a[338] & b[30])^(a[337] & b[31])^(a[336] & b[32])^(a[335] & b[33])^(a[334] & b[34])^(a[333] & b[35])^(a[332] & b[36])^(a[331] & b[37])^(a[330] & b[38])^(a[329] & b[39])^(a[328] & b[40])^(a[327] & b[41])^(a[326] & b[42])^(a[325] & b[43])^(a[324] & b[44])^(a[323] & b[45])^(a[322] & b[46])^(a[321] & b[47])^(a[320] & b[48])^(a[319] & b[49])^(a[318] & b[50])^(a[317] & b[51])^(a[316] & b[52])^(a[315] & b[53])^(a[314] & b[54])^(a[313] & b[55])^(a[312] & b[56])^(a[311] & b[57])^(a[310] & b[58])^(a[309] & b[59])^(a[308] & b[60])^(a[307] & b[61])^(a[306] & b[62])^(a[305] & b[63])^(a[304] & b[64])^(a[303] & b[65])^(a[302] & b[66])^(a[301] & b[67])^(a[300] & b[68])^(a[299] & b[69])^(a[298] & b[70])^(a[297] & b[71])^(a[296] & b[72])^(a[295] & b[73])^(a[294] & b[74])^(a[293] & b[75])^(a[292] & b[76])^(a[291] & b[77])^(a[290] & b[78])^(a[289] & b[79])^(a[288] & b[80])^(a[287] & b[81])^(a[286] & b[82])^(a[285] & b[83])^(a[284] & b[84])^(a[283] & b[85])^(a[282] & b[86])^(a[281] & b[87])^(a[280] & b[88])^(a[279] & b[89])^(a[278] & b[90])^(a[277] & b[91])^(a[276] & b[92])^(a[275] & b[93])^(a[274] & b[94])^(a[273] & b[95])^(a[272] & b[96])^(a[271] & b[97])^(a[270] & b[98])^(a[269] & b[99])^(a[268] & b[100])^(a[267] & b[101])^(a[266] & b[102])^(a[265] & b[103])^(a[264] & b[104])^(a[263] & b[105])^(a[262] & b[106])^(a[261] & b[107])^(a[260] & b[108])^(a[259] & b[109])^(a[258] & b[110])^(a[257] & b[111])^(a[256] & b[112])^(a[255] & b[113])^(a[254] & b[114])^(a[253] & b[115])^(a[252] & b[116])^(a[251] & b[117])^(a[250] & b[118])^(a[249] & b[119])^(a[248] & b[120])^(a[247] & b[121])^(a[246] & b[122])^(a[245] & b[123])^(a[244] & b[124])^(a[243] & b[125])^(a[242] & b[126])^(a[241] & b[127])^(a[240] & b[128])^(a[239] & b[129])^(a[238] & b[130])^(a[237] & b[131])^(a[236] & b[132])^(a[235] & b[133])^(a[234] & b[134])^(a[233] & b[135])^(a[232] & b[136])^(a[231] & b[137])^(a[230] & b[138])^(a[229] & b[139])^(a[228] & b[140])^(a[227] & b[141])^(a[226] & b[142])^(a[225] & b[143])^(a[224] & b[144])^(a[223] & b[145])^(a[222] & b[146])^(a[221] & b[147])^(a[220] & b[148])^(a[219] & b[149])^(a[218] & b[150])^(a[217] & b[151])^(a[216] & b[152])^(a[215] & b[153])^(a[214] & b[154])^(a[213] & b[155])^(a[212] & b[156])^(a[211] & b[157])^(a[210] & b[158])^(a[209] & b[159])^(a[208] & b[160])^(a[207] & b[161])^(a[206] & b[162])^(a[205] & b[163])^(a[204] & b[164])^(a[203] & b[165])^(a[202] & b[166])^(a[201] & b[167])^(a[200] & b[168])^(a[199] & b[169])^(a[198] & b[170])^(a[197] & b[171])^(a[196] & b[172])^(a[195] & b[173])^(a[194] & b[174])^(a[193] & b[175])^(a[192] & b[176])^(a[191] & b[177])^(a[190] & b[178])^(a[189] & b[179])^(a[188] & b[180])^(a[187] & b[181])^(a[186] & b[182])^(a[185] & b[183])^(a[184] & b[184])^(a[183] & b[185])^(a[182] & b[186])^(a[181] & b[187])^(a[180] & b[188])^(a[179] & b[189])^(a[178] & b[190])^(a[177] & b[191])^(a[176] & b[192])^(a[175] & b[193])^(a[174] & b[194])^(a[173] & b[195])^(a[172] & b[196])^(a[171] & b[197])^(a[170] & b[198])^(a[169] & b[199])^(a[168] & b[200])^(a[167] & b[201])^(a[166] & b[202])^(a[165] & b[203])^(a[164] & b[204])^(a[163] & b[205])^(a[162] & b[206])^(a[161] & b[207])^(a[160] & b[208])^(a[159] & b[209])^(a[158] & b[210])^(a[157] & b[211])^(a[156] & b[212])^(a[155] & b[213])^(a[154] & b[214])^(a[153] & b[215])^(a[152] & b[216])^(a[151] & b[217])^(a[150] & b[218])^(a[149] & b[219])^(a[148] & b[220])^(a[147] & b[221])^(a[146] & b[222])^(a[145] & b[223])^(a[144] & b[224])^(a[143] & b[225])^(a[142] & b[226])^(a[141] & b[227])^(a[140] & b[228])^(a[139] & b[229])^(a[138] & b[230])^(a[137] & b[231])^(a[136] & b[232])^(a[135] & b[233])^(a[134] & b[234])^(a[133] & b[235])^(a[132] & b[236])^(a[131] & b[237])^(a[130] & b[238])^(a[129] & b[239])^(a[128] & b[240])^(a[127] & b[241])^(a[126] & b[242])^(a[125] & b[243])^(a[124] & b[244])^(a[123] & b[245])^(a[122] & b[246])^(a[121] & b[247])^(a[120] & b[248])^(a[119] & b[249])^(a[118] & b[250])^(a[117] & b[251])^(a[116] & b[252])^(a[115] & b[253])^(a[114] & b[254])^(a[113] & b[255])^(a[112] & b[256])^(a[111] & b[257])^(a[110] & b[258])^(a[109] & b[259])^(a[108] & b[260])^(a[107] & b[261])^(a[106] & b[262])^(a[105] & b[263])^(a[104] & b[264])^(a[103] & b[265])^(a[102] & b[266])^(a[101] & b[267])^(a[100] & b[268])^(a[99] & b[269])^(a[98] & b[270])^(a[97] & b[271])^(a[96] & b[272])^(a[95] & b[273])^(a[94] & b[274])^(a[93] & b[275])^(a[92] & b[276])^(a[91] & b[277])^(a[90] & b[278])^(a[89] & b[279])^(a[88] & b[280])^(a[87] & b[281])^(a[86] & b[282])^(a[85] & b[283])^(a[84] & b[284])^(a[83] & b[285])^(a[82] & b[286])^(a[81] & b[287])^(a[80] & b[288])^(a[79] & b[289])^(a[78] & b[290])^(a[77] & b[291])^(a[76] & b[292])^(a[75] & b[293])^(a[74] & b[294])^(a[73] & b[295])^(a[72] & b[296])^(a[71] & b[297])^(a[70] & b[298])^(a[69] & b[299])^(a[68] & b[300])^(a[67] & b[301])^(a[66] & b[302])^(a[65] & b[303])^(a[64] & b[304])^(a[63] & b[305])^(a[62] & b[306])^(a[61] & b[307])^(a[60] & b[308])^(a[59] & b[309])^(a[58] & b[310])^(a[57] & b[311])^(a[56] & b[312])^(a[55] & b[313])^(a[54] & b[314])^(a[53] & b[315])^(a[52] & b[316])^(a[51] & b[317])^(a[50] & b[318])^(a[49] & b[319])^(a[48] & b[320])^(a[47] & b[321])^(a[46] & b[322])^(a[45] & b[323])^(a[44] & b[324])^(a[43] & b[325])^(a[42] & b[326])^(a[41] & b[327])^(a[40] & b[328])^(a[39] & b[329])^(a[38] & b[330])^(a[37] & b[331])^(a[36] & b[332])^(a[35] & b[333])^(a[34] & b[334])^(a[33] & b[335])^(a[32] & b[336])^(a[31] & b[337])^(a[30] & b[338])^(a[29] & b[339])^(a[28] & b[340])^(a[27] & b[341])^(a[26] & b[342])^(a[25] & b[343])^(a[24] & b[344])^(a[23] & b[345])^(a[22] & b[346])^(a[21] & b[347])^(a[20] & b[348])^(a[19] & b[349])^(a[18] & b[350])^(a[17] & b[351])^(a[16] & b[352])^(a[15] & b[353])^(a[14] & b[354])^(a[13] & b[355])^(a[12] & b[356])^(a[11] & b[357])^(a[10] & b[358])^(a[9] & b[359])^(a[8] & b[360])^(a[7] & b[361])^(a[6] & b[362])^(a[5] & b[363])^(a[4] & b[364])^(a[3] & b[365])^(a[2] & b[366])^(a[1] & b[367])^(a[0] & b[368]);
assign y[369] = (a[369] & b[0])^(a[368] & b[1])^(a[367] & b[2])^(a[366] & b[3])^(a[365] & b[4])^(a[364] & b[5])^(a[363] & b[6])^(a[362] & b[7])^(a[361] & b[8])^(a[360] & b[9])^(a[359] & b[10])^(a[358] & b[11])^(a[357] & b[12])^(a[356] & b[13])^(a[355] & b[14])^(a[354] & b[15])^(a[353] & b[16])^(a[352] & b[17])^(a[351] & b[18])^(a[350] & b[19])^(a[349] & b[20])^(a[348] & b[21])^(a[347] & b[22])^(a[346] & b[23])^(a[345] & b[24])^(a[344] & b[25])^(a[343] & b[26])^(a[342] & b[27])^(a[341] & b[28])^(a[340] & b[29])^(a[339] & b[30])^(a[338] & b[31])^(a[337] & b[32])^(a[336] & b[33])^(a[335] & b[34])^(a[334] & b[35])^(a[333] & b[36])^(a[332] & b[37])^(a[331] & b[38])^(a[330] & b[39])^(a[329] & b[40])^(a[328] & b[41])^(a[327] & b[42])^(a[326] & b[43])^(a[325] & b[44])^(a[324] & b[45])^(a[323] & b[46])^(a[322] & b[47])^(a[321] & b[48])^(a[320] & b[49])^(a[319] & b[50])^(a[318] & b[51])^(a[317] & b[52])^(a[316] & b[53])^(a[315] & b[54])^(a[314] & b[55])^(a[313] & b[56])^(a[312] & b[57])^(a[311] & b[58])^(a[310] & b[59])^(a[309] & b[60])^(a[308] & b[61])^(a[307] & b[62])^(a[306] & b[63])^(a[305] & b[64])^(a[304] & b[65])^(a[303] & b[66])^(a[302] & b[67])^(a[301] & b[68])^(a[300] & b[69])^(a[299] & b[70])^(a[298] & b[71])^(a[297] & b[72])^(a[296] & b[73])^(a[295] & b[74])^(a[294] & b[75])^(a[293] & b[76])^(a[292] & b[77])^(a[291] & b[78])^(a[290] & b[79])^(a[289] & b[80])^(a[288] & b[81])^(a[287] & b[82])^(a[286] & b[83])^(a[285] & b[84])^(a[284] & b[85])^(a[283] & b[86])^(a[282] & b[87])^(a[281] & b[88])^(a[280] & b[89])^(a[279] & b[90])^(a[278] & b[91])^(a[277] & b[92])^(a[276] & b[93])^(a[275] & b[94])^(a[274] & b[95])^(a[273] & b[96])^(a[272] & b[97])^(a[271] & b[98])^(a[270] & b[99])^(a[269] & b[100])^(a[268] & b[101])^(a[267] & b[102])^(a[266] & b[103])^(a[265] & b[104])^(a[264] & b[105])^(a[263] & b[106])^(a[262] & b[107])^(a[261] & b[108])^(a[260] & b[109])^(a[259] & b[110])^(a[258] & b[111])^(a[257] & b[112])^(a[256] & b[113])^(a[255] & b[114])^(a[254] & b[115])^(a[253] & b[116])^(a[252] & b[117])^(a[251] & b[118])^(a[250] & b[119])^(a[249] & b[120])^(a[248] & b[121])^(a[247] & b[122])^(a[246] & b[123])^(a[245] & b[124])^(a[244] & b[125])^(a[243] & b[126])^(a[242] & b[127])^(a[241] & b[128])^(a[240] & b[129])^(a[239] & b[130])^(a[238] & b[131])^(a[237] & b[132])^(a[236] & b[133])^(a[235] & b[134])^(a[234] & b[135])^(a[233] & b[136])^(a[232] & b[137])^(a[231] & b[138])^(a[230] & b[139])^(a[229] & b[140])^(a[228] & b[141])^(a[227] & b[142])^(a[226] & b[143])^(a[225] & b[144])^(a[224] & b[145])^(a[223] & b[146])^(a[222] & b[147])^(a[221] & b[148])^(a[220] & b[149])^(a[219] & b[150])^(a[218] & b[151])^(a[217] & b[152])^(a[216] & b[153])^(a[215] & b[154])^(a[214] & b[155])^(a[213] & b[156])^(a[212] & b[157])^(a[211] & b[158])^(a[210] & b[159])^(a[209] & b[160])^(a[208] & b[161])^(a[207] & b[162])^(a[206] & b[163])^(a[205] & b[164])^(a[204] & b[165])^(a[203] & b[166])^(a[202] & b[167])^(a[201] & b[168])^(a[200] & b[169])^(a[199] & b[170])^(a[198] & b[171])^(a[197] & b[172])^(a[196] & b[173])^(a[195] & b[174])^(a[194] & b[175])^(a[193] & b[176])^(a[192] & b[177])^(a[191] & b[178])^(a[190] & b[179])^(a[189] & b[180])^(a[188] & b[181])^(a[187] & b[182])^(a[186] & b[183])^(a[185] & b[184])^(a[184] & b[185])^(a[183] & b[186])^(a[182] & b[187])^(a[181] & b[188])^(a[180] & b[189])^(a[179] & b[190])^(a[178] & b[191])^(a[177] & b[192])^(a[176] & b[193])^(a[175] & b[194])^(a[174] & b[195])^(a[173] & b[196])^(a[172] & b[197])^(a[171] & b[198])^(a[170] & b[199])^(a[169] & b[200])^(a[168] & b[201])^(a[167] & b[202])^(a[166] & b[203])^(a[165] & b[204])^(a[164] & b[205])^(a[163] & b[206])^(a[162] & b[207])^(a[161] & b[208])^(a[160] & b[209])^(a[159] & b[210])^(a[158] & b[211])^(a[157] & b[212])^(a[156] & b[213])^(a[155] & b[214])^(a[154] & b[215])^(a[153] & b[216])^(a[152] & b[217])^(a[151] & b[218])^(a[150] & b[219])^(a[149] & b[220])^(a[148] & b[221])^(a[147] & b[222])^(a[146] & b[223])^(a[145] & b[224])^(a[144] & b[225])^(a[143] & b[226])^(a[142] & b[227])^(a[141] & b[228])^(a[140] & b[229])^(a[139] & b[230])^(a[138] & b[231])^(a[137] & b[232])^(a[136] & b[233])^(a[135] & b[234])^(a[134] & b[235])^(a[133] & b[236])^(a[132] & b[237])^(a[131] & b[238])^(a[130] & b[239])^(a[129] & b[240])^(a[128] & b[241])^(a[127] & b[242])^(a[126] & b[243])^(a[125] & b[244])^(a[124] & b[245])^(a[123] & b[246])^(a[122] & b[247])^(a[121] & b[248])^(a[120] & b[249])^(a[119] & b[250])^(a[118] & b[251])^(a[117] & b[252])^(a[116] & b[253])^(a[115] & b[254])^(a[114] & b[255])^(a[113] & b[256])^(a[112] & b[257])^(a[111] & b[258])^(a[110] & b[259])^(a[109] & b[260])^(a[108] & b[261])^(a[107] & b[262])^(a[106] & b[263])^(a[105] & b[264])^(a[104] & b[265])^(a[103] & b[266])^(a[102] & b[267])^(a[101] & b[268])^(a[100] & b[269])^(a[99] & b[270])^(a[98] & b[271])^(a[97] & b[272])^(a[96] & b[273])^(a[95] & b[274])^(a[94] & b[275])^(a[93] & b[276])^(a[92] & b[277])^(a[91] & b[278])^(a[90] & b[279])^(a[89] & b[280])^(a[88] & b[281])^(a[87] & b[282])^(a[86] & b[283])^(a[85] & b[284])^(a[84] & b[285])^(a[83] & b[286])^(a[82] & b[287])^(a[81] & b[288])^(a[80] & b[289])^(a[79] & b[290])^(a[78] & b[291])^(a[77] & b[292])^(a[76] & b[293])^(a[75] & b[294])^(a[74] & b[295])^(a[73] & b[296])^(a[72] & b[297])^(a[71] & b[298])^(a[70] & b[299])^(a[69] & b[300])^(a[68] & b[301])^(a[67] & b[302])^(a[66] & b[303])^(a[65] & b[304])^(a[64] & b[305])^(a[63] & b[306])^(a[62] & b[307])^(a[61] & b[308])^(a[60] & b[309])^(a[59] & b[310])^(a[58] & b[311])^(a[57] & b[312])^(a[56] & b[313])^(a[55] & b[314])^(a[54] & b[315])^(a[53] & b[316])^(a[52] & b[317])^(a[51] & b[318])^(a[50] & b[319])^(a[49] & b[320])^(a[48] & b[321])^(a[47] & b[322])^(a[46] & b[323])^(a[45] & b[324])^(a[44] & b[325])^(a[43] & b[326])^(a[42] & b[327])^(a[41] & b[328])^(a[40] & b[329])^(a[39] & b[330])^(a[38] & b[331])^(a[37] & b[332])^(a[36] & b[333])^(a[35] & b[334])^(a[34] & b[335])^(a[33] & b[336])^(a[32] & b[337])^(a[31] & b[338])^(a[30] & b[339])^(a[29] & b[340])^(a[28] & b[341])^(a[27] & b[342])^(a[26] & b[343])^(a[25] & b[344])^(a[24] & b[345])^(a[23] & b[346])^(a[22] & b[347])^(a[21] & b[348])^(a[20] & b[349])^(a[19] & b[350])^(a[18] & b[351])^(a[17] & b[352])^(a[16] & b[353])^(a[15] & b[354])^(a[14] & b[355])^(a[13] & b[356])^(a[12] & b[357])^(a[11] & b[358])^(a[10] & b[359])^(a[9] & b[360])^(a[8] & b[361])^(a[7] & b[362])^(a[6] & b[363])^(a[5] & b[364])^(a[4] & b[365])^(a[3] & b[366])^(a[2] & b[367])^(a[1] & b[368])^(a[0] & b[369]);
assign y[370] = (a[370] & b[0])^(a[369] & b[1])^(a[368] & b[2])^(a[367] & b[3])^(a[366] & b[4])^(a[365] & b[5])^(a[364] & b[6])^(a[363] & b[7])^(a[362] & b[8])^(a[361] & b[9])^(a[360] & b[10])^(a[359] & b[11])^(a[358] & b[12])^(a[357] & b[13])^(a[356] & b[14])^(a[355] & b[15])^(a[354] & b[16])^(a[353] & b[17])^(a[352] & b[18])^(a[351] & b[19])^(a[350] & b[20])^(a[349] & b[21])^(a[348] & b[22])^(a[347] & b[23])^(a[346] & b[24])^(a[345] & b[25])^(a[344] & b[26])^(a[343] & b[27])^(a[342] & b[28])^(a[341] & b[29])^(a[340] & b[30])^(a[339] & b[31])^(a[338] & b[32])^(a[337] & b[33])^(a[336] & b[34])^(a[335] & b[35])^(a[334] & b[36])^(a[333] & b[37])^(a[332] & b[38])^(a[331] & b[39])^(a[330] & b[40])^(a[329] & b[41])^(a[328] & b[42])^(a[327] & b[43])^(a[326] & b[44])^(a[325] & b[45])^(a[324] & b[46])^(a[323] & b[47])^(a[322] & b[48])^(a[321] & b[49])^(a[320] & b[50])^(a[319] & b[51])^(a[318] & b[52])^(a[317] & b[53])^(a[316] & b[54])^(a[315] & b[55])^(a[314] & b[56])^(a[313] & b[57])^(a[312] & b[58])^(a[311] & b[59])^(a[310] & b[60])^(a[309] & b[61])^(a[308] & b[62])^(a[307] & b[63])^(a[306] & b[64])^(a[305] & b[65])^(a[304] & b[66])^(a[303] & b[67])^(a[302] & b[68])^(a[301] & b[69])^(a[300] & b[70])^(a[299] & b[71])^(a[298] & b[72])^(a[297] & b[73])^(a[296] & b[74])^(a[295] & b[75])^(a[294] & b[76])^(a[293] & b[77])^(a[292] & b[78])^(a[291] & b[79])^(a[290] & b[80])^(a[289] & b[81])^(a[288] & b[82])^(a[287] & b[83])^(a[286] & b[84])^(a[285] & b[85])^(a[284] & b[86])^(a[283] & b[87])^(a[282] & b[88])^(a[281] & b[89])^(a[280] & b[90])^(a[279] & b[91])^(a[278] & b[92])^(a[277] & b[93])^(a[276] & b[94])^(a[275] & b[95])^(a[274] & b[96])^(a[273] & b[97])^(a[272] & b[98])^(a[271] & b[99])^(a[270] & b[100])^(a[269] & b[101])^(a[268] & b[102])^(a[267] & b[103])^(a[266] & b[104])^(a[265] & b[105])^(a[264] & b[106])^(a[263] & b[107])^(a[262] & b[108])^(a[261] & b[109])^(a[260] & b[110])^(a[259] & b[111])^(a[258] & b[112])^(a[257] & b[113])^(a[256] & b[114])^(a[255] & b[115])^(a[254] & b[116])^(a[253] & b[117])^(a[252] & b[118])^(a[251] & b[119])^(a[250] & b[120])^(a[249] & b[121])^(a[248] & b[122])^(a[247] & b[123])^(a[246] & b[124])^(a[245] & b[125])^(a[244] & b[126])^(a[243] & b[127])^(a[242] & b[128])^(a[241] & b[129])^(a[240] & b[130])^(a[239] & b[131])^(a[238] & b[132])^(a[237] & b[133])^(a[236] & b[134])^(a[235] & b[135])^(a[234] & b[136])^(a[233] & b[137])^(a[232] & b[138])^(a[231] & b[139])^(a[230] & b[140])^(a[229] & b[141])^(a[228] & b[142])^(a[227] & b[143])^(a[226] & b[144])^(a[225] & b[145])^(a[224] & b[146])^(a[223] & b[147])^(a[222] & b[148])^(a[221] & b[149])^(a[220] & b[150])^(a[219] & b[151])^(a[218] & b[152])^(a[217] & b[153])^(a[216] & b[154])^(a[215] & b[155])^(a[214] & b[156])^(a[213] & b[157])^(a[212] & b[158])^(a[211] & b[159])^(a[210] & b[160])^(a[209] & b[161])^(a[208] & b[162])^(a[207] & b[163])^(a[206] & b[164])^(a[205] & b[165])^(a[204] & b[166])^(a[203] & b[167])^(a[202] & b[168])^(a[201] & b[169])^(a[200] & b[170])^(a[199] & b[171])^(a[198] & b[172])^(a[197] & b[173])^(a[196] & b[174])^(a[195] & b[175])^(a[194] & b[176])^(a[193] & b[177])^(a[192] & b[178])^(a[191] & b[179])^(a[190] & b[180])^(a[189] & b[181])^(a[188] & b[182])^(a[187] & b[183])^(a[186] & b[184])^(a[185] & b[185])^(a[184] & b[186])^(a[183] & b[187])^(a[182] & b[188])^(a[181] & b[189])^(a[180] & b[190])^(a[179] & b[191])^(a[178] & b[192])^(a[177] & b[193])^(a[176] & b[194])^(a[175] & b[195])^(a[174] & b[196])^(a[173] & b[197])^(a[172] & b[198])^(a[171] & b[199])^(a[170] & b[200])^(a[169] & b[201])^(a[168] & b[202])^(a[167] & b[203])^(a[166] & b[204])^(a[165] & b[205])^(a[164] & b[206])^(a[163] & b[207])^(a[162] & b[208])^(a[161] & b[209])^(a[160] & b[210])^(a[159] & b[211])^(a[158] & b[212])^(a[157] & b[213])^(a[156] & b[214])^(a[155] & b[215])^(a[154] & b[216])^(a[153] & b[217])^(a[152] & b[218])^(a[151] & b[219])^(a[150] & b[220])^(a[149] & b[221])^(a[148] & b[222])^(a[147] & b[223])^(a[146] & b[224])^(a[145] & b[225])^(a[144] & b[226])^(a[143] & b[227])^(a[142] & b[228])^(a[141] & b[229])^(a[140] & b[230])^(a[139] & b[231])^(a[138] & b[232])^(a[137] & b[233])^(a[136] & b[234])^(a[135] & b[235])^(a[134] & b[236])^(a[133] & b[237])^(a[132] & b[238])^(a[131] & b[239])^(a[130] & b[240])^(a[129] & b[241])^(a[128] & b[242])^(a[127] & b[243])^(a[126] & b[244])^(a[125] & b[245])^(a[124] & b[246])^(a[123] & b[247])^(a[122] & b[248])^(a[121] & b[249])^(a[120] & b[250])^(a[119] & b[251])^(a[118] & b[252])^(a[117] & b[253])^(a[116] & b[254])^(a[115] & b[255])^(a[114] & b[256])^(a[113] & b[257])^(a[112] & b[258])^(a[111] & b[259])^(a[110] & b[260])^(a[109] & b[261])^(a[108] & b[262])^(a[107] & b[263])^(a[106] & b[264])^(a[105] & b[265])^(a[104] & b[266])^(a[103] & b[267])^(a[102] & b[268])^(a[101] & b[269])^(a[100] & b[270])^(a[99] & b[271])^(a[98] & b[272])^(a[97] & b[273])^(a[96] & b[274])^(a[95] & b[275])^(a[94] & b[276])^(a[93] & b[277])^(a[92] & b[278])^(a[91] & b[279])^(a[90] & b[280])^(a[89] & b[281])^(a[88] & b[282])^(a[87] & b[283])^(a[86] & b[284])^(a[85] & b[285])^(a[84] & b[286])^(a[83] & b[287])^(a[82] & b[288])^(a[81] & b[289])^(a[80] & b[290])^(a[79] & b[291])^(a[78] & b[292])^(a[77] & b[293])^(a[76] & b[294])^(a[75] & b[295])^(a[74] & b[296])^(a[73] & b[297])^(a[72] & b[298])^(a[71] & b[299])^(a[70] & b[300])^(a[69] & b[301])^(a[68] & b[302])^(a[67] & b[303])^(a[66] & b[304])^(a[65] & b[305])^(a[64] & b[306])^(a[63] & b[307])^(a[62] & b[308])^(a[61] & b[309])^(a[60] & b[310])^(a[59] & b[311])^(a[58] & b[312])^(a[57] & b[313])^(a[56] & b[314])^(a[55] & b[315])^(a[54] & b[316])^(a[53] & b[317])^(a[52] & b[318])^(a[51] & b[319])^(a[50] & b[320])^(a[49] & b[321])^(a[48] & b[322])^(a[47] & b[323])^(a[46] & b[324])^(a[45] & b[325])^(a[44] & b[326])^(a[43] & b[327])^(a[42] & b[328])^(a[41] & b[329])^(a[40] & b[330])^(a[39] & b[331])^(a[38] & b[332])^(a[37] & b[333])^(a[36] & b[334])^(a[35] & b[335])^(a[34] & b[336])^(a[33] & b[337])^(a[32] & b[338])^(a[31] & b[339])^(a[30] & b[340])^(a[29] & b[341])^(a[28] & b[342])^(a[27] & b[343])^(a[26] & b[344])^(a[25] & b[345])^(a[24] & b[346])^(a[23] & b[347])^(a[22] & b[348])^(a[21] & b[349])^(a[20] & b[350])^(a[19] & b[351])^(a[18] & b[352])^(a[17] & b[353])^(a[16] & b[354])^(a[15] & b[355])^(a[14] & b[356])^(a[13] & b[357])^(a[12] & b[358])^(a[11] & b[359])^(a[10] & b[360])^(a[9] & b[361])^(a[8] & b[362])^(a[7] & b[363])^(a[6] & b[364])^(a[5] & b[365])^(a[4] & b[366])^(a[3] & b[367])^(a[2] & b[368])^(a[1] & b[369])^(a[0] & b[370]);
assign y[371] = (a[371] & b[0])^(a[370] & b[1])^(a[369] & b[2])^(a[368] & b[3])^(a[367] & b[4])^(a[366] & b[5])^(a[365] & b[6])^(a[364] & b[7])^(a[363] & b[8])^(a[362] & b[9])^(a[361] & b[10])^(a[360] & b[11])^(a[359] & b[12])^(a[358] & b[13])^(a[357] & b[14])^(a[356] & b[15])^(a[355] & b[16])^(a[354] & b[17])^(a[353] & b[18])^(a[352] & b[19])^(a[351] & b[20])^(a[350] & b[21])^(a[349] & b[22])^(a[348] & b[23])^(a[347] & b[24])^(a[346] & b[25])^(a[345] & b[26])^(a[344] & b[27])^(a[343] & b[28])^(a[342] & b[29])^(a[341] & b[30])^(a[340] & b[31])^(a[339] & b[32])^(a[338] & b[33])^(a[337] & b[34])^(a[336] & b[35])^(a[335] & b[36])^(a[334] & b[37])^(a[333] & b[38])^(a[332] & b[39])^(a[331] & b[40])^(a[330] & b[41])^(a[329] & b[42])^(a[328] & b[43])^(a[327] & b[44])^(a[326] & b[45])^(a[325] & b[46])^(a[324] & b[47])^(a[323] & b[48])^(a[322] & b[49])^(a[321] & b[50])^(a[320] & b[51])^(a[319] & b[52])^(a[318] & b[53])^(a[317] & b[54])^(a[316] & b[55])^(a[315] & b[56])^(a[314] & b[57])^(a[313] & b[58])^(a[312] & b[59])^(a[311] & b[60])^(a[310] & b[61])^(a[309] & b[62])^(a[308] & b[63])^(a[307] & b[64])^(a[306] & b[65])^(a[305] & b[66])^(a[304] & b[67])^(a[303] & b[68])^(a[302] & b[69])^(a[301] & b[70])^(a[300] & b[71])^(a[299] & b[72])^(a[298] & b[73])^(a[297] & b[74])^(a[296] & b[75])^(a[295] & b[76])^(a[294] & b[77])^(a[293] & b[78])^(a[292] & b[79])^(a[291] & b[80])^(a[290] & b[81])^(a[289] & b[82])^(a[288] & b[83])^(a[287] & b[84])^(a[286] & b[85])^(a[285] & b[86])^(a[284] & b[87])^(a[283] & b[88])^(a[282] & b[89])^(a[281] & b[90])^(a[280] & b[91])^(a[279] & b[92])^(a[278] & b[93])^(a[277] & b[94])^(a[276] & b[95])^(a[275] & b[96])^(a[274] & b[97])^(a[273] & b[98])^(a[272] & b[99])^(a[271] & b[100])^(a[270] & b[101])^(a[269] & b[102])^(a[268] & b[103])^(a[267] & b[104])^(a[266] & b[105])^(a[265] & b[106])^(a[264] & b[107])^(a[263] & b[108])^(a[262] & b[109])^(a[261] & b[110])^(a[260] & b[111])^(a[259] & b[112])^(a[258] & b[113])^(a[257] & b[114])^(a[256] & b[115])^(a[255] & b[116])^(a[254] & b[117])^(a[253] & b[118])^(a[252] & b[119])^(a[251] & b[120])^(a[250] & b[121])^(a[249] & b[122])^(a[248] & b[123])^(a[247] & b[124])^(a[246] & b[125])^(a[245] & b[126])^(a[244] & b[127])^(a[243] & b[128])^(a[242] & b[129])^(a[241] & b[130])^(a[240] & b[131])^(a[239] & b[132])^(a[238] & b[133])^(a[237] & b[134])^(a[236] & b[135])^(a[235] & b[136])^(a[234] & b[137])^(a[233] & b[138])^(a[232] & b[139])^(a[231] & b[140])^(a[230] & b[141])^(a[229] & b[142])^(a[228] & b[143])^(a[227] & b[144])^(a[226] & b[145])^(a[225] & b[146])^(a[224] & b[147])^(a[223] & b[148])^(a[222] & b[149])^(a[221] & b[150])^(a[220] & b[151])^(a[219] & b[152])^(a[218] & b[153])^(a[217] & b[154])^(a[216] & b[155])^(a[215] & b[156])^(a[214] & b[157])^(a[213] & b[158])^(a[212] & b[159])^(a[211] & b[160])^(a[210] & b[161])^(a[209] & b[162])^(a[208] & b[163])^(a[207] & b[164])^(a[206] & b[165])^(a[205] & b[166])^(a[204] & b[167])^(a[203] & b[168])^(a[202] & b[169])^(a[201] & b[170])^(a[200] & b[171])^(a[199] & b[172])^(a[198] & b[173])^(a[197] & b[174])^(a[196] & b[175])^(a[195] & b[176])^(a[194] & b[177])^(a[193] & b[178])^(a[192] & b[179])^(a[191] & b[180])^(a[190] & b[181])^(a[189] & b[182])^(a[188] & b[183])^(a[187] & b[184])^(a[186] & b[185])^(a[185] & b[186])^(a[184] & b[187])^(a[183] & b[188])^(a[182] & b[189])^(a[181] & b[190])^(a[180] & b[191])^(a[179] & b[192])^(a[178] & b[193])^(a[177] & b[194])^(a[176] & b[195])^(a[175] & b[196])^(a[174] & b[197])^(a[173] & b[198])^(a[172] & b[199])^(a[171] & b[200])^(a[170] & b[201])^(a[169] & b[202])^(a[168] & b[203])^(a[167] & b[204])^(a[166] & b[205])^(a[165] & b[206])^(a[164] & b[207])^(a[163] & b[208])^(a[162] & b[209])^(a[161] & b[210])^(a[160] & b[211])^(a[159] & b[212])^(a[158] & b[213])^(a[157] & b[214])^(a[156] & b[215])^(a[155] & b[216])^(a[154] & b[217])^(a[153] & b[218])^(a[152] & b[219])^(a[151] & b[220])^(a[150] & b[221])^(a[149] & b[222])^(a[148] & b[223])^(a[147] & b[224])^(a[146] & b[225])^(a[145] & b[226])^(a[144] & b[227])^(a[143] & b[228])^(a[142] & b[229])^(a[141] & b[230])^(a[140] & b[231])^(a[139] & b[232])^(a[138] & b[233])^(a[137] & b[234])^(a[136] & b[235])^(a[135] & b[236])^(a[134] & b[237])^(a[133] & b[238])^(a[132] & b[239])^(a[131] & b[240])^(a[130] & b[241])^(a[129] & b[242])^(a[128] & b[243])^(a[127] & b[244])^(a[126] & b[245])^(a[125] & b[246])^(a[124] & b[247])^(a[123] & b[248])^(a[122] & b[249])^(a[121] & b[250])^(a[120] & b[251])^(a[119] & b[252])^(a[118] & b[253])^(a[117] & b[254])^(a[116] & b[255])^(a[115] & b[256])^(a[114] & b[257])^(a[113] & b[258])^(a[112] & b[259])^(a[111] & b[260])^(a[110] & b[261])^(a[109] & b[262])^(a[108] & b[263])^(a[107] & b[264])^(a[106] & b[265])^(a[105] & b[266])^(a[104] & b[267])^(a[103] & b[268])^(a[102] & b[269])^(a[101] & b[270])^(a[100] & b[271])^(a[99] & b[272])^(a[98] & b[273])^(a[97] & b[274])^(a[96] & b[275])^(a[95] & b[276])^(a[94] & b[277])^(a[93] & b[278])^(a[92] & b[279])^(a[91] & b[280])^(a[90] & b[281])^(a[89] & b[282])^(a[88] & b[283])^(a[87] & b[284])^(a[86] & b[285])^(a[85] & b[286])^(a[84] & b[287])^(a[83] & b[288])^(a[82] & b[289])^(a[81] & b[290])^(a[80] & b[291])^(a[79] & b[292])^(a[78] & b[293])^(a[77] & b[294])^(a[76] & b[295])^(a[75] & b[296])^(a[74] & b[297])^(a[73] & b[298])^(a[72] & b[299])^(a[71] & b[300])^(a[70] & b[301])^(a[69] & b[302])^(a[68] & b[303])^(a[67] & b[304])^(a[66] & b[305])^(a[65] & b[306])^(a[64] & b[307])^(a[63] & b[308])^(a[62] & b[309])^(a[61] & b[310])^(a[60] & b[311])^(a[59] & b[312])^(a[58] & b[313])^(a[57] & b[314])^(a[56] & b[315])^(a[55] & b[316])^(a[54] & b[317])^(a[53] & b[318])^(a[52] & b[319])^(a[51] & b[320])^(a[50] & b[321])^(a[49] & b[322])^(a[48] & b[323])^(a[47] & b[324])^(a[46] & b[325])^(a[45] & b[326])^(a[44] & b[327])^(a[43] & b[328])^(a[42] & b[329])^(a[41] & b[330])^(a[40] & b[331])^(a[39] & b[332])^(a[38] & b[333])^(a[37] & b[334])^(a[36] & b[335])^(a[35] & b[336])^(a[34] & b[337])^(a[33] & b[338])^(a[32] & b[339])^(a[31] & b[340])^(a[30] & b[341])^(a[29] & b[342])^(a[28] & b[343])^(a[27] & b[344])^(a[26] & b[345])^(a[25] & b[346])^(a[24] & b[347])^(a[23] & b[348])^(a[22] & b[349])^(a[21] & b[350])^(a[20] & b[351])^(a[19] & b[352])^(a[18] & b[353])^(a[17] & b[354])^(a[16] & b[355])^(a[15] & b[356])^(a[14] & b[357])^(a[13] & b[358])^(a[12] & b[359])^(a[11] & b[360])^(a[10] & b[361])^(a[9] & b[362])^(a[8] & b[363])^(a[7] & b[364])^(a[6] & b[365])^(a[5] & b[366])^(a[4] & b[367])^(a[3] & b[368])^(a[2] & b[369])^(a[1] & b[370])^(a[0] & b[371]);
assign y[372] = (a[372] & b[0])^(a[371] & b[1])^(a[370] & b[2])^(a[369] & b[3])^(a[368] & b[4])^(a[367] & b[5])^(a[366] & b[6])^(a[365] & b[7])^(a[364] & b[8])^(a[363] & b[9])^(a[362] & b[10])^(a[361] & b[11])^(a[360] & b[12])^(a[359] & b[13])^(a[358] & b[14])^(a[357] & b[15])^(a[356] & b[16])^(a[355] & b[17])^(a[354] & b[18])^(a[353] & b[19])^(a[352] & b[20])^(a[351] & b[21])^(a[350] & b[22])^(a[349] & b[23])^(a[348] & b[24])^(a[347] & b[25])^(a[346] & b[26])^(a[345] & b[27])^(a[344] & b[28])^(a[343] & b[29])^(a[342] & b[30])^(a[341] & b[31])^(a[340] & b[32])^(a[339] & b[33])^(a[338] & b[34])^(a[337] & b[35])^(a[336] & b[36])^(a[335] & b[37])^(a[334] & b[38])^(a[333] & b[39])^(a[332] & b[40])^(a[331] & b[41])^(a[330] & b[42])^(a[329] & b[43])^(a[328] & b[44])^(a[327] & b[45])^(a[326] & b[46])^(a[325] & b[47])^(a[324] & b[48])^(a[323] & b[49])^(a[322] & b[50])^(a[321] & b[51])^(a[320] & b[52])^(a[319] & b[53])^(a[318] & b[54])^(a[317] & b[55])^(a[316] & b[56])^(a[315] & b[57])^(a[314] & b[58])^(a[313] & b[59])^(a[312] & b[60])^(a[311] & b[61])^(a[310] & b[62])^(a[309] & b[63])^(a[308] & b[64])^(a[307] & b[65])^(a[306] & b[66])^(a[305] & b[67])^(a[304] & b[68])^(a[303] & b[69])^(a[302] & b[70])^(a[301] & b[71])^(a[300] & b[72])^(a[299] & b[73])^(a[298] & b[74])^(a[297] & b[75])^(a[296] & b[76])^(a[295] & b[77])^(a[294] & b[78])^(a[293] & b[79])^(a[292] & b[80])^(a[291] & b[81])^(a[290] & b[82])^(a[289] & b[83])^(a[288] & b[84])^(a[287] & b[85])^(a[286] & b[86])^(a[285] & b[87])^(a[284] & b[88])^(a[283] & b[89])^(a[282] & b[90])^(a[281] & b[91])^(a[280] & b[92])^(a[279] & b[93])^(a[278] & b[94])^(a[277] & b[95])^(a[276] & b[96])^(a[275] & b[97])^(a[274] & b[98])^(a[273] & b[99])^(a[272] & b[100])^(a[271] & b[101])^(a[270] & b[102])^(a[269] & b[103])^(a[268] & b[104])^(a[267] & b[105])^(a[266] & b[106])^(a[265] & b[107])^(a[264] & b[108])^(a[263] & b[109])^(a[262] & b[110])^(a[261] & b[111])^(a[260] & b[112])^(a[259] & b[113])^(a[258] & b[114])^(a[257] & b[115])^(a[256] & b[116])^(a[255] & b[117])^(a[254] & b[118])^(a[253] & b[119])^(a[252] & b[120])^(a[251] & b[121])^(a[250] & b[122])^(a[249] & b[123])^(a[248] & b[124])^(a[247] & b[125])^(a[246] & b[126])^(a[245] & b[127])^(a[244] & b[128])^(a[243] & b[129])^(a[242] & b[130])^(a[241] & b[131])^(a[240] & b[132])^(a[239] & b[133])^(a[238] & b[134])^(a[237] & b[135])^(a[236] & b[136])^(a[235] & b[137])^(a[234] & b[138])^(a[233] & b[139])^(a[232] & b[140])^(a[231] & b[141])^(a[230] & b[142])^(a[229] & b[143])^(a[228] & b[144])^(a[227] & b[145])^(a[226] & b[146])^(a[225] & b[147])^(a[224] & b[148])^(a[223] & b[149])^(a[222] & b[150])^(a[221] & b[151])^(a[220] & b[152])^(a[219] & b[153])^(a[218] & b[154])^(a[217] & b[155])^(a[216] & b[156])^(a[215] & b[157])^(a[214] & b[158])^(a[213] & b[159])^(a[212] & b[160])^(a[211] & b[161])^(a[210] & b[162])^(a[209] & b[163])^(a[208] & b[164])^(a[207] & b[165])^(a[206] & b[166])^(a[205] & b[167])^(a[204] & b[168])^(a[203] & b[169])^(a[202] & b[170])^(a[201] & b[171])^(a[200] & b[172])^(a[199] & b[173])^(a[198] & b[174])^(a[197] & b[175])^(a[196] & b[176])^(a[195] & b[177])^(a[194] & b[178])^(a[193] & b[179])^(a[192] & b[180])^(a[191] & b[181])^(a[190] & b[182])^(a[189] & b[183])^(a[188] & b[184])^(a[187] & b[185])^(a[186] & b[186])^(a[185] & b[187])^(a[184] & b[188])^(a[183] & b[189])^(a[182] & b[190])^(a[181] & b[191])^(a[180] & b[192])^(a[179] & b[193])^(a[178] & b[194])^(a[177] & b[195])^(a[176] & b[196])^(a[175] & b[197])^(a[174] & b[198])^(a[173] & b[199])^(a[172] & b[200])^(a[171] & b[201])^(a[170] & b[202])^(a[169] & b[203])^(a[168] & b[204])^(a[167] & b[205])^(a[166] & b[206])^(a[165] & b[207])^(a[164] & b[208])^(a[163] & b[209])^(a[162] & b[210])^(a[161] & b[211])^(a[160] & b[212])^(a[159] & b[213])^(a[158] & b[214])^(a[157] & b[215])^(a[156] & b[216])^(a[155] & b[217])^(a[154] & b[218])^(a[153] & b[219])^(a[152] & b[220])^(a[151] & b[221])^(a[150] & b[222])^(a[149] & b[223])^(a[148] & b[224])^(a[147] & b[225])^(a[146] & b[226])^(a[145] & b[227])^(a[144] & b[228])^(a[143] & b[229])^(a[142] & b[230])^(a[141] & b[231])^(a[140] & b[232])^(a[139] & b[233])^(a[138] & b[234])^(a[137] & b[235])^(a[136] & b[236])^(a[135] & b[237])^(a[134] & b[238])^(a[133] & b[239])^(a[132] & b[240])^(a[131] & b[241])^(a[130] & b[242])^(a[129] & b[243])^(a[128] & b[244])^(a[127] & b[245])^(a[126] & b[246])^(a[125] & b[247])^(a[124] & b[248])^(a[123] & b[249])^(a[122] & b[250])^(a[121] & b[251])^(a[120] & b[252])^(a[119] & b[253])^(a[118] & b[254])^(a[117] & b[255])^(a[116] & b[256])^(a[115] & b[257])^(a[114] & b[258])^(a[113] & b[259])^(a[112] & b[260])^(a[111] & b[261])^(a[110] & b[262])^(a[109] & b[263])^(a[108] & b[264])^(a[107] & b[265])^(a[106] & b[266])^(a[105] & b[267])^(a[104] & b[268])^(a[103] & b[269])^(a[102] & b[270])^(a[101] & b[271])^(a[100] & b[272])^(a[99] & b[273])^(a[98] & b[274])^(a[97] & b[275])^(a[96] & b[276])^(a[95] & b[277])^(a[94] & b[278])^(a[93] & b[279])^(a[92] & b[280])^(a[91] & b[281])^(a[90] & b[282])^(a[89] & b[283])^(a[88] & b[284])^(a[87] & b[285])^(a[86] & b[286])^(a[85] & b[287])^(a[84] & b[288])^(a[83] & b[289])^(a[82] & b[290])^(a[81] & b[291])^(a[80] & b[292])^(a[79] & b[293])^(a[78] & b[294])^(a[77] & b[295])^(a[76] & b[296])^(a[75] & b[297])^(a[74] & b[298])^(a[73] & b[299])^(a[72] & b[300])^(a[71] & b[301])^(a[70] & b[302])^(a[69] & b[303])^(a[68] & b[304])^(a[67] & b[305])^(a[66] & b[306])^(a[65] & b[307])^(a[64] & b[308])^(a[63] & b[309])^(a[62] & b[310])^(a[61] & b[311])^(a[60] & b[312])^(a[59] & b[313])^(a[58] & b[314])^(a[57] & b[315])^(a[56] & b[316])^(a[55] & b[317])^(a[54] & b[318])^(a[53] & b[319])^(a[52] & b[320])^(a[51] & b[321])^(a[50] & b[322])^(a[49] & b[323])^(a[48] & b[324])^(a[47] & b[325])^(a[46] & b[326])^(a[45] & b[327])^(a[44] & b[328])^(a[43] & b[329])^(a[42] & b[330])^(a[41] & b[331])^(a[40] & b[332])^(a[39] & b[333])^(a[38] & b[334])^(a[37] & b[335])^(a[36] & b[336])^(a[35] & b[337])^(a[34] & b[338])^(a[33] & b[339])^(a[32] & b[340])^(a[31] & b[341])^(a[30] & b[342])^(a[29] & b[343])^(a[28] & b[344])^(a[27] & b[345])^(a[26] & b[346])^(a[25] & b[347])^(a[24] & b[348])^(a[23] & b[349])^(a[22] & b[350])^(a[21] & b[351])^(a[20] & b[352])^(a[19] & b[353])^(a[18] & b[354])^(a[17] & b[355])^(a[16] & b[356])^(a[15] & b[357])^(a[14] & b[358])^(a[13] & b[359])^(a[12] & b[360])^(a[11] & b[361])^(a[10] & b[362])^(a[9] & b[363])^(a[8] & b[364])^(a[7] & b[365])^(a[6] & b[366])^(a[5] & b[367])^(a[4] & b[368])^(a[3] & b[369])^(a[2] & b[370])^(a[1] & b[371])^(a[0] & b[372]);
assign y[373] = (a[373] & b[0])^(a[372] & b[1])^(a[371] & b[2])^(a[370] & b[3])^(a[369] & b[4])^(a[368] & b[5])^(a[367] & b[6])^(a[366] & b[7])^(a[365] & b[8])^(a[364] & b[9])^(a[363] & b[10])^(a[362] & b[11])^(a[361] & b[12])^(a[360] & b[13])^(a[359] & b[14])^(a[358] & b[15])^(a[357] & b[16])^(a[356] & b[17])^(a[355] & b[18])^(a[354] & b[19])^(a[353] & b[20])^(a[352] & b[21])^(a[351] & b[22])^(a[350] & b[23])^(a[349] & b[24])^(a[348] & b[25])^(a[347] & b[26])^(a[346] & b[27])^(a[345] & b[28])^(a[344] & b[29])^(a[343] & b[30])^(a[342] & b[31])^(a[341] & b[32])^(a[340] & b[33])^(a[339] & b[34])^(a[338] & b[35])^(a[337] & b[36])^(a[336] & b[37])^(a[335] & b[38])^(a[334] & b[39])^(a[333] & b[40])^(a[332] & b[41])^(a[331] & b[42])^(a[330] & b[43])^(a[329] & b[44])^(a[328] & b[45])^(a[327] & b[46])^(a[326] & b[47])^(a[325] & b[48])^(a[324] & b[49])^(a[323] & b[50])^(a[322] & b[51])^(a[321] & b[52])^(a[320] & b[53])^(a[319] & b[54])^(a[318] & b[55])^(a[317] & b[56])^(a[316] & b[57])^(a[315] & b[58])^(a[314] & b[59])^(a[313] & b[60])^(a[312] & b[61])^(a[311] & b[62])^(a[310] & b[63])^(a[309] & b[64])^(a[308] & b[65])^(a[307] & b[66])^(a[306] & b[67])^(a[305] & b[68])^(a[304] & b[69])^(a[303] & b[70])^(a[302] & b[71])^(a[301] & b[72])^(a[300] & b[73])^(a[299] & b[74])^(a[298] & b[75])^(a[297] & b[76])^(a[296] & b[77])^(a[295] & b[78])^(a[294] & b[79])^(a[293] & b[80])^(a[292] & b[81])^(a[291] & b[82])^(a[290] & b[83])^(a[289] & b[84])^(a[288] & b[85])^(a[287] & b[86])^(a[286] & b[87])^(a[285] & b[88])^(a[284] & b[89])^(a[283] & b[90])^(a[282] & b[91])^(a[281] & b[92])^(a[280] & b[93])^(a[279] & b[94])^(a[278] & b[95])^(a[277] & b[96])^(a[276] & b[97])^(a[275] & b[98])^(a[274] & b[99])^(a[273] & b[100])^(a[272] & b[101])^(a[271] & b[102])^(a[270] & b[103])^(a[269] & b[104])^(a[268] & b[105])^(a[267] & b[106])^(a[266] & b[107])^(a[265] & b[108])^(a[264] & b[109])^(a[263] & b[110])^(a[262] & b[111])^(a[261] & b[112])^(a[260] & b[113])^(a[259] & b[114])^(a[258] & b[115])^(a[257] & b[116])^(a[256] & b[117])^(a[255] & b[118])^(a[254] & b[119])^(a[253] & b[120])^(a[252] & b[121])^(a[251] & b[122])^(a[250] & b[123])^(a[249] & b[124])^(a[248] & b[125])^(a[247] & b[126])^(a[246] & b[127])^(a[245] & b[128])^(a[244] & b[129])^(a[243] & b[130])^(a[242] & b[131])^(a[241] & b[132])^(a[240] & b[133])^(a[239] & b[134])^(a[238] & b[135])^(a[237] & b[136])^(a[236] & b[137])^(a[235] & b[138])^(a[234] & b[139])^(a[233] & b[140])^(a[232] & b[141])^(a[231] & b[142])^(a[230] & b[143])^(a[229] & b[144])^(a[228] & b[145])^(a[227] & b[146])^(a[226] & b[147])^(a[225] & b[148])^(a[224] & b[149])^(a[223] & b[150])^(a[222] & b[151])^(a[221] & b[152])^(a[220] & b[153])^(a[219] & b[154])^(a[218] & b[155])^(a[217] & b[156])^(a[216] & b[157])^(a[215] & b[158])^(a[214] & b[159])^(a[213] & b[160])^(a[212] & b[161])^(a[211] & b[162])^(a[210] & b[163])^(a[209] & b[164])^(a[208] & b[165])^(a[207] & b[166])^(a[206] & b[167])^(a[205] & b[168])^(a[204] & b[169])^(a[203] & b[170])^(a[202] & b[171])^(a[201] & b[172])^(a[200] & b[173])^(a[199] & b[174])^(a[198] & b[175])^(a[197] & b[176])^(a[196] & b[177])^(a[195] & b[178])^(a[194] & b[179])^(a[193] & b[180])^(a[192] & b[181])^(a[191] & b[182])^(a[190] & b[183])^(a[189] & b[184])^(a[188] & b[185])^(a[187] & b[186])^(a[186] & b[187])^(a[185] & b[188])^(a[184] & b[189])^(a[183] & b[190])^(a[182] & b[191])^(a[181] & b[192])^(a[180] & b[193])^(a[179] & b[194])^(a[178] & b[195])^(a[177] & b[196])^(a[176] & b[197])^(a[175] & b[198])^(a[174] & b[199])^(a[173] & b[200])^(a[172] & b[201])^(a[171] & b[202])^(a[170] & b[203])^(a[169] & b[204])^(a[168] & b[205])^(a[167] & b[206])^(a[166] & b[207])^(a[165] & b[208])^(a[164] & b[209])^(a[163] & b[210])^(a[162] & b[211])^(a[161] & b[212])^(a[160] & b[213])^(a[159] & b[214])^(a[158] & b[215])^(a[157] & b[216])^(a[156] & b[217])^(a[155] & b[218])^(a[154] & b[219])^(a[153] & b[220])^(a[152] & b[221])^(a[151] & b[222])^(a[150] & b[223])^(a[149] & b[224])^(a[148] & b[225])^(a[147] & b[226])^(a[146] & b[227])^(a[145] & b[228])^(a[144] & b[229])^(a[143] & b[230])^(a[142] & b[231])^(a[141] & b[232])^(a[140] & b[233])^(a[139] & b[234])^(a[138] & b[235])^(a[137] & b[236])^(a[136] & b[237])^(a[135] & b[238])^(a[134] & b[239])^(a[133] & b[240])^(a[132] & b[241])^(a[131] & b[242])^(a[130] & b[243])^(a[129] & b[244])^(a[128] & b[245])^(a[127] & b[246])^(a[126] & b[247])^(a[125] & b[248])^(a[124] & b[249])^(a[123] & b[250])^(a[122] & b[251])^(a[121] & b[252])^(a[120] & b[253])^(a[119] & b[254])^(a[118] & b[255])^(a[117] & b[256])^(a[116] & b[257])^(a[115] & b[258])^(a[114] & b[259])^(a[113] & b[260])^(a[112] & b[261])^(a[111] & b[262])^(a[110] & b[263])^(a[109] & b[264])^(a[108] & b[265])^(a[107] & b[266])^(a[106] & b[267])^(a[105] & b[268])^(a[104] & b[269])^(a[103] & b[270])^(a[102] & b[271])^(a[101] & b[272])^(a[100] & b[273])^(a[99] & b[274])^(a[98] & b[275])^(a[97] & b[276])^(a[96] & b[277])^(a[95] & b[278])^(a[94] & b[279])^(a[93] & b[280])^(a[92] & b[281])^(a[91] & b[282])^(a[90] & b[283])^(a[89] & b[284])^(a[88] & b[285])^(a[87] & b[286])^(a[86] & b[287])^(a[85] & b[288])^(a[84] & b[289])^(a[83] & b[290])^(a[82] & b[291])^(a[81] & b[292])^(a[80] & b[293])^(a[79] & b[294])^(a[78] & b[295])^(a[77] & b[296])^(a[76] & b[297])^(a[75] & b[298])^(a[74] & b[299])^(a[73] & b[300])^(a[72] & b[301])^(a[71] & b[302])^(a[70] & b[303])^(a[69] & b[304])^(a[68] & b[305])^(a[67] & b[306])^(a[66] & b[307])^(a[65] & b[308])^(a[64] & b[309])^(a[63] & b[310])^(a[62] & b[311])^(a[61] & b[312])^(a[60] & b[313])^(a[59] & b[314])^(a[58] & b[315])^(a[57] & b[316])^(a[56] & b[317])^(a[55] & b[318])^(a[54] & b[319])^(a[53] & b[320])^(a[52] & b[321])^(a[51] & b[322])^(a[50] & b[323])^(a[49] & b[324])^(a[48] & b[325])^(a[47] & b[326])^(a[46] & b[327])^(a[45] & b[328])^(a[44] & b[329])^(a[43] & b[330])^(a[42] & b[331])^(a[41] & b[332])^(a[40] & b[333])^(a[39] & b[334])^(a[38] & b[335])^(a[37] & b[336])^(a[36] & b[337])^(a[35] & b[338])^(a[34] & b[339])^(a[33] & b[340])^(a[32] & b[341])^(a[31] & b[342])^(a[30] & b[343])^(a[29] & b[344])^(a[28] & b[345])^(a[27] & b[346])^(a[26] & b[347])^(a[25] & b[348])^(a[24] & b[349])^(a[23] & b[350])^(a[22] & b[351])^(a[21] & b[352])^(a[20] & b[353])^(a[19] & b[354])^(a[18] & b[355])^(a[17] & b[356])^(a[16] & b[357])^(a[15] & b[358])^(a[14] & b[359])^(a[13] & b[360])^(a[12] & b[361])^(a[11] & b[362])^(a[10] & b[363])^(a[9] & b[364])^(a[8] & b[365])^(a[7] & b[366])^(a[6] & b[367])^(a[5] & b[368])^(a[4] & b[369])^(a[3] & b[370])^(a[2] & b[371])^(a[1] & b[372])^(a[0] & b[373]);
assign y[374] = (a[374] & b[0])^(a[373] & b[1])^(a[372] & b[2])^(a[371] & b[3])^(a[370] & b[4])^(a[369] & b[5])^(a[368] & b[6])^(a[367] & b[7])^(a[366] & b[8])^(a[365] & b[9])^(a[364] & b[10])^(a[363] & b[11])^(a[362] & b[12])^(a[361] & b[13])^(a[360] & b[14])^(a[359] & b[15])^(a[358] & b[16])^(a[357] & b[17])^(a[356] & b[18])^(a[355] & b[19])^(a[354] & b[20])^(a[353] & b[21])^(a[352] & b[22])^(a[351] & b[23])^(a[350] & b[24])^(a[349] & b[25])^(a[348] & b[26])^(a[347] & b[27])^(a[346] & b[28])^(a[345] & b[29])^(a[344] & b[30])^(a[343] & b[31])^(a[342] & b[32])^(a[341] & b[33])^(a[340] & b[34])^(a[339] & b[35])^(a[338] & b[36])^(a[337] & b[37])^(a[336] & b[38])^(a[335] & b[39])^(a[334] & b[40])^(a[333] & b[41])^(a[332] & b[42])^(a[331] & b[43])^(a[330] & b[44])^(a[329] & b[45])^(a[328] & b[46])^(a[327] & b[47])^(a[326] & b[48])^(a[325] & b[49])^(a[324] & b[50])^(a[323] & b[51])^(a[322] & b[52])^(a[321] & b[53])^(a[320] & b[54])^(a[319] & b[55])^(a[318] & b[56])^(a[317] & b[57])^(a[316] & b[58])^(a[315] & b[59])^(a[314] & b[60])^(a[313] & b[61])^(a[312] & b[62])^(a[311] & b[63])^(a[310] & b[64])^(a[309] & b[65])^(a[308] & b[66])^(a[307] & b[67])^(a[306] & b[68])^(a[305] & b[69])^(a[304] & b[70])^(a[303] & b[71])^(a[302] & b[72])^(a[301] & b[73])^(a[300] & b[74])^(a[299] & b[75])^(a[298] & b[76])^(a[297] & b[77])^(a[296] & b[78])^(a[295] & b[79])^(a[294] & b[80])^(a[293] & b[81])^(a[292] & b[82])^(a[291] & b[83])^(a[290] & b[84])^(a[289] & b[85])^(a[288] & b[86])^(a[287] & b[87])^(a[286] & b[88])^(a[285] & b[89])^(a[284] & b[90])^(a[283] & b[91])^(a[282] & b[92])^(a[281] & b[93])^(a[280] & b[94])^(a[279] & b[95])^(a[278] & b[96])^(a[277] & b[97])^(a[276] & b[98])^(a[275] & b[99])^(a[274] & b[100])^(a[273] & b[101])^(a[272] & b[102])^(a[271] & b[103])^(a[270] & b[104])^(a[269] & b[105])^(a[268] & b[106])^(a[267] & b[107])^(a[266] & b[108])^(a[265] & b[109])^(a[264] & b[110])^(a[263] & b[111])^(a[262] & b[112])^(a[261] & b[113])^(a[260] & b[114])^(a[259] & b[115])^(a[258] & b[116])^(a[257] & b[117])^(a[256] & b[118])^(a[255] & b[119])^(a[254] & b[120])^(a[253] & b[121])^(a[252] & b[122])^(a[251] & b[123])^(a[250] & b[124])^(a[249] & b[125])^(a[248] & b[126])^(a[247] & b[127])^(a[246] & b[128])^(a[245] & b[129])^(a[244] & b[130])^(a[243] & b[131])^(a[242] & b[132])^(a[241] & b[133])^(a[240] & b[134])^(a[239] & b[135])^(a[238] & b[136])^(a[237] & b[137])^(a[236] & b[138])^(a[235] & b[139])^(a[234] & b[140])^(a[233] & b[141])^(a[232] & b[142])^(a[231] & b[143])^(a[230] & b[144])^(a[229] & b[145])^(a[228] & b[146])^(a[227] & b[147])^(a[226] & b[148])^(a[225] & b[149])^(a[224] & b[150])^(a[223] & b[151])^(a[222] & b[152])^(a[221] & b[153])^(a[220] & b[154])^(a[219] & b[155])^(a[218] & b[156])^(a[217] & b[157])^(a[216] & b[158])^(a[215] & b[159])^(a[214] & b[160])^(a[213] & b[161])^(a[212] & b[162])^(a[211] & b[163])^(a[210] & b[164])^(a[209] & b[165])^(a[208] & b[166])^(a[207] & b[167])^(a[206] & b[168])^(a[205] & b[169])^(a[204] & b[170])^(a[203] & b[171])^(a[202] & b[172])^(a[201] & b[173])^(a[200] & b[174])^(a[199] & b[175])^(a[198] & b[176])^(a[197] & b[177])^(a[196] & b[178])^(a[195] & b[179])^(a[194] & b[180])^(a[193] & b[181])^(a[192] & b[182])^(a[191] & b[183])^(a[190] & b[184])^(a[189] & b[185])^(a[188] & b[186])^(a[187] & b[187])^(a[186] & b[188])^(a[185] & b[189])^(a[184] & b[190])^(a[183] & b[191])^(a[182] & b[192])^(a[181] & b[193])^(a[180] & b[194])^(a[179] & b[195])^(a[178] & b[196])^(a[177] & b[197])^(a[176] & b[198])^(a[175] & b[199])^(a[174] & b[200])^(a[173] & b[201])^(a[172] & b[202])^(a[171] & b[203])^(a[170] & b[204])^(a[169] & b[205])^(a[168] & b[206])^(a[167] & b[207])^(a[166] & b[208])^(a[165] & b[209])^(a[164] & b[210])^(a[163] & b[211])^(a[162] & b[212])^(a[161] & b[213])^(a[160] & b[214])^(a[159] & b[215])^(a[158] & b[216])^(a[157] & b[217])^(a[156] & b[218])^(a[155] & b[219])^(a[154] & b[220])^(a[153] & b[221])^(a[152] & b[222])^(a[151] & b[223])^(a[150] & b[224])^(a[149] & b[225])^(a[148] & b[226])^(a[147] & b[227])^(a[146] & b[228])^(a[145] & b[229])^(a[144] & b[230])^(a[143] & b[231])^(a[142] & b[232])^(a[141] & b[233])^(a[140] & b[234])^(a[139] & b[235])^(a[138] & b[236])^(a[137] & b[237])^(a[136] & b[238])^(a[135] & b[239])^(a[134] & b[240])^(a[133] & b[241])^(a[132] & b[242])^(a[131] & b[243])^(a[130] & b[244])^(a[129] & b[245])^(a[128] & b[246])^(a[127] & b[247])^(a[126] & b[248])^(a[125] & b[249])^(a[124] & b[250])^(a[123] & b[251])^(a[122] & b[252])^(a[121] & b[253])^(a[120] & b[254])^(a[119] & b[255])^(a[118] & b[256])^(a[117] & b[257])^(a[116] & b[258])^(a[115] & b[259])^(a[114] & b[260])^(a[113] & b[261])^(a[112] & b[262])^(a[111] & b[263])^(a[110] & b[264])^(a[109] & b[265])^(a[108] & b[266])^(a[107] & b[267])^(a[106] & b[268])^(a[105] & b[269])^(a[104] & b[270])^(a[103] & b[271])^(a[102] & b[272])^(a[101] & b[273])^(a[100] & b[274])^(a[99] & b[275])^(a[98] & b[276])^(a[97] & b[277])^(a[96] & b[278])^(a[95] & b[279])^(a[94] & b[280])^(a[93] & b[281])^(a[92] & b[282])^(a[91] & b[283])^(a[90] & b[284])^(a[89] & b[285])^(a[88] & b[286])^(a[87] & b[287])^(a[86] & b[288])^(a[85] & b[289])^(a[84] & b[290])^(a[83] & b[291])^(a[82] & b[292])^(a[81] & b[293])^(a[80] & b[294])^(a[79] & b[295])^(a[78] & b[296])^(a[77] & b[297])^(a[76] & b[298])^(a[75] & b[299])^(a[74] & b[300])^(a[73] & b[301])^(a[72] & b[302])^(a[71] & b[303])^(a[70] & b[304])^(a[69] & b[305])^(a[68] & b[306])^(a[67] & b[307])^(a[66] & b[308])^(a[65] & b[309])^(a[64] & b[310])^(a[63] & b[311])^(a[62] & b[312])^(a[61] & b[313])^(a[60] & b[314])^(a[59] & b[315])^(a[58] & b[316])^(a[57] & b[317])^(a[56] & b[318])^(a[55] & b[319])^(a[54] & b[320])^(a[53] & b[321])^(a[52] & b[322])^(a[51] & b[323])^(a[50] & b[324])^(a[49] & b[325])^(a[48] & b[326])^(a[47] & b[327])^(a[46] & b[328])^(a[45] & b[329])^(a[44] & b[330])^(a[43] & b[331])^(a[42] & b[332])^(a[41] & b[333])^(a[40] & b[334])^(a[39] & b[335])^(a[38] & b[336])^(a[37] & b[337])^(a[36] & b[338])^(a[35] & b[339])^(a[34] & b[340])^(a[33] & b[341])^(a[32] & b[342])^(a[31] & b[343])^(a[30] & b[344])^(a[29] & b[345])^(a[28] & b[346])^(a[27] & b[347])^(a[26] & b[348])^(a[25] & b[349])^(a[24] & b[350])^(a[23] & b[351])^(a[22] & b[352])^(a[21] & b[353])^(a[20] & b[354])^(a[19] & b[355])^(a[18] & b[356])^(a[17] & b[357])^(a[16] & b[358])^(a[15] & b[359])^(a[14] & b[360])^(a[13] & b[361])^(a[12] & b[362])^(a[11] & b[363])^(a[10] & b[364])^(a[9] & b[365])^(a[8] & b[366])^(a[7] & b[367])^(a[6] & b[368])^(a[5] & b[369])^(a[4] & b[370])^(a[3] & b[371])^(a[2] & b[372])^(a[1] & b[373])^(a[0] & b[374]);
assign y[375] = (a[375] & b[0])^(a[374] & b[1])^(a[373] & b[2])^(a[372] & b[3])^(a[371] & b[4])^(a[370] & b[5])^(a[369] & b[6])^(a[368] & b[7])^(a[367] & b[8])^(a[366] & b[9])^(a[365] & b[10])^(a[364] & b[11])^(a[363] & b[12])^(a[362] & b[13])^(a[361] & b[14])^(a[360] & b[15])^(a[359] & b[16])^(a[358] & b[17])^(a[357] & b[18])^(a[356] & b[19])^(a[355] & b[20])^(a[354] & b[21])^(a[353] & b[22])^(a[352] & b[23])^(a[351] & b[24])^(a[350] & b[25])^(a[349] & b[26])^(a[348] & b[27])^(a[347] & b[28])^(a[346] & b[29])^(a[345] & b[30])^(a[344] & b[31])^(a[343] & b[32])^(a[342] & b[33])^(a[341] & b[34])^(a[340] & b[35])^(a[339] & b[36])^(a[338] & b[37])^(a[337] & b[38])^(a[336] & b[39])^(a[335] & b[40])^(a[334] & b[41])^(a[333] & b[42])^(a[332] & b[43])^(a[331] & b[44])^(a[330] & b[45])^(a[329] & b[46])^(a[328] & b[47])^(a[327] & b[48])^(a[326] & b[49])^(a[325] & b[50])^(a[324] & b[51])^(a[323] & b[52])^(a[322] & b[53])^(a[321] & b[54])^(a[320] & b[55])^(a[319] & b[56])^(a[318] & b[57])^(a[317] & b[58])^(a[316] & b[59])^(a[315] & b[60])^(a[314] & b[61])^(a[313] & b[62])^(a[312] & b[63])^(a[311] & b[64])^(a[310] & b[65])^(a[309] & b[66])^(a[308] & b[67])^(a[307] & b[68])^(a[306] & b[69])^(a[305] & b[70])^(a[304] & b[71])^(a[303] & b[72])^(a[302] & b[73])^(a[301] & b[74])^(a[300] & b[75])^(a[299] & b[76])^(a[298] & b[77])^(a[297] & b[78])^(a[296] & b[79])^(a[295] & b[80])^(a[294] & b[81])^(a[293] & b[82])^(a[292] & b[83])^(a[291] & b[84])^(a[290] & b[85])^(a[289] & b[86])^(a[288] & b[87])^(a[287] & b[88])^(a[286] & b[89])^(a[285] & b[90])^(a[284] & b[91])^(a[283] & b[92])^(a[282] & b[93])^(a[281] & b[94])^(a[280] & b[95])^(a[279] & b[96])^(a[278] & b[97])^(a[277] & b[98])^(a[276] & b[99])^(a[275] & b[100])^(a[274] & b[101])^(a[273] & b[102])^(a[272] & b[103])^(a[271] & b[104])^(a[270] & b[105])^(a[269] & b[106])^(a[268] & b[107])^(a[267] & b[108])^(a[266] & b[109])^(a[265] & b[110])^(a[264] & b[111])^(a[263] & b[112])^(a[262] & b[113])^(a[261] & b[114])^(a[260] & b[115])^(a[259] & b[116])^(a[258] & b[117])^(a[257] & b[118])^(a[256] & b[119])^(a[255] & b[120])^(a[254] & b[121])^(a[253] & b[122])^(a[252] & b[123])^(a[251] & b[124])^(a[250] & b[125])^(a[249] & b[126])^(a[248] & b[127])^(a[247] & b[128])^(a[246] & b[129])^(a[245] & b[130])^(a[244] & b[131])^(a[243] & b[132])^(a[242] & b[133])^(a[241] & b[134])^(a[240] & b[135])^(a[239] & b[136])^(a[238] & b[137])^(a[237] & b[138])^(a[236] & b[139])^(a[235] & b[140])^(a[234] & b[141])^(a[233] & b[142])^(a[232] & b[143])^(a[231] & b[144])^(a[230] & b[145])^(a[229] & b[146])^(a[228] & b[147])^(a[227] & b[148])^(a[226] & b[149])^(a[225] & b[150])^(a[224] & b[151])^(a[223] & b[152])^(a[222] & b[153])^(a[221] & b[154])^(a[220] & b[155])^(a[219] & b[156])^(a[218] & b[157])^(a[217] & b[158])^(a[216] & b[159])^(a[215] & b[160])^(a[214] & b[161])^(a[213] & b[162])^(a[212] & b[163])^(a[211] & b[164])^(a[210] & b[165])^(a[209] & b[166])^(a[208] & b[167])^(a[207] & b[168])^(a[206] & b[169])^(a[205] & b[170])^(a[204] & b[171])^(a[203] & b[172])^(a[202] & b[173])^(a[201] & b[174])^(a[200] & b[175])^(a[199] & b[176])^(a[198] & b[177])^(a[197] & b[178])^(a[196] & b[179])^(a[195] & b[180])^(a[194] & b[181])^(a[193] & b[182])^(a[192] & b[183])^(a[191] & b[184])^(a[190] & b[185])^(a[189] & b[186])^(a[188] & b[187])^(a[187] & b[188])^(a[186] & b[189])^(a[185] & b[190])^(a[184] & b[191])^(a[183] & b[192])^(a[182] & b[193])^(a[181] & b[194])^(a[180] & b[195])^(a[179] & b[196])^(a[178] & b[197])^(a[177] & b[198])^(a[176] & b[199])^(a[175] & b[200])^(a[174] & b[201])^(a[173] & b[202])^(a[172] & b[203])^(a[171] & b[204])^(a[170] & b[205])^(a[169] & b[206])^(a[168] & b[207])^(a[167] & b[208])^(a[166] & b[209])^(a[165] & b[210])^(a[164] & b[211])^(a[163] & b[212])^(a[162] & b[213])^(a[161] & b[214])^(a[160] & b[215])^(a[159] & b[216])^(a[158] & b[217])^(a[157] & b[218])^(a[156] & b[219])^(a[155] & b[220])^(a[154] & b[221])^(a[153] & b[222])^(a[152] & b[223])^(a[151] & b[224])^(a[150] & b[225])^(a[149] & b[226])^(a[148] & b[227])^(a[147] & b[228])^(a[146] & b[229])^(a[145] & b[230])^(a[144] & b[231])^(a[143] & b[232])^(a[142] & b[233])^(a[141] & b[234])^(a[140] & b[235])^(a[139] & b[236])^(a[138] & b[237])^(a[137] & b[238])^(a[136] & b[239])^(a[135] & b[240])^(a[134] & b[241])^(a[133] & b[242])^(a[132] & b[243])^(a[131] & b[244])^(a[130] & b[245])^(a[129] & b[246])^(a[128] & b[247])^(a[127] & b[248])^(a[126] & b[249])^(a[125] & b[250])^(a[124] & b[251])^(a[123] & b[252])^(a[122] & b[253])^(a[121] & b[254])^(a[120] & b[255])^(a[119] & b[256])^(a[118] & b[257])^(a[117] & b[258])^(a[116] & b[259])^(a[115] & b[260])^(a[114] & b[261])^(a[113] & b[262])^(a[112] & b[263])^(a[111] & b[264])^(a[110] & b[265])^(a[109] & b[266])^(a[108] & b[267])^(a[107] & b[268])^(a[106] & b[269])^(a[105] & b[270])^(a[104] & b[271])^(a[103] & b[272])^(a[102] & b[273])^(a[101] & b[274])^(a[100] & b[275])^(a[99] & b[276])^(a[98] & b[277])^(a[97] & b[278])^(a[96] & b[279])^(a[95] & b[280])^(a[94] & b[281])^(a[93] & b[282])^(a[92] & b[283])^(a[91] & b[284])^(a[90] & b[285])^(a[89] & b[286])^(a[88] & b[287])^(a[87] & b[288])^(a[86] & b[289])^(a[85] & b[290])^(a[84] & b[291])^(a[83] & b[292])^(a[82] & b[293])^(a[81] & b[294])^(a[80] & b[295])^(a[79] & b[296])^(a[78] & b[297])^(a[77] & b[298])^(a[76] & b[299])^(a[75] & b[300])^(a[74] & b[301])^(a[73] & b[302])^(a[72] & b[303])^(a[71] & b[304])^(a[70] & b[305])^(a[69] & b[306])^(a[68] & b[307])^(a[67] & b[308])^(a[66] & b[309])^(a[65] & b[310])^(a[64] & b[311])^(a[63] & b[312])^(a[62] & b[313])^(a[61] & b[314])^(a[60] & b[315])^(a[59] & b[316])^(a[58] & b[317])^(a[57] & b[318])^(a[56] & b[319])^(a[55] & b[320])^(a[54] & b[321])^(a[53] & b[322])^(a[52] & b[323])^(a[51] & b[324])^(a[50] & b[325])^(a[49] & b[326])^(a[48] & b[327])^(a[47] & b[328])^(a[46] & b[329])^(a[45] & b[330])^(a[44] & b[331])^(a[43] & b[332])^(a[42] & b[333])^(a[41] & b[334])^(a[40] & b[335])^(a[39] & b[336])^(a[38] & b[337])^(a[37] & b[338])^(a[36] & b[339])^(a[35] & b[340])^(a[34] & b[341])^(a[33] & b[342])^(a[32] & b[343])^(a[31] & b[344])^(a[30] & b[345])^(a[29] & b[346])^(a[28] & b[347])^(a[27] & b[348])^(a[26] & b[349])^(a[25] & b[350])^(a[24] & b[351])^(a[23] & b[352])^(a[22] & b[353])^(a[21] & b[354])^(a[20] & b[355])^(a[19] & b[356])^(a[18] & b[357])^(a[17] & b[358])^(a[16] & b[359])^(a[15] & b[360])^(a[14] & b[361])^(a[13] & b[362])^(a[12] & b[363])^(a[11] & b[364])^(a[10] & b[365])^(a[9] & b[366])^(a[8] & b[367])^(a[7] & b[368])^(a[6] & b[369])^(a[5] & b[370])^(a[4] & b[371])^(a[3] & b[372])^(a[2] & b[373])^(a[1] & b[374])^(a[0] & b[375]);
assign y[376] = (a[376] & b[0])^(a[375] & b[1])^(a[374] & b[2])^(a[373] & b[3])^(a[372] & b[4])^(a[371] & b[5])^(a[370] & b[6])^(a[369] & b[7])^(a[368] & b[8])^(a[367] & b[9])^(a[366] & b[10])^(a[365] & b[11])^(a[364] & b[12])^(a[363] & b[13])^(a[362] & b[14])^(a[361] & b[15])^(a[360] & b[16])^(a[359] & b[17])^(a[358] & b[18])^(a[357] & b[19])^(a[356] & b[20])^(a[355] & b[21])^(a[354] & b[22])^(a[353] & b[23])^(a[352] & b[24])^(a[351] & b[25])^(a[350] & b[26])^(a[349] & b[27])^(a[348] & b[28])^(a[347] & b[29])^(a[346] & b[30])^(a[345] & b[31])^(a[344] & b[32])^(a[343] & b[33])^(a[342] & b[34])^(a[341] & b[35])^(a[340] & b[36])^(a[339] & b[37])^(a[338] & b[38])^(a[337] & b[39])^(a[336] & b[40])^(a[335] & b[41])^(a[334] & b[42])^(a[333] & b[43])^(a[332] & b[44])^(a[331] & b[45])^(a[330] & b[46])^(a[329] & b[47])^(a[328] & b[48])^(a[327] & b[49])^(a[326] & b[50])^(a[325] & b[51])^(a[324] & b[52])^(a[323] & b[53])^(a[322] & b[54])^(a[321] & b[55])^(a[320] & b[56])^(a[319] & b[57])^(a[318] & b[58])^(a[317] & b[59])^(a[316] & b[60])^(a[315] & b[61])^(a[314] & b[62])^(a[313] & b[63])^(a[312] & b[64])^(a[311] & b[65])^(a[310] & b[66])^(a[309] & b[67])^(a[308] & b[68])^(a[307] & b[69])^(a[306] & b[70])^(a[305] & b[71])^(a[304] & b[72])^(a[303] & b[73])^(a[302] & b[74])^(a[301] & b[75])^(a[300] & b[76])^(a[299] & b[77])^(a[298] & b[78])^(a[297] & b[79])^(a[296] & b[80])^(a[295] & b[81])^(a[294] & b[82])^(a[293] & b[83])^(a[292] & b[84])^(a[291] & b[85])^(a[290] & b[86])^(a[289] & b[87])^(a[288] & b[88])^(a[287] & b[89])^(a[286] & b[90])^(a[285] & b[91])^(a[284] & b[92])^(a[283] & b[93])^(a[282] & b[94])^(a[281] & b[95])^(a[280] & b[96])^(a[279] & b[97])^(a[278] & b[98])^(a[277] & b[99])^(a[276] & b[100])^(a[275] & b[101])^(a[274] & b[102])^(a[273] & b[103])^(a[272] & b[104])^(a[271] & b[105])^(a[270] & b[106])^(a[269] & b[107])^(a[268] & b[108])^(a[267] & b[109])^(a[266] & b[110])^(a[265] & b[111])^(a[264] & b[112])^(a[263] & b[113])^(a[262] & b[114])^(a[261] & b[115])^(a[260] & b[116])^(a[259] & b[117])^(a[258] & b[118])^(a[257] & b[119])^(a[256] & b[120])^(a[255] & b[121])^(a[254] & b[122])^(a[253] & b[123])^(a[252] & b[124])^(a[251] & b[125])^(a[250] & b[126])^(a[249] & b[127])^(a[248] & b[128])^(a[247] & b[129])^(a[246] & b[130])^(a[245] & b[131])^(a[244] & b[132])^(a[243] & b[133])^(a[242] & b[134])^(a[241] & b[135])^(a[240] & b[136])^(a[239] & b[137])^(a[238] & b[138])^(a[237] & b[139])^(a[236] & b[140])^(a[235] & b[141])^(a[234] & b[142])^(a[233] & b[143])^(a[232] & b[144])^(a[231] & b[145])^(a[230] & b[146])^(a[229] & b[147])^(a[228] & b[148])^(a[227] & b[149])^(a[226] & b[150])^(a[225] & b[151])^(a[224] & b[152])^(a[223] & b[153])^(a[222] & b[154])^(a[221] & b[155])^(a[220] & b[156])^(a[219] & b[157])^(a[218] & b[158])^(a[217] & b[159])^(a[216] & b[160])^(a[215] & b[161])^(a[214] & b[162])^(a[213] & b[163])^(a[212] & b[164])^(a[211] & b[165])^(a[210] & b[166])^(a[209] & b[167])^(a[208] & b[168])^(a[207] & b[169])^(a[206] & b[170])^(a[205] & b[171])^(a[204] & b[172])^(a[203] & b[173])^(a[202] & b[174])^(a[201] & b[175])^(a[200] & b[176])^(a[199] & b[177])^(a[198] & b[178])^(a[197] & b[179])^(a[196] & b[180])^(a[195] & b[181])^(a[194] & b[182])^(a[193] & b[183])^(a[192] & b[184])^(a[191] & b[185])^(a[190] & b[186])^(a[189] & b[187])^(a[188] & b[188])^(a[187] & b[189])^(a[186] & b[190])^(a[185] & b[191])^(a[184] & b[192])^(a[183] & b[193])^(a[182] & b[194])^(a[181] & b[195])^(a[180] & b[196])^(a[179] & b[197])^(a[178] & b[198])^(a[177] & b[199])^(a[176] & b[200])^(a[175] & b[201])^(a[174] & b[202])^(a[173] & b[203])^(a[172] & b[204])^(a[171] & b[205])^(a[170] & b[206])^(a[169] & b[207])^(a[168] & b[208])^(a[167] & b[209])^(a[166] & b[210])^(a[165] & b[211])^(a[164] & b[212])^(a[163] & b[213])^(a[162] & b[214])^(a[161] & b[215])^(a[160] & b[216])^(a[159] & b[217])^(a[158] & b[218])^(a[157] & b[219])^(a[156] & b[220])^(a[155] & b[221])^(a[154] & b[222])^(a[153] & b[223])^(a[152] & b[224])^(a[151] & b[225])^(a[150] & b[226])^(a[149] & b[227])^(a[148] & b[228])^(a[147] & b[229])^(a[146] & b[230])^(a[145] & b[231])^(a[144] & b[232])^(a[143] & b[233])^(a[142] & b[234])^(a[141] & b[235])^(a[140] & b[236])^(a[139] & b[237])^(a[138] & b[238])^(a[137] & b[239])^(a[136] & b[240])^(a[135] & b[241])^(a[134] & b[242])^(a[133] & b[243])^(a[132] & b[244])^(a[131] & b[245])^(a[130] & b[246])^(a[129] & b[247])^(a[128] & b[248])^(a[127] & b[249])^(a[126] & b[250])^(a[125] & b[251])^(a[124] & b[252])^(a[123] & b[253])^(a[122] & b[254])^(a[121] & b[255])^(a[120] & b[256])^(a[119] & b[257])^(a[118] & b[258])^(a[117] & b[259])^(a[116] & b[260])^(a[115] & b[261])^(a[114] & b[262])^(a[113] & b[263])^(a[112] & b[264])^(a[111] & b[265])^(a[110] & b[266])^(a[109] & b[267])^(a[108] & b[268])^(a[107] & b[269])^(a[106] & b[270])^(a[105] & b[271])^(a[104] & b[272])^(a[103] & b[273])^(a[102] & b[274])^(a[101] & b[275])^(a[100] & b[276])^(a[99] & b[277])^(a[98] & b[278])^(a[97] & b[279])^(a[96] & b[280])^(a[95] & b[281])^(a[94] & b[282])^(a[93] & b[283])^(a[92] & b[284])^(a[91] & b[285])^(a[90] & b[286])^(a[89] & b[287])^(a[88] & b[288])^(a[87] & b[289])^(a[86] & b[290])^(a[85] & b[291])^(a[84] & b[292])^(a[83] & b[293])^(a[82] & b[294])^(a[81] & b[295])^(a[80] & b[296])^(a[79] & b[297])^(a[78] & b[298])^(a[77] & b[299])^(a[76] & b[300])^(a[75] & b[301])^(a[74] & b[302])^(a[73] & b[303])^(a[72] & b[304])^(a[71] & b[305])^(a[70] & b[306])^(a[69] & b[307])^(a[68] & b[308])^(a[67] & b[309])^(a[66] & b[310])^(a[65] & b[311])^(a[64] & b[312])^(a[63] & b[313])^(a[62] & b[314])^(a[61] & b[315])^(a[60] & b[316])^(a[59] & b[317])^(a[58] & b[318])^(a[57] & b[319])^(a[56] & b[320])^(a[55] & b[321])^(a[54] & b[322])^(a[53] & b[323])^(a[52] & b[324])^(a[51] & b[325])^(a[50] & b[326])^(a[49] & b[327])^(a[48] & b[328])^(a[47] & b[329])^(a[46] & b[330])^(a[45] & b[331])^(a[44] & b[332])^(a[43] & b[333])^(a[42] & b[334])^(a[41] & b[335])^(a[40] & b[336])^(a[39] & b[337])^(a[38] & b[338])^(a[37] & b[339])^(a[36] & b[340])^(a[35] & b[341])^(a[34] & b[342])^(a[33] & b[343])^(a[32] & b[344])^(a[31] & b[345])^(a[30] & b[346])^(a[29] & b[347])^(a[28] & b[348])^(a[27] & b[349])^(a[26] & b[350])^(a[25] & b[351])^(a[24] & b[352])^(a[23] & b[353])^(a[22] & b[354])^(a[21] & b[355])^(a[20] & b[356])^(a[19] & b[357])^(a[18] & b[358])^(a[17] & b[359])^(a[16] & b[360])^(a[15] & b[361])^(a[14] & b[362])^(a[13] & b[363])^(a[12] & b[364])^(a[11] & b[365])^(a[10] & b[366])^(a[9] & b[367])^(a[8] & b[368])^(a[7] & b[369])^(a[6] & b[370])^(a[5] & b[371])^(a[4] & b[372])^(a[3] & b[373])^(a[2] & b[374])^(a[1] & b[375])^(a[0] & b[376]);
assign y[377] = (a[377] & b[0])^(a[376] & b[1])^(a[375] & b[2])^(a[374] & b[3])^(a[373] & b[4])^(a[372] & b[5])^(a[371] & b[6])^(a[370] & b[7])^(a[369] & b[8])^(a[368] & b[9])^(a[367] & b[10])^(a[366] & b[11])^(a[365] & b[12])^(a[364] & b[13])^(a[363] & b[14])^(a[362] & b[15])^(a[361] & b[16])^(a[360] & b[17])^(a[359] & b[18])^(a[358] & b[19])^(a[357] & b[20])^(a[356] & b[21])^(a[355] & b[22])^(a[354] & b[23])^(a[353] & b[24])^(a[352] & b[25])^(a[351] & b[26])^(a[350] & b[27])^(a[349] & b[28])^(a[348] & b[29])^(a[347] & b[30])^(a[346] & b[31])^(a[345] & b[32])^(a[344] & b[33])^(a[343] & b[34])^(a[342] & b[35])^(a[341] & b[36])^(a[340] & b[37])^(a[339] & b[38])^(a[338] & b[39])^(a[337] & b[40])^(a[336] & b[41])^(a[335] & b[42])^(a[334] & b[43])^(a[333] & b[44])^(a[332] & b[45])^(a[331] & b[46])^(a[330] & b[47])^(a[329] & b[48])^(a[328] & b[49])^(a[327] & b[50])^(a[326] & b[51])^(a[325] & b[52])^(a[324] & b[53])^(a[323] & b[54])^(a[322] & b[55])^(a[321] & b[56])^(a[320] & b[57])^(a[319] & b[58])^(a[318] & b[59])^(a[317] & b[60])^(a[316] & b[61])^(a[315] & b[62])^(a[314] & b[63])^(a[313] & b[64])^(a[312] & b[65])^(a[311] & b[66])^(a[310] & b[67])^(a[309] & b[68])^(a[308] & b[69])^(a[307] & b[70])^(a[306] & b[71])^(a[305] & b[72])^(a[304] & b[73])^(a[303] & b[74])^(a[302] & b[75])^(a[301] & b[76])^(a[300] & b[77])^(a[299] & b[78])^(a[298] & b[79])^(a[297] & b[80])^(a[296] & b[81])^(a[295] & b[82])^(a[294] & b[83])^(a[293] & b[84])^(a[292] & b[85])^(a[291] & b[86])^(a[290] & b[87])^(a[289] & b[88])^(a[288] & b[89])^(a[287] & b[90])^(a[286] & b[91])^(a[285] & b[92])^(a[284] & b[93])^(a[283] & b[94])^(a[282] & b[95])^(a[281] & b[96])^(a[280] & b[97])^(a[279] & b[98])^(a[278] & b[99])^(a[277] & b[100])^(a[276] & b[101])^(a[275] & b[102])^(a[274] & b[103])^(a[273] & b[104])^(a[272] & b[105])^(a[271] & b[106])^(a[270] & b[107])^(a[269] & b[108])^(a[268] & b[109])^(a[267] & b[110])^(a[266] & b[111])^(a[265] & b[112])^(a[264] & b[113])^(a[263] & b[114])^(a[262] & b[115])^(a[261] & b[116])^(a[260] & b[117])^(a[259] & b[118])^(a[258] & b[119])^(a[257] & b[120])^(a[256] & b[121])^(a[255] & b[122])^(a[254] & b[123])^(a[253] & b[124])^(a[252] & b[125])^(a[251] & b[126])^(a[250] & b[127])^(a[249] & b[128])^(a[248] & b[129])^(a[247] & b[130])^(a[246] & b[131])^(a[245] & b[132])^(a[244] & b[133])^(a[243] & b[134])^(a[242] & b[135])^(a[241] & b[136])^(a[240] & b[137])^(a[239] & b[138])^(a[238] & b[139])^(a[237] & b[140])^(a[236] & b[141])^(a[235] & b[142])^(a[234] & b[143])^(a[233] & b[144])^(a[232] & b[145])^(a[231] & b[146])^(a[230] & b[147])^(a[229] & b[148])^(a[228] & b[149])^(a[227] & b[150])^(a[226] & b[151])^(a[225] & b[152])^(a[224] & b[153])^(a[223] & b[154])^(a[222] & b[155])^(a[221] & b[156])^(a[220] & b[157])^(a[219] & b[158])^(a[218] & b[159])^(a[217] & b[160])^(a[216] & b[161])^(a[215] & b[162])^(a[214] & b[163])^(a[213] & b[164])^(a[212] & b[165])^(a[211] & b[166])^(a[210] & b[167])^(a[209] & b[168])^(a[208] & b[169])^(a[207] & b[170])^(a[206] & b[171])^(a[205] & b[172])^(a[204] & b[173])^(a[203] & b[174])^(a[202] & b[175])^(a[201] & b[176])^(a[200] & b[177])^(a[199] & b[178])^(a[198] & b[179])^(a[197] & b[180])^(a[196] & b[181])^(a[195] & b[182])^(a[194] & b[183])^(a[193] & b[184])^(a[192] & b[185])^(a[191] & b[186])^(a[190] & b[187])^(a[189] & b[188])^(a[188] & b[189])^(a[187] & b[190])^(a[186] & b[191])^(a[185] & b[192])^(a[184] & b[193])^(a[183] & b[194])^(a[182] & b[195])^(a[181] & b[196])^(a[180] & b[197])^(a[179] & b[198])^(a[178] & b[199])^(a[177] & b[200])^(a[176] & b[201])^(a[175] & b[202])^(a[174] & b[203])^(a[173] & b[204])^(a[172] & b[205])^(a[171] & b[206])^(a[170] & b[207])^(a[169] & b[208])^(a[168] & b[209])^(a[167] & b[210])^(a[166] & b[211])^(a[165] & b[212])^(a[164] & b[213])^(a[163] & b[214])^(a[162] & b[215])^(a[161] & b[216])^(a[160] & b[217])^(a[159] & b[218])^(a[158] & b[219])^(a[157] & b[220])^(a[156] & b[221])^(a[155] & b[222])^(a[154] & b[223])^(a[153] & b[224])^(a[152] & b[225])^(a[151] & b[226])^(a[150] & b[227])^(a[149] & b[228])^(a[148] & b[229])^(a[147] & b[230])^(a[146] & b[231])^(a[145] & b[232])^(a[144] & b[233])^(a[143] & b[234])^(a[142] & b[235])^(a[141] & b[236])^(a[140] & b[237])^(a[139] & b[238])^(a[138] & b[239])^(a[137] & b[240])^(a[136] & b[241])^(a[135] & b[242])^(a[134] & b[243])^(a[133] & b[244])^(a[132] & b[245])^(a[131] & b[246])^(a[130] & b[247])^(a[129] & b[248])^(a[128] & b[249])^(a[127] & b[250])^(a[126] & b[251])^(a[125] & b[252])^(a[124] & b[253])^(a[123] & b[254])^(a[122] & b[255])^(a[121] & b[256])^(a[120] & b[257])^(a[119] & b[258])^(a[118] & b[259])^(a[117] & b[260])^(a[116] & b[261])^(a[115] & b[262])^(a[114] & b[263])^(a[113] & b[264])^(a[112] & b[265])^(a[111] & b[266])^(a[110] & b[267])^(a[109] & b[268])^(a[108] & b[269])^(a[107] & b[270])^(a[106] & b[271])^(a[105] & b[272])^(a[104] & b[273])^(a[103] & b[274])^(a[102] & b[275])^(a[101] & b[276])^(a[100] & b[277])^(a[99] & b[278])^(a[98] & b[279])^(a[97] & b[280])^(a[96] & b[281])^(a[95] & b[282])^(a[94] & b[283])^(a[93] & b[284])^(a[92] & b[285])^(a[91] & b[286])^(a[90] & b[287])^(a[89] & b[288])^(a[88] & b[289])^(a[87] & b[290])^(a[86] & b[291])^(a[85] & b[292])^(a[84] & b[293])^(a[83] & b[294])^(a[82] & b[295])^(a[81] & b[296])^(a[80] & b[297])^(a[79] & b[298])^(a[78] & b[299])^(a[77] & b[300])^(a[76] & b[301])^(a[75] & b[302])^(a[74] & b[303])^(a[73] & b[304])^(a[72] & b[305])^(a[71] & b[306])^(a[70] & b[307])^(a[69] & b[308])^(a[68] & b[309])^(a[67] & b[310])^(a[66] & b[311])^(a[65] & b[312])^(a[64] & b[313])^(a[63] & b[314])^(a[62] & b[315])^(a[61] & b[316])^(a[60] & b[317])^(a[59] & b[318])^(a[58] & b[319])^(a[57] & b[320])^(a[56] & b[321])^(a[55] & b[322])^(a[54] & b[323])^(a[53] & b[324])^(a[52] & b[325])^(a[51] & b[326])^(a[50] & b[327])^(a[49] & b[328])^(a[48] & b[329])^(a[47] & b[330])^(a[46] & b[331])^(a[45] & b[332])^(a[44] & b[333])^(a[43] & b[334])^(a[42] & b[335])^(a[41] & b[336])^(a[40] & b[337])^(a[39] & b[338])^(a[38] & b[339])^(a[37] & b[340])^(a[36] & b[341])^(a[35] & b[342])^(a[34] & b[343])^(a[33] & b[344])^(a[32] & b[345])^(a[31] & b[346])^(a[30] & b[347])^(a[29] & b[348])^(a[28] & b[349])^(a[27] & b[350])^(a[26] & b[351])^(a[25] & b[352])^(a[24] & b[353])^(a[23] & b[354])^(a[22] & b[355])^(a[21] & b[356])^(a[20] & b[357])^(a[19] & b[358])^(a[18] & b[359])^(a[17] & b[360])^(a[16] & b[361])^(a[15] & b[362])^(a[14] & b[363])^(a[13] & b[364])^(a[12] & b[365])^(a[11] & b[366])^(a[10] & b[367])^(a[9] & b[368])^(a[8] & b[369])^(a[7] & b[370])^(a[6] & b[371])^(a[5] & b[372])^(a[4] & b[373])^(a[3] & b[374])^(a[2] & b[375])^(a[1] & b[376])^(a[0] & b[377]);
assign y[378] = (a[378] & b[0])^(a[377] & b[1])^(a[376] & b[2])^(a[375] & b[3])^(a[374] & b[4])^(a[373] & b[5])^(a[372] & b[6])^(a[371] & b[7])^(a[370] & b[8])^(a[369] & b[9])^(a[368] & b[10])^(a[367] & b[11])^(a[366] & b[12])^(a[365] & b[13])^(a[364] & b[14])^(a[363] & b[15])^(a[362] & b[16])^(a[361] & b[17])^(a[360] & b[18])^(a[359] & b[19])^(a[358] & b[20])^(a[357] & b[21])^(a[356] & b[22])^(a[355] & b[23])^(a[354] & b[24])^(a[353] & b[25])^(a[352] & b[26])^(a[351] & b[27])^(a[350] & b[28])^(a[349] & b[29])^(a[348] & b[30])^(a[347] & b[31])^(a[346] & b[32])^(a[345] & b[33])^(a[344] & b[34])^(a[343] & b[35])^(a[342] & b[36])^(a[341] & b[37])^(a[340] & b[38])^(a[339] & b[39])^(a[338] & b[40])^(a[337] & b[41])^(a[336] & b[42])^(a[335] & b[43])^(a[334] & b[44])^(a[333] & b[45])^(a[332] & b[46])^(a[331] & b[47])^(a[330] & b[48])^(a[329] & b[49])^(a[328] & b[50])^(a[327] & b[51])^(a[326] & b[52])^(a[325] & b[53])^(a[324] & b[54])^(a[323] & b[55])^(a[322] & b[56])^(a[321] & b[57])^(a[320] & b[58])^(a[319] & b[59])^(a[318] & b[60])^(a[317] & b[61])^(a[316] & b[62])^(a[315] & b[63])^(a[314] & b[64])^(a[313] & b[65])^(a[312] & b[66])^(a[311] & b[67])^(a[310] & b[68])^(a[309] & b[69])^(a[308] & b[70])^(a[307] & b[71])^(a[306] & b[72])^(a[305] & b[73])^(a[304] & b[74])^(a[303] & b[75])^(a[302] & b[76])^(a[301] & b[77])^(a[300] & b[78])^(a[299] & b[79])^(a[298] & b[80])^(a[297] & b[81])^(a[296] & b[82])^(a[295] & b[83])^(a[294] & b[84])^(a[293] & b[85])^(a[292] & b[86])^(a[291] & b[87])^(a[290] & b[88])^(a[289] & b[89])^(a[288] & b[90])^(a[287] & b[91])^(a[286] & b[92])^(a[285] & b[93])^(a[284] & b[94])^(a[283] & b[95])^(a[282] & b[96])^(a[281] & b[97])^(a[280] & b[98])^(a[279] & b[99])^(a[278] & b[100])^(a[277] & b[101])^(a[276] & b[102])^(a[275] & b[103])^(a[274] & b[104])^(a[273] & b[105])^(a[272] & b[106])^(a[271] & b[107])^(a[270] & b[108])^(a[269] & b[109])^(a[268] & b[110])^(a[267] & b[111])^(a[266] & b[112])^(a[265] & b[113])^(a[264] & b[114])^(a[263] & b[115])^(a[262] & b[116])^(a[261] & b[117])^(a[260] & b[118])^(a[259] & b[119])^(a[258] & b[120])^(a[257] & b[121])^(a[256] & b[122])^(a[255] & b[123])^(a[254] & b[124])^(a[253] & b[125])^(a[252] & b[126])^(a[251] & b[127])^(a[250] & b[128])^(a[249] & b[129])^(a[248] & b[130])^(a[247] & b[131])^(a[246] & b[132])^(a[245] & b[133])^(a[244] & b[134])^(a[243] & b[135])^(a[242] & b[136])^(a[241] & b[137])^(a[240] & b[138])^(a[239] & b[139])^(a[238] & b[140])^(a[237] & b[141])^(a[236] & b[142])^(a[235] & b[143])^(a[234] & b[144])^(a[233] & b[145])^(a[232] & b[146])^(a[231] & b[147])^(a[230] & b[148])^(a[229] & b[149])^(a[228] & b[150])^(a[227] & b[151])^(a[226] & b[152])^(a[225] & b[153])^(a[224] & b[154])^(a[223] & b[155])^(a[222] & b[156])^(a[221] & b[157])^(a[220] & b[158])^(a[219] & b[159])^(a[218] & b[160])^(a[217] & b[161])^(a[216] & b[162])^(a[215] & b[163])^(a[214] & b[164])^(a[213] & b[165])^(a[212] & b[166])^(a[211] & b[167])^(a[210] & b[168])^(a[209] & b[169])^(a[208] & b[170])^(a[207] & b[171])^(a[206] & b[172])^(a[205] & b[173])^(a[204] & b[174])^(a[203] & b[175])^(a[202] & b[176])^(a[201] & b[177])^(a[200] & b[178])^(a[199] & b[179])^(a[198] & b[180])^(a[197] & b[181])^(a[196] & b[182])^(a[195] & b[183])^(a[194] & b[184])^(a[193] & b[185])^(a[192] & b[186])^(a[191] & b[187])^(a[190] & b[188])^(a[189] & b[189])^(a[188] & b[190])^(a[187] & b[191])^(a[186] & b[192])^(a[185] & b[193])^(a[184] & b[194])^(a[183] & b[195])^(a[182] & b[196])^(a[181] & b[197])^(a[180] & b[198])^(a[179] & b[199])^(a[178] & b[200])^(a[177] & b[201])^(a[176] & b[202])^(a[175] & b[203])^(a[174] & b[204])^(a[173] & b[205])^(a[172] & b[206])^(a[171] & b[207])^(a[170] & b[208])^(a[169] & b[209])^(a[168] & b[210])^(a[167] & b[211])^(a[166] & b[212])^(a[165] & b[213])^(a[164] & b[214])^(a[163] & b[215])^(a[162] & b[216])^(a[161] & b[217])^(a[160] & b[218])^(a[159] & b[219])^(a[158] & b[220])^(a[157] & b[221])^(a[156] & b[222])^(a[155] & b[223])^(a[154] & b[224])^(a[153] & b[225])^(a[152] & b[226])^(a[151] & b[227])^(a[150] & b[228])^(a[149] & b[229])^(a[148] & b[230])^(a[147] & b[231])^(a[146] & b[232])^(a[145] & b[233])^(a[144] & b[234])^(a[143] & b[235])^(a[142] & b[236])^(a[141] & b[237])^(a[140] & b[238])^(a[139] & b[239])^(a[138] & b[240])^(a[137] & b[241])^(a[136] & b[242])^(a[135] & b[243])^(a[134] & b[244])^(a[133] & b[245])^(a[132] & b[246])^(a[131] & b[247])^(a[130] & b[248])^(a[129] & b[249])^(a[128] & b[250])^(a[127] & b[251])^(a[126] & b[252])^(a[125] & b[253])^(a[124] & b[254])^(a[123] & b[255])^(a[122] & b[256])^(a[121] & b[257])^(a[120] & b[258])^(a[119] & b[259])^(a[118] & b[260])^(a[117] & b[261])^(a[116] & b[262])^(a[115] & b[263])^(a[114] & b[264])^(a[113] & b[265])^(a[112] & b[266])^(a[111] & b[267])^(a[110] & b[268])^(a[109] & b[269])^(a[108] & b[270])^(a[107] & b[271])^(a[106] & b[272])^(a[105] & b[273])^(a[104] & b[274])^(a[103] & b[275])^(a[102] & b[276])^(a[101] & b[277])^(a[100] & b[278])^(a[99] & b[279])^(a[98] & b[280])^(a[97] & b[281])^(a[96] & b[282])^(a[95] & b[283])^(a[94] & b[284])^(a[93] & b[285])^(a[92] & b[286])^(a[91] & b[287])^(a[90] & b[288])^(a[89] & b[289])^(a[88] & b[290])^(a[87] & b[291])^(a[86] & b[292])^(a[85] & b[293])^(a[84] & b[294])^(a[83] & b[295])^(a[82] & b[296])^(a[81] & b[297])^(a[80] & b[298])^(a[79] & b[299])^(a[78] & b[300])^(a[77] & b[301])^(a[76] & b[302])^(a[75] & b[303])^(a[74] & b[304])^(a[73] & b[305])^(a[72] & b[306])^(a[71] & b[307])^(a[70] & b[308])^(a[69] & b[309])^(a[68] & b[310])^(a[67] & b[311])^(a[66] & b[312])^(a[65] & b[313])^(a[64] & b[314])^(a[63] & b[315])^(a[62] & b[316])^(a[61] & b[317])^(a[60] & b[318])^(a[59] & b[319])^(a[58] & b[320])^(a[57] & b[321])^(a[56] & b[322])^(a[55] & b[323])^(a[54] & b[324])^(a[53] & b[325])^(a[52] & b[326])^(a[51] & b[327])^(a[50] & b[328])^(a[49] & b[329])^(a[48] & b[330])^(a[47] & b[331])^(a[46] & b[332])^(a[45] & b[333])^(a[44] & b[334])^(a[43] & b[335])^(a[42] & b[336])^(a[41] & b[337])^(a[40] & b[338])^(a[39] & b[339])^(a[38] & b[340])^(a[37] & b[341])^(a[36] & b[342])^(a[35] & b[343])^(a[34] & b[344])^(a[33] & b[345])^(a[32] & b[346])^(a[31] & b[347])^(a[30] & b[348])^(a[29] & b[349])^(a[28] & b[350])^(a[27] & b[351])^(a[26] & b[352])^(a[25] & b[353])^(a[24] & b[354])^(a[23] & b[355])^(a[22] & b[356])^(a[21] & b[357])^(a[20] & b[358])^(a[19] & b[359])^(a[18] & b[360])^(a[17] & b[361])^(a[16] & b[362])^(a[15] & b[363])^(a[14] & b[364])^(a[13] & b[365])^(a[12] & b[366])^(a[11] & b[367])^(a[10] & b[368])^(a[9] & b[369])^(a[8] & b[370])^(a[7] & b[371])^(a[6] & b[372])^(a[5] & b[373])^(a[4] & b[374])^(a[3] & b[375])^(a[2] & b[376])^(a[1] & b[377])^(a[0] & b[378]);
assign y[379] = (a[379] & b[0])^(a[378] & b[1])^(a[377] & b[2])^(a[376] & b[3])^(a[375] & b[4])^(a[374] & b[5])^(a[373] & b[6])^(a[372] & b[7])^(a[371] & b[8])^(a[370] & b[9])^(a[369] & b[10])^(a[368] & b[11])^(a[367] & b[12])^(a[366] & b[13])^(a[365] & b[14])^(a[364] & b[15])^(a[363] & b[16])^(a[362] & b[17])^(a[361] & b[18])^(a[360] & b[19])^(a[359] & b[20])^(a[358] & b[21])^(a[357] & b[22])^(a[356] & b[23])^(a[355] & b[24])^(a[354] & b[25])^(a[353] & b[26])^(a[352] & b[27])^(a[351] & b[28])^(a[350] & b[29])^(a[349] & b[30])^(a[348] & b[31])^(a[347] & b[32])^(a[346] & b[33])^(a[345] & b[34])^(a[344] & b[35])^(a[343] & b[36])^(a[342] & b[37])^(a[341] & b[38])^(a[340] & b[39])^(a[339] & b[40])^(a[338] & b[41])^(a[337] & b[42])^(a[336] & b[43])^(a[335] & b[44])^(a[334] & b[45])^(a[333] & b[46])^(a[332] & b[47])^(a[331] & b[48])^(a[330] & b[49])^(a[329] & b[50])^(a[328] & b[51])^(a[327] & b[52])^(a[326] & b[53])^(a[325] & b[54])^(a[324] & b[55])^(a[323] & b[56])^(a[322] & b[57])^(a[321] & b[58])^(a[320] & b[59])^(a[319] & b[60])^(a[318] & b[61])^(a[317] & b[62])^(a[316] & b[63])^(a[315] & b[64])^(a[314] & b[65])^(a[313] & b[66])^(a[312] & b[67])^(a[311] & b[68])^(a[310] & b[69])^(a[309] & b[70])^(a[308] & b[71])^(a[307] & b[72])^(a[306] & b[73])^(a[305] & b[74])^(a[304] & b[75])^(a[303] & b[76])^(a[302] & b[77])^(a[301] & b[78])^(a[300] & b[79])^(a[299] & b[80])^(a[298] & b[81])^(a[297] & b[82])^(a[296] & b[83])^(a[295] & b[84])^(a[294] & b[85])^(a[293] & b[86])^(a[292] & b[87])^(a[291] & b[88])^(a[290] & b[89])^(a[289] & b[90])^(a[288] & b[91])^(a[287] & b[92])^(a[286] & b[93])^(a[285] & b[94])^(a[284] & b[95])^(a[283] & b[96])^(a[282] & b[97])^(a[281] & b[98])^(a[280] & b[99])^(a[279] & b[100])^(a[278] & b[101])^(a[277] & b[102])^(a[276] & b[103])^(a[275] & b[104])^(a[274] & b[105])^(a[273] & b[106])^(a[272] & b[107])^(a[271] & b[108])^(a[270] & b[109])^(a[269] & b[110])^(a[268] & b[111])^(a[267] & b[112])^(a[266] & b[113])^(a[265] & b[114])^(a[264] & b[115])^(a[263] & b[116])^(a[262] & b[117])^(a[261] & b[118])^(a[260] & b[119])^(a[259] & b[120])^(a[258] & b[121])^(a[257] & b[122])^(a[256] & b[123])^(a[255] & b[124])^(a[254] & b[125])^(a[253] & b[126])^(a[252] & b[127])^(a[251] & b[128])^(a[250] & b[129])^(a[249] & b[130])^(a[248] & b[131])^(a[247] & b[132])^(a[246] & b[133])^(a[245] & b[134])^(a[244] & b[135])^(a[243] & b[136])^(a[242] & b[137])^(a[241] & b[138])^(a[240] & b[139])^(a[239] & b[140])^(a[238] & b[141])^(a[237] & b[142])^(a[236] & b[143])^(a[235] & b[144])^(a[234] & b[145])^(a[233] & b[146])^(a[232] & b[147])^(a[231] & b[148])^(a[230] & b[149])^(a[229] & b[150])^(a[228] & b[151])^(a[227] & b[152])^(a[226] & b[153])^(a[225] & b[154])^(a[224] & b[155])^(a[223] & b[156])^(a[222] & b[157])^(a[221] & b[158])^(a[220] & b[159])^(a[219] & b[160])^(a[218] & b[161])^(a[217] & b[162])^(a[216] & b[163])^(a[215] & b[164])^(a[214] & b[165])^(a[213] & b[166])^(a[212] & b[167])^(a[211] & b[168])^(a[210] & b[169])^(a[209] & b[170])^(a[208] & b[171])^(a[207] & b[172])^(a[206] & b[173])^(a[205] & b[174])^(a[204] & b[175])^(a[203] & b[176])^(a[202] & b[177])^(a[201] & b[178])^(a[200] & b[179])^(a[199] & b[180])^(a[198] & b[181])^(a[197] & b[182])^(a[196] & b[183])^(a[195] & b[184])^(a[194] & b[185])^(a[193] & b[186])^(a[192] & b[187])^(a[191] & b[188])^(a[190] & b[189])^(a[189] & b[190])^(a[188] & b[191])^(a[187] & b[192])^(a[186] & b[193])^(a[185] & b[194])^(a[184] & b[195])^(a[183] & b[196])^(a[182] & b[197])^(a[181] & b[198])^(a[180] & b[199])^(a[179] & b[200])^(a[178] & b[201])^(a[177] & b[202])^(a[176] & b[203])^(a[175] & b[204])^(a[174] & b[205])^(a[173] & b[206])^(a[172] & b[207])^(a[171] & b[208])^(a[170] & b[209])^(a[169] & b[210])^(a[168] & b[211])^(a[167] & b[212])^(a[166] & b[213])^(a[165] & b[214])^(a[164] & b[215])^(a[163] & b[216])^(a[162] & b[217])^(a[161] & b[218])^(a[160] & b[219])^(a[159] & b[220])^(a[158] & b[221])^(a[157] & b[222])^(a[156] & b[223])^(a[155] & b[224])^(a[154] & b[225])^(a[153] & b[226])^(a[152] & b[227])^(a[151] & b[228])^(a[150] & b[229])^(a[149] & b[230])^(a[148] & b[231])^(a[147] & b[232])^(a[146] & b[233])^(a[145] & b[234])^(a[144] & b[235])^(a[143] & b[236])^(a[142] & b[237])^(a[141] & b[238])^(a[140] & b[239])^(a[139] & b[240])^(a[138] & b[241])^(a[137] & b[242])^(a[136] & b[243])^(a[135] & b[244])^(a[134] & b[245])^(a[133] & b[246])^(a[132] & b[247])^(a[131] & b[248])^(a[130] & b[249])^(a[129] & b[250])^(a[128] & b[251])^(a[127] & b[252])^(a[126] & b[253])^(a[125] & b[254])^(a[124] & b[255])^(a[123] & b[256])^(a[122] & b[257])^(a[121] & b[258])^(a[120] & b[259])^(a[119] & b[260])^(a[118] & b[261])^(a[117] & b[262])^(a[116] & b[263])^(a[115] & b[264])^(a[114] & b[265])^(a[113] & b[266])^(a[112] & b[267])^(a[111] & b[268])^(a[110] & b[269])^(a[109] & b[270])^(a[108] & b[271])^(a[107] & b[272])^(a[106] & b[273])^(a[105] & b[274])^(a[104] & b[275])^(a[103] & b[276])^(a[102] & b[277])^(a[101] & b[278])^(a[100] & b[279])^(a[99] & b[280])^(a[98] & b[281])^(a[97] & b[282])^(a[96] & b[283])^(a[95] & b[284])^(a[94] & b[285])^(a[93] & b[286])^(a[92] & b[287])^(a[91] & b[288])^(a[90] & b[289])^(a[89] & b[290])^(a[88] & b[291])^(a[87] & b[292])^(a[86] & b[293])^(a[85] & b[294])^(a[84] & b[295])^(a[83] & b[296])^(a[82] & b[297])^(a[81] & b[298])^(a[80] & b[299])^(a[79] & b[300])^(a[78] & b[301])^(a[77] & b[302])^(a[76] & b[303])^(a[75] & b[304])^(a[74] & b[305])^(a[73] & b[306])^(a[72] & b[307])^(a[71] & b[308])^(a[70] & b[309])^(a[69] & b[310])^(a[68] & b[311])^(a[67] & b[312])^(a[66] & b[313])^(a[65] & b[314])^(a[64] & b[315])^(a[63] & b[316])^(a[62] & b[317])^(a[61] & b[318])^(a[60] & b[319])^(a[59] & b[320])^(a[58] & b[321])^(a[57] & b[322])^(a[56] & b[323])^(a[55] & b[324])^(a[54] & b[325])^(a[53] & b[326])^(a[52] & b[327])^(a[51] & b[328])^(a[50] & b[329])^(a[49] & b[330])^(a[48] & b[331])^(a[47] & b[332])^(a[46] & b[333])^(a[45] & b[334])^(a[44] & b[335])^(a[43] & b[336])^(a[42] & b[337])^(a[41] & b[338])^(a[40] & b[339])^(a[39] & b[340])^(a[38] & b[341])^(a[37] & b[342])^(a[36] & b[343])^(a[35] & b[344])^(a[34] & b[345])^(a[33] & b[346])^(a[32] & b[347])^(a[31] & b[348])^(a[30] & b[349])^(a[29] & b[350])^(a[28] & b[351])^(a[27] & b[352])^(a[26] & b[353])^(a[25] & b[354])^(a[24] & b[355])^(a[23] & b[356])^(a[22] & b[357])^(a[21] & b[358])^(a[20] & b[359])^(a[19] & b[360])^(a[18] & b[361])^(a[17] & b[362])^(a[16] & b[363])^(a[15] & b[364])^(a[14] & b[365])^(a[13] & b[366])^(a[12] & b[367])^(a[11] & b[368])^(a[10] & b[369])^(a[9] & b[370])^(a[8] & b[371])^(a[7] & b[372])^(a[6] & b[373])^(a[5] & b[374])^(a[4] & b[375])^(a[3] & b[376])^(a[2] & b[377])^(a[1] & b[378])^(a[0] & b[379]);
assign y[380] = (a[380] & b[0])^(a[379] & b[1])^(a[378] & b[2])^(a[377] & b[3])^(a[376] & b[4])^(a[375] & b[5])^(a[374] & b[6])^(a[373] & b[7])^(a[372] & b[8])^(a[371] & b[9])^(a[370] & b[10])^(a[369] & b[11])^(a[368] & b[12])^(a[367] & b[13])^(a[366] & b[14])^(a[365] & b[15])^(a[364] & b[16])^(a[363] & b[17])^(a[362] & b[18])^(a[361] & b[19])^(a[360] & b[20])^(a[359] & b[21])^(a[358] & b[22])^(a[357] & b[23])^(a[356] & b[24])^(a[355] & b[25])^(a[354] & b[26])^(a[353] & b[27])^(a[352] & b[28])^(a[351] & b[29])^(a[350] & b[30])^(a[349] & b[31])^(a[348] & b[32])^(a[347] & b[33])^(a[346] & b[34])^(a[345] & b[35])^(a[344] & b[36])^(a[343] & b[37])^(a[342] & b[38])^(a[341] & b[39])^(a[340] & b[40])^(a[339] & b[41])^(a[338] & b[42])^(a[337] & b[43])^(a[336] & b[44])^(a[335] & b[45])^(a[334] & b[46])^(a[333] & b[47])^(a[332] & b[48])^(a[331] & b[49])^(a[330] & b[50])^(a[329] & b[51])^(a[328] & b[52])^(a[327] & b[53])^(a[326] & b[54])^(a[325] & b[55])^(a[324] & b[56])^(a[323] & b[57])^(a[322] & b[58])^(a[321] & b[59])^(a[320] & b[60])^(a[319] & b[61])^(a[318] & b[62])^(a[317] & b[63])^(a[316] & b[64])^(a[315] & b[65])^(a[314] & b[66])^(a[313] & b[67])^(a[312] & b[68])^(a[311] & b[69])^(a[310] & b[70])^(a[309] & b[71])^(a[308] & b[72])^(a[307] & b[73])^(a[306] & b[74])^(a[305] & b[75])^(a[304] & b[76])^(a[303] & b[77])^(a[302] & b[78])^(a[301] & b[79])^(a[300] & b[80])^(a[299] & b[81])^(a[298] & b[82])^(a[297] & b[83])^(a[296] & b[84])^(a[295] & b[85])^(a[294] & b[86])^(a[293] & b[87])^(a[292] & b[88])^(a[291] & b[89])^(a[290] & b[90])^(a[289] & b[91])^(a[288] & b[92])^(a[287] & b[93])^(a[286] & b[94])^(a[285] & b[95])^(a[284] & b[96])^(a[283] & b[97])^(a[282] & b[98])^(a[281] & b[99])^(a[280] & b[100])^(a[279] & b[101])^(a[278] & b[102])^(a[277] & b[103])^(a[276] & b[104])^(a[275] & b[105])^(a[274] & b[106])^(a[273] & b[107])^(a[272] & b[108])^(a[271] & b[109])^(a[270] & b[110])^(a[269] & b[111])^(a[268] & b[112])^(a[267] & b[113])^(a[266] & b[114])^(a[265] & b[115])^(a[264] & b[116])^(a[263] & b[117])^(a[262] & b[118])^(a[261] & b[119])^(a[260] & b[120])^(a[259] & b[121])^(a[258] & b[122])^(a[257] & b[123])^(a[256] & b[124])^(a[255] & b[125])^(a[254] & b[126])^(a[253] & b[127])^(a[252] & b[128])^(a[251] & b[129])^(a[250] & b[130])^(a[249] & b[131])^(a[248] & b[132])^(a[247] & b[133])^(a[246] & b[134])^(a[245] & b[135])^(a[244] & b[136])^(a[243] & b[137])^(a[242] & b[138])^(a[241] & b[139])^(a[240] & b[140])^(a[239] & b[141])^(a[238] & b[142])^(a[237] & b[143])^(a[236] & b[144])^(a[235] & b[145])^(a[234] & b[146])^(a[233] & b[147])^(a[232] & b[148])^(a[231] & b[149])^(a[230] & b[150])^(a[229] & b[151])^(a[228] & b[152])^(a[227] & b[153])^(a[226] & b[154])^(a[225] & b[155])^(a[224] & b[156])^(a[223] & b[157])^(a[222] & b[158])^(a[221] & b[159])^(a[220] & b[160])^(a[219] & b[161])^(a[218] & b[162])^(a[217] & b[163])^(a[216] & b[164])^(a[215] & b[165])^(a[214] & b[166])^(a[213] & b[167])^(a[212] & b[168])^(a[211] & b[169])^(a[210] & b[170])^(a[209] & b[171])^(a[208] & b[172])^(a[207] & b[173])^(a[206] & b[174])^(a[205] & b[175])^(a[204] & b[176])^(a[203] & b[177])^(a[202] & b[178])^(a[201] & b[179])^(a[200] & b[180])^(a[199] & b[181])^(a[198] & b[182])^(a[197] & b[183])^(a[196] & b[184])^(a[195] & b[185])^(a[194] & b[186])^(a[193] & b[187])^(a[192] & b[188])^(a[191] & b[189])^(a[190] & b[190])^(a[189] & b[191])^(a[188] & b[192])^(a[187] & b[193])^(a[186] & b[194])^(a[185] & b[195])^(a[184] & b[196])^(a[183] & b[197])^(a[182] & b[198])^(a[181] & b[199])^(a[180] & b[200])^(a[179] & b[201])^(a[178] & b[202])^(a[177] & b[203])^(a[176] & b[204])^(a[175] & b[205])^(a[174] & b[206])^(a[173] & b[207])^(a[172] & b[208])^(a[171] & b[209])^(a[170] & b[210])^(a[169] & b[211])^(a[168] & b[212])^(a[167] & b[213])^(a[166] & b[214])^(a[165] & b[215])^(a[164] & b[216])^(a[163] & b[217])^(a[162] & b[218])^(a[161] & b[219])^(a[160] & b[220])^(a[159] & b[221])^(a[158] & b[222])^(a[157] & b[223])^(a[156] & b[224])^(a[155] & b[225])^(a[154] & b[226])^(a[153] & b[227])^(a[152] & b[228])^(a[151] & b[229])^(a[150] & b[230])^(a[149] & b[231])^(a[148] & b[232])^(a[147] & b[233])^(a[146] & b[234])^(a[145] & b[235])^(a[144] & b[236])^(a[143] & b[237])^(a[142] & b[238])^(a[141] & b[239])^(a[140] & b[240])^(a[139] & b[241])^(a[138] & b[242])^(a[137] & b[243])^(a[136] & b[244])^(a[135] & b[245])^(a[134] & b[246])^(a[133] & b[247])^(a[132] & b[248])^(a[131] & b[249])^(a[130] & b[250])^(a[129] & b[251])^(a[128] & b[252])^(a[127] & b[253])^(a[126] & b[254])^(a[125] & b[255])^(a[124] & b[256])^(a[123] & b[257])^(a[122] & b[258])^(a[121] & b[259])^(a[120] & b[260])^(a[119] & b[261])^(a[118] & b[262])^(a[117] & b[263])^(a[116] & b[264])^(a[115] & b[265])^(a[114] & b[266])^(a[113] & b[267])^(a[112] & b[268])^(a[111] & b[269])^(a[110] & b[270])^(a[109] & b[271])^(a[108] & b[272])^(a[107] & b[273])^(a[106] & b[274])^(a[105] & b[275])^(a[104] & b[276])^(a[103] & b[277])^(a[102] & b[278])^(a[101] & b[279])^(a[100] & b[280])^(a[99] & b[281])^(a[98] & b[282])^(a[97] & b[283])^(a[96] & b[284])^(a[95] & b[285])^(a[94] & b[286])^(a[93] & b[287])^(a[92] & b[288])^(a[91] & b[289])^(a[90] & b[290])^(a[89] & b[291])^(a[88] & b[292])^(a[87] & b[293])^(a[86] & b[294])^(a[85] & b[295])^(a[84] & b[296])^(a[83] & b[297])^(a[82] & b[298])^(a[81] & b[299])^(a[80] & b[300])^(a[79] & b[301])^(a[78] & b[302])^(a[77] & b[303])^(a[76] & b[304])^(a[75] & b[305])^(a[74] & b[306])^(a[73] & b[307])^(a[72] & b[308])^(a[71] & b[309])^(a[70] & b[310])^(a[69] & b[311])^(a[68] & b[312])^(a[67] & b[313])^(a[66] & b[314])^(a[65] & b[315])^(a[64] & b[316])^(a[63] & b[317])^(a[62] & b[318])^(a[61] & b[319])^(a[60] & b[320])^(a[59] & b[321])^(a[58] & b[322])^(a[57] & b[323])^(a[56] & b[324])^(a[55] & b[325])^(a[54] & b[326])^(a[53] & b[327])^(a[52] & b[328])^(a[51] & b[329])^(a[50] & b[330])^(a[49] & b[331])^(a[48] & b[332])^(a[47] & b[333])^(a[46] & b[334])^(a[45] & b[335])^(a[44] & b[336])^(a[43] & b[337])^(a[42] & b[338])^(a[41] & b[339])^(a[40] & b[340])^(a[39] & b[341])^(a[38] & b[342])^(a[37] & b[343])^(a[36] & b[344])^(a[35] & b[345])^(a[34] & b[346])^(a[33] & b[347])^(a[32] & b[348])^(a[31] & b[349])^(a[30] & b[350])^(a[29] & b[351])^(a[28] & b[352])^(a[27] & b[353])^(a[26] & b[354])^(a[25] & b[355])^(a[24] & b[356])^(a[23] & b[357])^(a[22] & b[358])^(a[21] & b[359])^(a[20] & b[360])^(a[19] & b[361])^(a[18] & b[362])^(a[17] & b[363])^(a[16] & b[364])^(a[15] & b[365])^(a[14] & b[366])^(a[13] & b[367])^(a[12] & b[368])^(a[11] & b[369])^(a[10] & b[370])^(a[9] & b[371])^(a[8] & b[372])^(a[7] & b[373])^(a[6] & b[374])^(a[5] & b[375])^(a[4] & b[376])^(a[3] & b[377])^(a[2] & b[378])^(a[1] & b[379])^(a[0] & b[380]);
assign y[381] = (a[381] & b[0])^(a[380] & b[1])^(a[379] & b[2])^(a[378] & b[3])^(a[377] & b[4])^(a[376] & b[5])^(a[375] & b[6])^(a[374] & b[7])^(a[373] & b[8])^(a[372] & b[9])^(a[371] & b[10])^(a[370] & b[11])^(a[369] & b[12])^(a[368] & b[13])^(a[367] & b[14])^(a[366] & b[15])^(a[365] & b[16])^(a[364] & b[17])^(a[363] & b[18])^(a[362] & b[19])^(a[361] & b[20])^(a[360] & b[21])^(a[359] & b[22])^(a[358] & b[23])^(a[357] & b[24])^(a[356] & b[25])^(a[355] & b[26])^(a[354] & b[27])^(a[353] & b[28])^(a[352] & b[29])^(a[351] & b[30])^(a[350] & b[31])^(a[349] & b[32])^(a[348] & b[33])^(a[347] & b[34])^(a[346] & b[35])^(a[345] & b[36])^(a[344] & b[37])^(a[343] & b[38])^(a[342] & b[39])^(a[341] & b[40])^(a[340] & b[41])^(a[339] & b[42])^(a[338] & b[43])^(a[337] & b[44])^(a[336] & b[45])^(a[335] & b[46])^(a[334] & b[47])^(a[333] & b[48])^(a[332] & b[49])^(a[331] & b[50])^(a[330] & b[51])^(a[329] & b[52])^(a[328] & b[53])^(a[327] & b[54])^(a[326] & b[55])^(a[325] & b[56])^(a[324] & b[57])^(a[323] & b[58])^(a[322] & b[59])^(a[321] & b[60])^(a[320] & b[61])^(a[319] & b[62])^(a[318] & b[63])^(a[317] & b[64])^(a[316] & b[65])^(a[315] & b[66])^(a[314] & b[67])^(a[313] & b[68])^(a[312] & b[69])^(a[311] & b[70])^(a[310] & b[71])^(a[309] & b[72])^(a[308] & b[73])^(a[307] & b[74])^(a[306] & b[75])^(a[305] & b[76])^(a[304] & b[77])^(a[303] & b[78])^(a[302] & b[79])^(a[301] & b[80])^(a[300] & b[81])^(a[299] & b[82])^(a[298] & b[83])^(a[297] & b[84])^(a[296] & b[85])^(a[295] & b[86])^(a[294] & b[87])^(a[293] & b[88])^(a[292] & b[89])^(a[291] & b[90])^(a[290] & b[91])^(a[289] & b[92])^(a[288] & b[93])^(a[287] & b[94])^(a[286] & b[95])^(a[285] & b[96])^(a[284] & b[97])^(a[283] & b[98])^(a[282] & b[99])^(a[281] & b[100])^(a[280] & b[101])^(a[279] & b[102])^(a[278] & b[103])^(a[277] & b[104])^(a[276] & b[105])^(a[275] & b[106])^(a[274] & b[107])^(a[273] & b[108])^(a[272] & b[109])^(a[271] & b[110])^(a[270] & b[111])^(a[269] & b[112])^(a[268] & b[113])^(a[267] & b[114])^(a[266] & b[115])^(a[265] & b[116])^(a[264] & b[117])^(a[263] & b[118])^(a[262] & b[119])^(a[261] & b[120])^(a[260] & b[121])^(a[259] & b[122])^(a[258] & b[123])^(a[257] & b[124])^(a[256] & b[125])^(a[255] & b[126])^(a[254] & b[127])^(a[253] & b[128])^(a[252] & b[129])^(a[251] & b[130])^(a[250] & b[131])^(a[249] & b[132])^(a[248] & b[133])^(a[247] & b[134])^(a[246] & b[135])^(a[245] & b[136])^(a[244] & b[137])^(a[243] & b[138])^(a[242] & b[139])^(a[241] & b[140])^(a[240] & b[141])^(a[239] & b[142])^(a[238] & b[143])^(a[237] & b[144])^(a[236] & b[145])^(a[235] & b[146])^(a[234] & b[147])^(a[233] & b[148])^(a[232] & b[149])^(a[231] & b[150])^(a[230] & b[151])^(a[229] & b[152])^(a[228] & b[153])^(a[227] & b[154])^(a[226] & b[155])^(a[225] & b[156])^(a[224] & b[157])^(a[223] & b[158])^(a[222] & b[159])^(a[221] & b[160])^(a[220] & b[161])^(a[219] & b[162])^(a[218] & b[163])^(a[217] & b[164])^(a[216] & b[165])^(a[215] & b[166])^(a[214] & b[167])^(a[213] & b[168])^(a[212] & b[169])^(a[211] & b[170])^(a[210] & b[171])^(a[209] & b[172])^(a[208] & b[173])^(a[207] & b[174])^(a[206] & b[175])^(a[205] & b[176])^(a[204] & b[177])^(a[203] & b[178])^(a[202] & b[179])^(a[201] & b[180])^(a[200] & b[181])^(a[199] & b[182])^(a[198] & b[183])^(a[197] & b[184])^(a[196] & b[185])^(a[195] & b[186])^(a[194] & b[187])^(a[193] & b[188])^(a[192] & b[189])^(a[191] & b[190])^(a[190] & b[191])^(a[189] & b[192])^(a[188] & b[193])^(a[187] & b[194])^(a[186] & b[195])^(a[185] & b[196])^(a[184] & b[197])^(a[183] & b[198])^(a[182] & b[199])^(a[181] & b[200])^(a[180] & b[201])^(a[179] & b[202])^(a[178] & b[203])^(a[177] & b[204])^(a[176] & b[205])^(a[175] & b[206])^(a[174] & b[207])^(a[173] & b[208])^(a[172] & b[209])^(a[171] & b[210])^(a[170] & b[211])^(a[169] & b[212])^(a[168] & b[213])^(a[167] & b[214])^(a[166] & b[215])^(a[165] & b[216])^(a[164] & b[217])^(a[163] & b[218])^(a[162] & b[219])^(a[161] & b[220])^(a[160] & b[221])^(a[159] & b[222])^(a[158] & b[223])^(a[157] & b[224])^(a[156] & b[225])^(a[155] & b[226])^(a[154] & b[227])^(a[153] & b[228])^(a[152] & b[229])^(a[151] & b[230])^(a[150] & b[231])^(a[149] & b[232])^(a[148] & b[233])^(a[147] & b[234])^(a[146] & b[235])^(a[145] & b[236])^(a[144] & b[237])^(a[143] & b[238])^(a[142] & b[239])^(a[141] & b[240])^(a[140] & b[241])^(a[139] & b[242])^(a[138] & b[243])^(a[137] & b[244])^(a[136] & b[245])^(a[135] & b[246])^(a[134] & b[247])^(a[133] & b[248])^(a[132] & b[249])^(a[131] & b[250])^(a[130] & b[251])^(a[129] & b[252])^(a[128] & b[253])^(a[127] & b[254])^(a[126] & b[255])^(a[125] & b[256])^(a[124] & b[257])^(a[123] & b[258])^(a[122] & b[259])^(a[121] & b[260])^(a[120] & b[261])^(a[119] & b[262])^(a[118] & b[263])^(a[117] & b[264])^(a[116] & b[265])^(a[115] & b[266])^(a[114] & b[267])^(a[113] & b[268])^(a[112] & b[269])^(a[111] & b[270])^(a[110] & b[271])^(a[109] & b[272])^(a[108] & b[273])^(a[107] & b[274])^(a[106] & b[275])^(a[105] & b[276])^(a[104] & b[277])^(a[103] & b[278])^(a[102] & b[279])^(a[101] & b[280])^(a[100] & b[281])^(a[99] & b[282])^(a[98] & b[283])^(a[97] & b[284])^(a[96] & b[285])^(a[95] & b[286])^(a[94] & b[287])^(a[93] & b[288])^(a[92] & b[289])^(a[91] & b[290])^(a[90] & b[291])^(a[89] & b[292])^(a[88] & b[293])^(a[87] & b[294])^(a[86] & b[295])^(a[85] & b[296])^(a[84] & b[297])^(a[83] & b[298])^(a[82] & b[299])^(a[81] & b[300])^(a[80] & b[301])^(a[79] & b[302])^(a[78] & b[303])^(a[77] & b[304])^(a[76] & b[305])^(a[75] & b[306])^(a[74] & b[307])^(a[73] & b[308])^(a[72] & b[309])^(a[71] & b[310])^(a[70] & b[311])^(a[69] & b[312])^(a[68] & b[313])^(a[67] & b[314])^(a[66] & b[315])^(a[65] & b[316])^(a[64] & b[317])^(a[63] & b[318])^(a[62] & b[319])^(a[61] & b[320])^(a[60] & b[321])^(a[59] & b[322])^(a[58] & b[323])^(a[57] & b[324])^(a[56] & b[325])^(a[55] & b[326])^(a[54] & b[327])^(a[53] & b[328])^(a[52] & b[329])^(a[51] & b[330])^(a[50] & b[331])^(a[49] & b[332])^(a[48] & b[333])^(a[47] & b[334])^(a[46] & b[335])^(a[45] & b[336])^(a[44] & b[337])^(a[43] & b[338])^(a[42] & b[339])^(a[41] & b[340])^(a[40] & b[341])^(a[39] & b[342])^(a[38] & b[343])^(a[37] & b[344])^(a[36] & b[345])^(a[35] & b[346])^(a[34] & b[347])^(a[33] & b[348])^(a[32] & b[349])^(a[31] & b[350])^(a[30] & b[351])^(a[29] & b[352])^(a[28] & b[353])^(a[27] & b[354])^(a[26] & b[355])^(a[25] & b[356])^(a[24] & b[357])^(a[23] & b[358])^(a[22] & b[359])^(a[21] & b[360])^(a[20] & b[361])^(a[19] & b[362])^(a[18] & b[363])^(a[17] & b[364])^(a[16] & b[365])^(a[15] & b[366])^(a[14] & b[367])^(a[13] & b[368])^(a[12] & b[369])^(a[11] & b[370])^(a[10] & b[371])^(a[9] & b[372])^(a[8] & b[373])^(a[7] & b[374])^(a[6] & b[375])^(a[5] & b[376])^(a[4] & b[377])^(a[3] & b[378])^(a[2] & b[379])^(a[1] & b[380])^(a[0] & b[381]);
assign y[382] = (a[382] & b[0])^(a[381] & b[1])^(a[380] & b[2])^(a[379] & b[3])^(a[378] & b[4])^(a[377] & b[5])^(a[376] & b[6])^(a[375] & b[7])^(a[374] & b[8])^(a[373] & b[9])^(a[372] & b[10])^(a[371] & b[11])^(a[370] & b[12])^(a[369] & b[13])^(a[368] & b[14])^(a[367] & b[15])^(a[366] & b[16])^(a[365] & b[17])^(a[364] & b[18])^(a[363] & b[19])^(a[362] & b[20])^(a[361] & b[21])^(a[360] & b[22])^(a[359] & b[23])^(a[358] & b[24])^(a[357] & b[25])^(a[356] & b[26])^(a[355] & b[27])^(a[354] & b[28])^(a[353] & b[29])^(a[352] & b[30])^(a[351] & b[31])^(a[350] & b[32])^(a[349] & b[33])^(a[348] & b[34])^(a[347] & b[35])^(a[346] & b[36])^(a[345] & b[37])^(a[344] & b[38])^(a[343] & b[39])^(a[342] & b[40])^(a[341] & b[41])^(a[340] & b[42])^(a[339] & b[43])^(a[338] & b[44])^(a[337] & b[45])^(a[336] & b[46])^(a[335] & b[47])^(a[334] & b[48])^(a[333] & b[49])^(a[332] & b[50])^(a[331] & b[51])^(a[330] & b[52])^(a[329] & b[53])^(a[328] & b[54])^(a[327] & b[55])^(a[326] & b[56])^(a[325] & b[57])^(a[324] & b[58])^(a[323] & b[59])^(a[322] & b[60])^(a[321] & b[61])^(a[320] & b[62])^(a[319] & b[63])^(a[318] & b[64])^(a[317] & b[65])^(a[316] & b[66])^(a[315] & b[67])^(a[314] & b[68])^(a[313] & b[69])^(a[312] & b[70])^(a[311] & b[71])^(a[310] & b[72])^(a[309] & b[73])^(a[308] & b[74])^(a[307] & b[75])^(a[306] & b[76])^(a[305] & b[77])^(a[304] & b[78])^(a[303] & b[79])^(a[302] & b[80])^(a[301] & b[81])^(a[300] & b[82])^(a[299] & b[83])^(a[298] & b[84])^(a[297] & b[85])^(a[296] & b[86])^(a[295] & b[87])^(a[294] & b[88])^(a[293] & b[89])^(a[292] & b[90])^(a[291] & b[91])^(a[290] & b[92])^(a[289] & b[93])^(a[288] & b[94])^(a[287] & b[95])^(a[286] & b[96])^(a[285] & b[97])^(a[284] & b[98])^(a[283] & b[99])^(a[282] & b[100])^(a[281] & b[101])^(a[280] & b[102])^(a[279] & b[103])^(a[278] & b[104])^(a[277] & b[105])^(a[276] & b[106])^(a[275] & b[107])^(a[274] & b[108])^(a[273] & b[109])^(a[272] & b[110])^(a[271] & b[111])^(a[270] & b[112])^(a[269] & b[113])^(a[268] & b[114])^(a[267] & b[115])^(a[266] & b[116])^(a[265] & b[117])^(a[264] & b[118])^(a[263] & b[119])^(a[262] & b[120])^(a[261] & b[121])^(a[260] & b[122])^(a[259] & b[123])^(a[258] & b[124])^(a[257] & b[125])^(a[256] & b[126])^(a[255] & b[127])^(a[254] & b[128])^(a[253] & b[129])^(a[252] & b[130])^(a[251] & b[131])^(a[250] & b[132])^(a[249] & b[133])^(a[248] & b[134])^(a[247] & b[135])^(a[246] & b[136])^(a[245] & b[137])^(a[244] & b[138])^(a[243] & b[139])^(a[242] & b[140])^(a[241] & b[141])^(a[240] & b[142])^(a[239] & b[143])^(a[238] & b[144])^(a[237] & b[145])^(a[236] & b[146])^(a[235] & b[147])^(a[234] & b[148])^(a[233] & b[149])^(a[232] & b[150])^(a[231] & b[151])^(a[230] & b[152])^(a[229] & b[153])^(a[228] & b[154])^(a[227] & b[155])^(a[226] & b[156])^(a[225] & b[157])^(a[224] & b[158])^(a[223] & b[159])^(a[222] & b[160])^(a[221] & b[161])^(a[220] & b[162])^(a[219] & b[163])^(a[218] & b[164])^(a[217] & b[165])^(a[216] & b[166])^(a[215] & b[167])^(a[214] & b[168])^(a[213] & b[169])^(a[212] & b[170])^(a[211] & b[171])^(a[210] & b[172])^(a[209] & b[173])^(a[208] & b[174])^(a[207] & b[175])^(a[206] & b[176])^(a[205] & b[177])^(a[204] & b[178])^(a[203] & b[179])^(a[202] & b[180])^(a[201] & b[181])^(a[200] & b[182])^(a[199] & b[183])^(a[198] & b[184])^(a[197] & b[185])^(a[196] & b[186])^(a[195] & b[187])^(a[194] & b[188])^(a[193] & b[189])^(a[192] & b[190])^(a[191] & b[191])^(a[190] & b[192])^(a[189] & b[193])^(a[188] & b[194])^(a[187] & b[195])^(a[186] & b[196])^(a[185] & b[197])^(a[184] & b[198])^(a[183] & b[199])^(a[182] & b[200])^(a[181] & b[201])^(a[180] & b[202])^(a[179] & b[203])^(a[178] & b[204])^(a[177] & b[205])^(a[176] & b[206])^(a[175] & b[207])^(a[174] & b[208])^(a[173] & b[209])^(a[172] & b[210])^(a[171] & b[211])^(a[170] & b[212])^(a[169] & b[213])^(a[168] & b[214])^(a[167] & b[215])^(a[166] & b[216])^(a[165] & b[217])^(a[164] & b[218])^(a[163] & b[219])^(a[162] & b[220])^(a[161] & b[221])^(a[160] & b[222])^(a[159] & b[223])^(a[158] & b[224])^(a[157] & b[225])^(a[156] & b[226])^(a[155] & b[227])^(a[154] & b[228])^(a[153] & b[229])^(a[152] & b[230])^(a[151] & b[231])^(a[150] & b[232])^(a[149] & b[233])^(a[148] & b[234])^(a[147] & b[235])^(a[146] & b[236])^(a[145] & b[237])^(a[144] & b[238])^(a[143] & b[239])^(a[142] & b[240])^(a[141] & b[241])^(a[140] & b[242])^(a[139] & b[243])^(a[138] & b[244])^(a[137] & b[245])^(a[136] & b[246])^(a[135] & b[247])^(a[134] & b[248])^(a[133] & b[249])^(a[132] & b[250])^(a[131] & b[251])^(a[130] & b[252])^(a[129] & b[253])^(a[128] & b[254])^(a[127] & b[255])^(a[126] & b[256])^(a[125] & b[257])^(a[124] & b[258])^(a[123] & b[259])^(a[122] & b[260])^(a[121] & b[261])^(a[120] & b[262])^(a[119] & b[263])^(a[118] & b[264])^(a[117] & b[265])^(a[116] & b[266])^(a[115] & b[267])^(a[114] & b[268])^(a[113] & b[269])^(a[112] & b[270])^(a[111] & b[271])^(a[110] & b[272])^(a[109] & b[273])^(a[108] & b[274])^(a[107] & b[275])^(a[106] & b[276])^(a[105] & b[277])^(a[104] & b[278])^(a[103] & b[279])^(a[102] & b[280])^(a[101] & b[281])^(a[100] & b[282])^(a[99] & b[283])^(a[98] & b[284])^(a[97] & b[285])^(a[96] & b[286])^(a[95] & b[287])^(a[94] & b[288])^(a[93] & b[289])^(a[92] & b[290])^(a[91] & b[291])^(a[90] & b[292])^(a[89] & b[293])^(a[88] & b[294])^(a[87] & b[295])^(a[86] & b[296])^(a[85] & b[297])^(a[84] & b[298])^(a[83] & b[299])^(a[82] & b[300])^(a[81] & b[301])^(a[80] & b[302])^(a[79] & b[303])^(a[78] & b[304])^(a[77] & b[305])^(a[76] & b[306])^(a[75] & b[307])^(a[74] & b[308])^(a[73] & b[309])^(a[72] & b[310])^(a[71] & b[311])^(a[70] & b[312])^(a[69] & b[313])^(a[68] & b[314])^(a[67] & b[315])^(a[66] & b[316])^(a[65] & b[317])^(a[64] & b[318])^(a[63] & b[319])^(a[62] & b[320])^(a[61] & b[321])^(a[60] & b[322])^(a[59] & b[323])^(a[58] & b[324])^(a[57] & b[325])^(a[56] & b[326])^(a[55] & b[327])^(a[54] & b[328])^(a[53] & b[329])^(a[52] & b[330])^(a[51] & b[331])^(a[50] & b[332])^(a[49] & b[333])^(a[48] & b[334])^(a[47] & b[335])^(a[46] & b[336])^(a[45] & b[337])^(a[44] & b[338])^(a[43] & b[339])^(a[42] & b[340])^(a[41] & b[341])^(a[40] & b[342])^(a[39] & b[343])^(a[38] & b[344])^(a[37] & b[345])^(a[36] & b[346])^(a[35] & b[347])^(a[34] & b[348])^(a[33] & b[349])^(a[32] & b[350])^(a[31] & b[351])^(a[30] & b[352])^(a[29] & b[353])^(a[28] & b[354])^(a[27] & b[355])^(a[26] & b[356])^(a[25] & b[357])^(a[24] & b[358])^(a[23] & b[359])^(a[22] & b[360])^(a[21] & b[361])^(a[20] & b[362])^(a[19] & b[363])^(a[18] & b[364])^(a[17] & b[365])^(a[16] & b[366])^(a[15] & b[367])^(a[14] & b[368])^(a[13] & b[369])^(a[12] & b[370])^(a[11] & b[371])^(a[10] & b[372])^(a[9] & b[373])^(a[8] & b[374])^(a[7] & b[375])^(a[6] & b[376])^(a[5] & b[377])^(a[4] & b[378])^(a[3] & b[379])^(a[2] & b[380])^(a[1] & b[381])^(a[0] & b[382]);
assign y[383] = (a[383] & b[0])^(a[382] & b[1])^(a[381] & b[2])^(a[380] & b[3])^(a[379] & b[4])^(a[378] & b[5])^(a[377] & b[6])^(a[376] & b[7])^(a[375] & b[8])^(a[374] & b[9])^(a[373] & b[10])^(a[372] & b[11])^(a[371] & b[12])^(a[370] & b[13])^(a[369] & b[14])^(a[368] & b[15])^(a[367] & b[16])^(a[366] & b[17])^(a[365] & b[18])^(a[364] & b[19])^(a[363] & b[20])^(a[362] & b[21])^(a[361] & b[22])^(a[360] & b[23])^(a[359] & b[24])^(a[358] & b[25])^(a[357] & b[26])^(a[356] & b[27])^(a[355] & b[28])^(a[354] & b[29])^(a[353] & b[30])^(a[352] & b[31])^(a[351] & b[32])^(a[350] & b[33])^(a[349] & b[34])^(a[348] & b[35])^(a[347] & b[36])^(a[346] & b[37])^(a[345] & b[38])^(a[344] & b[39])^(a[343] & b[40])^(a[342] & b[41])^(a[341] & b[42])^(a[340] & b[43])^(a[339] & b[44])^(a[338] & b[45])^(a[337] & b[46])^(a[336] & b[47])^(a[335] & b[48])^(a[334] & b[49])^(a[333] & b[50])^(a[332] & b[51])^(a[331] & b[52])^(a[330] & b[53])^(a[329] & b[54])^(a[328] & b[55])^(a[327] & b[56])^(a[326] & b[57])^(a[325] & b[58])^(a[324] & b[59])^(a[323] & b[60])^(a[322] & b[61])^(a[321] & b[62])^(a[320] & b[63])^(a[319] & b[64])^(a[318] & b[65])^(a[317] & b[66])^(a[316] & b[67])^(a[315] & b[68])^(a[314] & b[69])^(a[313] & b[70])^(a[312] & b[71])^(a[311] & b[72])^(a[310] & b[73])^(a[309] & b[74])^(a[308] & b[75])^(a[307] & b[76])^(a[306] & b[77])^(a[305] & b[78])^(a[304] & b[79])^(a[303] & b[80])^(a[302] & b[81])^(a[301] & b[82])^(a[300] & b[83])^(a[299] & b[84])^(a[298] & b[85])^(a[297] & b[86])^(a[296] & b[87])^(a[295] & b[88])^(a[294] & b[89])^(a[293] & b[90])^(a[292] & b[91])^(a[291] & b[92])^(a[290] & b[93])^(a[289] & b[94])^(a[288] & b[95])^(a[287] & b[96])^(a[286] & b[97])^(a[285] & b[98])^(a[284] & b[99])^(a[283] & b[100])^(a[282] & b[101])^(a[281] & b[102])^(a[280] & b[103])^(a[279] & b[104])^(a[278] & b[105])^(a[277] & b[106])^(a[276] & b[107])^(a[275] & b[108])^(a[274] & b[109])^(a[273] & b[110])^(a[272] & b[111])^(a[271] & b[112])^(a[270] & b[113])^(a[269] & b[114])^(a[268] & b[115])^(a[267] & b[116])^(a[266] & b[117])^(a[265] & b[118])^(a[264] & b[119])^(a[263] & b[120])^(a[262] & b[121])^(a[261] & b[122])^(a[260] & b[123])^(a[259] & b[124])^(a[258] & b[125])^(a[257] & b[126])^(a[256] & b[127])^(a[255] & b[128])^(a[254] & b[129])^(a[253] & b[130])^(a[252] & b[131])^(a[251] & b[132])^(a[250] & b[133])^(a[249] & b[134])^(a[248] & b[135])^(a[247] & b[136])^(a[246] & b[137])^(a[245] & b[138])^(a[244] & b[139])^(a[243] & b[140])^(a[242] & b[141])^(a[241] & b[142])^(a[240] & b[143])^(a[239] & b[144])^(a[238] & b[145])^(a[237] & b[146])^(a[236] & b[147])^(a[235] & b[148])^(a[234] & b[149])^(a[233] & b[150])^(a[232] & b[151])^(a[231] & b[152])^(a[230] & b[153])^(a[229] & b[154])^(a[228] & b[155])^(a[227] & b[156])^(a[226] & b[157])^(a[225] & b[158])^(a[224] & b[159])^(a[223] & b[160])^(a[222] & b[161])^(a[221] & b[162])^(a[220] & b[163])^(a[219] & b[164])^(a[218] & b[165])^(a[217] & b[166])^(a[216] & b[167])^(a[215] & b[168])^(a[214] & b[169])^(a[213] & b[170])^(a[212] & b[171])^(a[211] & b[172])^(a[210] & b[173])^(a[209] & b[174])^(a[208] & b[175])^(a[207] & b[176])^(a[206] & b[177])^(a[205] & b[178])^(a[204] & b[179])^(a[203] & b[180])^(a[202] & b[181])^(a[201] & b[182])^(a[200] & b[183])^(a[199] & b[184])^(a[198] & b[185])^(a[197] & b[186])^(a[196] & b[187])^(a[195] & b[188])^(a[194] & b[189])^(a[193] & b[190])^(a[192] & b[191])^(a[191] & b[192])^(a[190] & b[193])^(a[189] & b[194])^(a[188] & b[195])^(a[187] & b[196])^(a[186] & b[197])^(a[185] & b[198])^(a[184] & b[199])^(a[183] & b[200])^(a[182] & b[201])^(a[181] & b[202])^(a[180] & b[203])^(a[179] & b[204])^(a[178] & b[205])^(a[177] & b[206])^(a[176] & b[207])^(a[175] & b[208])^(a[174] & b[209])^(a[173] & b[210])^(a[172] & b[211])^(a[171] & b[212])^(a[170] & b[213])^(a[169] & b[214])^(a[168] & b[215])^(a[167] & b[216])^(a[166] & b[217])^(a[165] & b[218])^(a[164] & b[219])^(a[163] & b[220])^(a[162] & b[221])^(a[161] & b[222])^(a[160] & b[223])^(a[159] & b[224])^(a[158] & b[225])^(a[157] & b[226])^(a[156] & b[227])^(a[155] & b[228])^(a[154] & b[229])^(a[153] & b[230])^(a[152] & b[231])^(a[151] & b[232])^(a[150] & b[233])^(a[149] & b[234])^(a[148] & b[235])^(a[147] & b[236])^(a[146] & b[237])^(a[145] & b[238])^(a[144] & b[239])^(a[143] & b[240])^(a[142] & b[241])^(a[141] & b[242])^(a[140] & b[243])^(a[139] & b[244])^(a[138] & b[245])^(a[137] & b[246])^(a[136] & b[247])^(a[135] & b[248])^(a[134] & b[249])^(a[133] & b[250])^(a[132] & b[251])^(a[131] & b[252])^(a[130] & b[253])^(a[129] & b[254])^(a[128] & b[255])^(a[127] & b[256])^(a[126] & b[257])^(a[125] & b[258])^(a[124] & b[259])^(a[123] & b[260])^(a[122] & b[261])^(a[121] & b[262])^(a[120] & b[263])^(a[119] & b[264])^(a[118] & b[265])^(a[117] & b[266])^(a[116] & b[267])^(a[115] & b[268])^(a[114] & b[269])^(a[113] & b[270])^(a[112] & b[271])^(a[111] & b[272])^(a[110] & b[273])^(a[109] & b[274])^(a[108] & b[275])^(a[107] & b[276])^(a[106] & b[277])^(a[105] & b[278])^(a[104] & b[279])^(a[103] & b[280])^(a[102] & b[281])^(a[101] & b[282])^(a[100] & b[283])^(a[99] & b[284])^(a[98] & b[285])^(a[97] & b[286])^(a[96] & b[287])^(a[95] & b[288])^(a[94] & b[289])^(a[93] & b[290])^(a[92] & b[291])^(a[91] & b[292])^(a[90] & b[293])^(a[89] & b[294])^(a[88] & b[295])^(a[87] & b[296])^(a[86] & b[297])^(a[85] & b[298])^(a[84] & b[299])^(a[83] & b[300])^(a[82] & b[301])^(a[81] & b[302])^(a[80] & b[303])^(a[79] & b[304])^(a[78] & b[305])^(a[77] & b[306])^(a[76] & b[307])^(a[75] & b[308])^(a[74] & b[309])^(a[73] & b[310])^(a[72] & b[311])^(a[71] & b[312])^(a[70] & b[313])^(a[69] & b[314])^(a[68] & b[315])^(a[67] & b[316])^(a[66] & b[317])^(a[65] & b[318])^(a[64] & b[319])^(a[63] & b[320])^(a[62] & b[321])^(a[61] & b[322])^(a[60] & b[323])^(a[59] & b[324])^(a[58] & b[325])^(a[57] & b[326])^(a[56] & b[327])^(a[55] & b[328])^(a[54] & b[329])^(a[53] & b[330])^(a[52] & b[331])^(a[51] & b[332])^(a[50] & b[333])^(a[49] & b[334])^(a[48] & b[335])^(a[47] & b[336])^(a[46] & b[337])^(a[45] & b[338])^(a[44] & b[339])^(a[43] & b[340])^(a[42] & b[341])^(a[41] & b[342])^(a[40] & b[343])^(a[39] & b[344])^(a[38] & b[345])^(a[37] & b[346])^(a[36] & b[347])^(a[35] & b[348])^(a[34] & b[349])^(a[33] & b[350])^(a[32] & b[351])^(a[31] & b[352])^(a[30] & b[353])^(a[29] & b[354])^(a[28] & b[355])^(a[27] & b[356])^(a[26] & b[357])^(a[25] & b[358])^(a[24] & b[359])^(a[23] & b[360])^(a[22] & b[361])^(a[21] & b[362])^(a[20] & b[363])^(a[19] & b[364])^(a[18] & b[365])^(a[17] & b[366])^(a[16] & b[367])^(a[15] & b[368])^(a[14] & b[369])^(a[13] & b[370])^(a[12] & b[371])^(a[11] & b[372])^(a[10] & b[373])^(a[9] & b[374])^(a[8] & b[375])^(a[7] & b[376])^(a[6] & b[377])^(a[5] & b[378])^(a[4] & b[379])^(a[3] & b[380])^(a[2] & b[381])^(a[1] & b[382])^(a[0] & b[383]);
assign y[384] = (a[384] & b[0])^(a[383] & b[1])^(a[382] & b[2])^(a[381] & b[3])^(a[380] & b[4])^(a[379] & b[5])^(a[378] & b[6])^(a[377] & b[7])^(a[376] & b[8])^(a[375] & b[9])^(a[374] & b[10])^(a[373] & b[11])^(a[372] & b[12])^(a[371] & b[13])^(a[370] & b[14])^(a[369] & b[15])^(a[368] & b[16])^(a[367] & b[17])^(a[366] & b[18])^(a[365] & b[19])^(a[364] & b[20])^(a[363] & b[21])^(a[362] & b[22])^(a[361] & b[23])^(a[360] & b[24])^(a[359] & b[25])^(a[358] & b[26])^(a[357] & b[27])^(a[356] & b[28])^(a[355] & b[29])^(a[354] & b[30])^(a[353] & b[31])^(a[352] & b[32])^(a[351] & b[33])^(a[350] & b[34])^(a[349] & b[35])^(a[348] & b[36])^(a[347] & b[37])^(a[346] & b[38])^(a[345] & b[39])^(a[344] & b[40])^(a[343] & b[41])^(a[342] & b[42])^(a[341] & b[43])^(a[340] & b[44])^(a[339] & b[45])^(a[338] & b[46])^(a[337] & b[47])^(a[336] & b[48])^(a[335] & b[49])^(a[334] & b[50])^(a[333] & b[51])^(a[332] & b[52])^(a[331] & b[53])^(a[330] & b[54])^(a[329] & b[55])^(a[328] & b[56])^(a[327] & b[57])^(a[326] & b[58])^(a[325] & b[59])^(a[324] & b[60])^(a[323] & b[61])^(a[322] & b[62])^(a[321] & b[63])^(a[320] & b[64])^(a[319] & b[65])^(a[318] & b[66])^(a[317] & b[67])^(a[316] & b[68])^(a[315] & b[69])^(a[314] & b[70])^(a[313] & b[71])^(a[312] & b[72])^(a[311] & b[73])^(a[310] & b[74])^(a[309] & b[75])^(a[308] & b[76])^(a[307] & b[77])^(a[306] & b[78])^(a[305] & b[79])^(a[304] & b[80])^(a[303] & b[81])^(a[302] & b[82])^(a[301] & b[83])^(a[300] & b[84])^(a[299] & b[85])^(a[298] & b[86])^(a[297] & b[87])^(a[296] & b[88])^(a[295] & b[89])^(a[294] & b[90])^(a[293] & b[91])^(a[292] & b[92])^(a[291] & b[93])^(a[290] & b[94])^(a[289] & b[95])^(a[288] & b[96])^(a[287] & b[97])^(a[286] & b[98])^(a[285] & b[99])^(a[284] & b[100])^(a[283] & b[101])^(a[282] & b[102])^(a[281] & b[103])^(a[280] & b[104])^(a[279] & b[105])^(a[278] & b[106])^(a[277] & b[107])^(a[276] & b[108])^(a[275] & b[109])^(a[274] & b[110])^(a[273] & b[111])^(a[272] & b[112])^(a[271] & b[113])^(a[270] & b[114])^(a[269] & b[115])^(a[268] & b[116])^(a[267] & b[117])^(a[266] & b[118])^(a[265] & b[119])^(a[264] & b[120])^(a[263] & b[121])^(a[262] & b[122])^(a[261] & b[123])^(a[260] & b[124])^(a[259] & b[125])^(a[258] & b[126])^(a[257] & b[127])^(a[256] & b[128])^(a[255] & b[129])^(a[254] & b[130])^(a[253] & b[131])^(a[252] & b[132])^(a[251] & b[133])^(a[250] & b[134])^(a[249] & b[135])^(a[248] & b[136])^(a[247] & b[137])^(a[246] & b[138])^(a[245] & b[139])^(a[244] & b[140])^(a[243] & b[141])^(a[242] & b[142])^(a[241] & b[143])^(a[240] & b[144])^(a[239] & b[145])^(a[238] & b[146])^(a[237] & b[147])^(a[236] & b[148])^(a[235] & b[149])^(a[234] & b[150])^(a[233] & b[151])^(a[232] & b[152])^(a[231] & b[153])^(a[230] & b[154])^(a[229] & b[155])^(a[228] & b[156])^(a[227] & b[157])^(a[226] & b[158])^(a[225] & b[159])^(a[224] & b[160])^(a[223] & b[161])^(a[222] & b[162])^(a[221] & b[163])^(a[220] & b[164])^(a[219] & b[165])^(a[218] & b[166])^(a[217] & b[167])^(a[216] & b[168])^(a[215] & b[169])^(a[214] & b[170])^(a[213] & b[171])^(a[212] & b[172])^(a[211] & b[173])^(a[210] & b[174])^(a[209] & b[175])^(a[208] & b[176])^(a[207] & b[177])^(a[206] & b[178])^(a[205] & b[179])^(a[204] & b[180])^(a[203] & b[181])^(a[202] & b[182])^(a[201] & b[183])^(a[200] & b[184])^(a[199] & b[185])^(a[198] & b[186])^(a[197] & b[187])^(a[196] & b[188])^(a[195] & b[189])^(a[194] & b[190])^(a[193] & b[191])^(a[192] & b[192])^(a[191] & b[193])^(a[190] & b[194])^(a[189] & b[195])^(a[188] & b[196])^(a[187] & b[197])^(a[186] & b[198])^(a[185] & b[199])^(a[184] & b[200])^(a[183] & b[201])^(a[182] & b[202])^(a[181] & b[203])^(a[180] & b[204])^(a[179] & b[205])^(a[178] & b[206])^(a[177] & b[207])^(a[176] & b[208])^(a[175] & b[209])^(a[174] & b[210])^(a[173] & b[211])^(a[172] & b[212])^(a[171] & b[213])^(a[170] & b[214])^(a[169] & b[215])^(a[168] & b[216])^(a[167] & b[217])^(a[166] & b[218])^(a[165] & b[219])^(a[164] & b[220])^(a[163] & b[221])^(a[162] & b[222])^(a[161] & b[223])^(a[160] & b[224])^(a[159] & b[225])^(a[158] & b[226])^(a[157] & b[227])^(a[156] & b[228])^(a[155] & b[229])^(a[154] & b[230])^(a[153] & b[231])^(a[152] & b[232])^(a[151] & b[233])^(a[150] & b[234])^(a[149] & b[235])^(a[148] & b[236])^(a[147] & b[237])^(a[146] & b[238])^(a[145] & b[239])^(a[144] & b[240])^(a[143] & b[241])^(a[142] & b[242])^(a[141] & b[243])^(a[140] & b[244])^(a[139] & b[245])^(a[138] & b[246])^(a[137] & b[247])^(a[136] & b[248])^(a[135] & b[249])^(a[134] & b[250])^(a[133] & b[251])^(a[132] & b[252])^(a[131] & b[253])^(a[130] & b[254])^(a[129] & b[255])^(a[128] & b[256])^(a[127] & b[257])^(a[126] & b[258])^(a[125] & b[259])^(a[124] & b[260])^(a[123] & b[261])^(a[122] & b[262])^(a[121] & b[263])^(a[120] & b[264])^(a[119] & b[265])^(a[118] & b[266])^(a[117] & b[267])^(a[116] & b[268])^(a[115] & b[269])^(a[114] & b[270])^(a[113] & b[271])^(a[112] & b[272])^(a[111] & b[273])^(a[110] & b[274])^(a[109] & b[275])^(a[108] & b[276])^(a[107] & b[277])^(a[106] & b[278])^(a[105] & b[279])^(a[104] & b[280])^(a[103] & b[281])^(a[102] & b[282])^(a[101] & b[283])^(a[100] & b[284])^(a[99] & b[285])^(a[98] & b[286])^(a[97] & b[287])^(a[96] & b[288])^(a[95] & b[289])^(a[94] & b[290])^(a[93] & b[291])^(a[92] & b[292])^(a[91] & b[293])^(a[90] & b[294])^(a[89] & b[295])^(a[88] & b[296])^(a[87] & b[297])^(a[86] & b[298])^(a[85] & b[299])^(a[84] & b[300])^(a[83] & b[301])^(a[82] & b[302])^(a[81] & b[303])^(a[80] & b[304])^(a[79] & b[305])^(a[78] & b[306])^(a[77] & b[307])^(a[76] & b[308])^(a[75] & b[309])^(a[74] & b[310])^(a[73] & b[311])^(a[72] & b[312])^(a[71] & b[313])^(a[70] & b[314])^(a[69] & b[315])^(a[68] & b[316])^(a[67] & b[317])^(a[66] & b[318])^(a[65] & b[319])^(a[64] & b[320])^(a[63] & b[321])^(a[62] & b[322])^(a[61] & b[323])^(a[60] & b[324])^(a[59] & b[325])^(a[58] & b[326])^(a[57] & b[327])^(a[56] & b[328])^(a[55] & b[329])^(a[54] & b[330])^(a[53] & b[331])^(a[52] & b[332])^(a[51] & b[333])^(a[50] & b[334])^(a[49] & b[335])^(a[48] & b[336])^(a[47] & b[337])^(a[46] & b[338])^(a[45] & b[339])^(a[44] & b[340])^(a[43] & b[341])^(a[42] & b[342])^(a[41] & b[343])^(a[40] & b[344])^(a[39] & b[345])^(a[38] & b[346])^(a[37] & b[347])^(a[36] & b[348])^(a[35] & b[349])^(a[34] & b[350])^(a[33] & b[351])^(a[32] & b[352])^(a[31] & b[353])^(a[30] & b[354])^(a[29] & b[355])^(a[28] & b[356])^(a[27] & b[357])^(a[26] & b[358])^(a[25] & b[359])^(a[24] & b[360])^(a[23] & b[361])^(a[22] & b[362])^(a[21] & b[363])^(a[20] & b[364])^(a[19] & b[365])^(a[18] & b[366])^(a[17] & b[367])^(a[16] & b[368])^(a[15] & b[369])^(a[14] & b[370])^(a[13] & b[371])^(a[12] & b[372])^(a[11] & b[373])^(a[10] & b[374])^(a[9] & b[375])^(a[8] & b[376])^(a[7] & b[377])^(a[6] & b[378])^(a[5] & b[379])^(a[4] & b[380])^(a[3] & b[381])^(a[2] & b[382])^(a[1] & b[383])^(a[0] & b[384]);
assign y[385] = (a[385] & b[0])^(a[384] & b[1])^(a[383] & b[2])^(a[382] & b[3])^(a[381] & b[4])^(a[380] & b[5])^(a[379] & b[6])^(a[378] & b[7])^(a[377] & b[8])^(a[376] & b[9])^(a[375] & b[10])^(a[374] & b[11])^(a[373] & b[12])^(a[372] & b[13])^(a[371] & b[14])^(a[370] & b[15])^(a[369] & b[16])^(a[368] & b[17])^(a[367] & b[18])^(a[366] & b[19])^(a[365] & b[20])^(a[364] & b[21])^(a[363] & b[22])^(a[362] & b[23])^(a[361] & b[24])^(a[360] & b[25])^(a[359] & b[26])^(a[358] & b[27])^(a[357] & b[28])^(a[356] & b[29])^(a[355] & b[30])^(a[354] & b[31])^(a[353] & b[32])^(a[352] & b[33])^(a[351] & b[34])^(a[350] & b[35])^(a[349] & b[36])^(a[348] & b[37])^(a[347] & b[38])^(a[346] & b[39])^(a[345] & b[40])^(a[344] & b[41])^(a[343] & b[42])^(a[342] & b[43])^(a[341] & b[44])^(a[340] & b[45])^(a[339] & b[46])^(a[338] & b[47])^(a[337] & b[48])^(a[336] & b[49])^(a[335] & b[50])^(a[334] & b[51])^(a[333] & b[52])^(a[332] & b[53])^(a[331] & b[54])^(a[330] & b[55])^(a[329] & b[56])^(a[328] & b[57])^(a[327] & b[58])^(a[326] & b[59])^(a[325] & b[60])^(a[324] & b[61])^(a[323] & b[62])^(a[322] & b[63])^(a[321] & b[64])^(a[320] & b[65])^(a[319] & b[66])^(a[318] & b[67])^(a[317] & b[68])^(a[316] & b[69])^(a[315] & b[70])^(a[314] & b[71])^(a[313] & b[72])^(a[312] & b[73])^(a[311] & b[74])^(a[310] & b[75])^(a[309] & b[76])^(a[308] & b[77])^(a[307] & b[78])^(a[306] & b[79])^(a[305] & b[80])^(a[304] & b[81])^(a[303] & b[82])^(a[302] & b[83])^(a[301] & b[84])^(a[300] & b[85])^(a[299] & b[86])^(a[298] & b[87])^(a[297] & b[88])^(a[296] & b[89])^(a[295] & b[90])^(a[294] & b[91])^(a[293] & b[92])^(a[292] & b[93])^(a[291] & b[94])^(a[290] & b[95])^(a[289] & b[96])^(a[288] & b[97])^(a[287] & b[98])^(a[286] & b[99])^(a[285] & b[100])^(a[284] & b[101])^(a[283] & b[102])^(a[282] & b[103])^(a[281] & b[104])^(a[280] & b[105])^(a[279] & b[106])^(a[278] & b[107])^(a[277] & b[108])^(a[276] & b[109])^(a[275] & b[110])^(a[274] & b[111])^(a[273] & b[112])^(a[272] & b[113])^(a[271] & b[114])^(a[270] & b[115])^(a[269] & b[116])^(a[268] & b[117])^(a[267] & b[118])^(a[266] & b[119])^(a[265] & b[120])^(a[264] & b[121])^(a[263] & b[122])^(a[262] & b[123])^(a[261] & b[124])^(a[260] & b[125])^(a[259] & b[126])^(a[258] & b[127])^(a[257] & b[128])^(a[256] & b[129])^(a[255] & b[130])^(a[254] & b[131])^(a[253] & b[132])^(a[252] & b[133])^(a[251] & b[134])^(a[250] & b[135])^(a[249] & b[136])^(a[248] & b[137])^(a[247] & b[138])^(a[246] & b[139])^(a[245] & b[140])^(a[244] & b[141])^(a[243] & b[142])^(a[242] & b[143])^(a[241] & b[144])^(a[240] & b[145])^(a[239] & b[146])^(a[238] & b[147])^(a[237] & b[148])^(a[236] & b[149])^(a[235] & b[150])^(a[234] & b[151])^(a[233] & b[152])^(a[232] & b[153])^(a[231] & b[154])^(a[230] & b[155])^(a[229] & b[156])^(a[228] & b[157])^(a[227] & b[158])^(a[226] & b[159])^(a[225] & b[160])^(a[224] & b[161])^(a[223] & b[162])^(a[222] & b[163])^(a[221] & b[164])^(a[220] & b[165])^(a[219] & b[166])^(a[218] & b[167])^(a[217] & b[168])^(a[216] & b[169])^(a[215] & b[170])^(a[214] & b[171])^(a[213] & b[172])^(a[212] & b[173])^(a[211] & b[174])^(a[210] & b[175])^(a[209] & b[176])^(a[208] & b[177])^(a[207] & b[178])^(a[206] & b[179])^(a[205] & b[180])^(a[204] & b[181])^(a[203] & b[182])^(a[202] & b[183])^(a[201] & b[184])^(a[200] & b[185])^(a[199] & b[186])^(a[198] & b[187])^(a[197] & b[188])^(a[196] & b[189])^(a[195] & b[190])^(a[194] & b[191])^(a[193] & b[192])^(a[192] & b[193])^(a[191] & b[194])^(a[190] & b[195])^(a[189] & b[196])^(a[188] & b[197])^(a[187] & b[198])^(a[186] & b[199])^(a[185] & b[200])^(a[184] & b[201])^(a[183] & b[202])^(a[182] & b[203])^(a[181] & b[204])^(a[180] & b[205])^(a[179] & b[206])^(a[178] & b[207])^(a[177] & b[208])^(a[176] & b[209])^(a[175] & b[210])^(a[174] & b[211])^(a[173] & b[212])^(a[172] & b[213])^(a[171] & b[214])^(a[170] & b[215])^(a[169] & b[216])^(a[168] & b[217])^(a[167] & b[218])^(a[166] & b[219])^(a[165] & b[220])^(a[164] & b[221])^(a[163] & b[222])^(a[162] & b[223])^(a[161] & b[224])^(a[160] & b[225])^(a[159] & b[226])^(a[158] & b[227])^(a[157] & b[228])^(a[156] & b[229])^(a[155] & b[230])^(a[154] & b[231])^(a[153] & b[232])^(a[152] & b[233])^(a[151] & b[234])^(a[150] & b[235])^(a[149] & b[236])^(a[148] & b[237])^(a[147] & b[238])^(a[146] & b[239])^(a[145] & b[240])^(a[144] & b[241])^(a[143] & b[242])^(a[142] & b[243])^(a[141] & b[244])^(a[140] & b[245])^(a[139] & b[246])^(a[138] & b[247])^(a[137] & b[248])^(a[136] & b[249])^(a[135] & b[250])^(a[134] & b[251])^(a[133] & b[252])^(a[132] & b[253])^(a[131] & b[254])^(a[130] & b[255])^(a[129] & b[256])^(a[128] & b[257])^(a[127] & b[258])^(a[126] & b[259])^(a[125] & b[260])^(a[124] & b[261])^(a[123] & b[262])^(a[122] & b[263])^(a[121] & b[264])^(a[120] & b[265])^(a[119] & b[266])^(a[118] & b[267])^(a[117] & b[268])^(a[116] & b[269])^(a[115] & b[270])^(a[114] & b[271])^(a[113] & b[272])^(a[112] & b[273])^(a[111] & b[274])^(a[110] & b[275])^(a[109] & b[276])^(a[108] & b[277])^(a[107] & b[278])^(a[106] & b[279])^(a[105] & b[280])^(a[104] & b[281])^(a[103] & b[282])^(a[102] & b[283])^(a[101] & b[284])^(a[100] & b[285])^(a[99] & b[286])^(a[98] & b[287])^(a[97] & b[288])^(a[96] & b[289])^(a[95] & b[290])^(a[94] & b[291])^(a[93] & b[292])^(a[92] & b[293])^(a[91] & b[294])^(a[90] & b[295])^(a[89] & b[296])^(a[88] & b[297])^(a[87] & b[298])^(a[86] & b[299])^(a[85] & b[300])^(a[84] & b[301])^(a[83] & b[302])^(a[82] & b[303])^(a[81] & b[304])^(a[80] & b[305])^(a[79] & b[306])^(a[78] & b[307])^(a[77] & b[308])^(a[76] & b[309])^(a[75] & b[310])^(a[74] & b[311])^(a[73] & b[312])^(a[72] & b[313])^(a[71] & b[314])^(a[70] & b[315])^(a[69] & b[316])^(a[68] & b[317])^(a[67] & b[318])^(a[66] & b[319])^(a[65] & b[320])^(a[64] & b[321])^(a[63] & b[322])^(a[62] & b[323])^(a[61] & b[324])^(a[60] & b[325])^(a[59] & b[326])^(a[58] & b[327])^(a[57] & b[328])^(a[56] & b[329])^(a[55] & b[330])^(a[54] & b[331])^(a[53] & b[332])^(a[52] & b[333])^(a[51] & b[334])^(a[50] & b[335])^(a[49] & b[336])^(a[48] & b[337])^(a[47] & b[338])^(a[46] & b[339])^(a[45] & b[340])^(a[44] & b[341])^(a[43] & b[342])^(a[42] & b[343])^(a[41] & b[344])^(a[40] & b[345])^(a[39] & b[346])^(a[38] & b[347])^(a[37] & b[348])^(a[36] & b[349])^(a[35] & b[350])^(a[34] & b[351])^(a[33] & b[352])^(a[32] & b[353])^(a[31] & b[354])^(a[30] & b[355])^(a[29] & b[356])^(a[28] & b[357])^(a[27] & b[358])^(a[26] & b[359])^(a[25] & b[360])^(a[24] & b[361])^(a[23] & b[362])^(a[22] & b[363])^(a[21] & b[364])^(a[20] & b[365])^(a[19] & b[366])^(a[18] & b[367])^(a[17] & b[368])^(a[16] & b[369])^(a[15] & b[370])^(a[14] & b[371])^(a[13] & b[372])^(a[12] & b[373])^(a[11] & b[374])^(a[10] & b[375])^(a[9] & b[376])^(a[8] & b[377])^(a[7] & b[378])^(a[6] & b[379])^(a[5] & b[380])^(a[4] & b[381])^(a[3] & b[382])^(a[2] & b[383])^(a[1] & b[384])^(a[0] & b[385]);
assign y[386] = (a[386] & b[0])^(a[385] & b[1])^(a[384] & b[2])^(a[383] & b[3])^(a[382] & b[4])^(a[381] & b[5])^(a[380] & b[6])^(a[379] & b[7])^(a[378] & b[8])^(a[377] & b[9])^(a[376] & b[10])^(a[375] & b[11])^(a[374] & b[12])^(a[373] & b[13])^(a[372] & b[14])^(a[371] & b[15])^(a[370] & b[16])^(a[369] & b[17])^(a[368] & b[18])^(a[367] & b[19])^(a[366] & b[20])^(a[365] & b[21])^(a[364] & b[22])^(a[363] & b[23])^(a[362] & b[24])^(a[361] & b[25])^(a[360] & b[26])^(a[359] & b[27])^(a[358] & b[28])^(a[357] & b[29])^(a[356] & b[30])^(a[355] & b[31])^(a[354] & b[32])^(a[353] & b[33])^(a[352] & b[34])^(a[351] & b[35])^(a[350] & b[36])^(a[349] & b[37])^(a[348] & b[38])^(a[347] & b[39])^(a[346] & b[40])^(a[345] & b[41])^(a[344] & b[42])^(a[343] & b[43])^(a[342] & b[44])^(a[341] & b[45])^(a[340] & b[46])^(a[339] & b[47])^(a[338] & b[48])^(a[337] & b[49])^(a[336] & b[50])^(a[335] & b[51])^(a[334] & b[52])^(a[333] & b[53])^(a[332] & b[54])^(a[331] & b[55])^(a[330] & b[56])^(a[329] & b[57])^(a[328] & b[58])^(a[327] & b[59])^(a[326] & b[60])^(a[325] & b[61])^(a[324] & b[62])^(a[323] & b[63])^(a[322] & b[64])^(a[321] & b[65])^(a[320] & b[66])^(a[319] & b[67])^(a[318] & b[68])^(a[317] & b[69])^(a[316] & b[70])^(a[315] & b[71])^(a[314] & b[72])^(a[313] & b[73])^(a[312] & b[74])^(a[311] & b[75])^(a[310] & b[76])^(a[309] & b[77])^(a[308] & b[78])^(a[307] & b[79])^(a[306] & b[80])^(a[305] & b[81])^(a[304] & b[82])^(a[303] & b[83])^(a[302] & b[84])^(a[301] & b[85])^(a[300] & b[86])^(a[299] & b[87])^(a[298] & b[88])^(a[297] & b[89])^(a[296] & b[90])^(a[295] & b[91])^(a[294] & b[92])^(a[293] & b[93])^(a[292] & b[94])^(a[291] & b[95])^(a[290] & b[96])^(a[289] & b[97])^(a[288] & b[98])^(a[287] & b[99])^(a[286] & b[100])^(a[285] & b[101])^(a[284] & b[102])^(a[283] & b[103])^(a[282] & b[104])^(a[281] & b[105])^(a[280] & b[106])^(a[279] & b[107])^(a[278] & b[108])^(a[277] & b[109])^(a[276] & b[110])^(a[275] & b[111])^(a[274] & b[112])^(a[273] & b[113])^(a[272] & b[114])^(a[271] & b[115])^(a[270] & b[116])^(a[269] & b[117])^(a[268] & b[118])^(a[267] & b[119])^(a[266] & b[120])^(a[265] & b[121])^(a[264] & b[122])^(a[263] & b[123])^(a[262] & b[124])^(a[261] & b[125])^(a[260] & b[126])^(a[259] & b[127])^(a[258] & b[128])^(a[257] & b[129])^(a[256] & b[130])^(a[255] & b[131])^(a[254] & b[132])^(a[253] & b[133])^(a[252] & b[134])^(a[251] & b[135])^(a[250] & b[136])^(a[249] & b[137])^(a[248] & b[138])^(a[247] & b[139])^(a[246] & b[140])^(a[245] & b[141])^(a[244] & b[142])^(a[243] & b[143])^(a[242] & b[144])^(a[241] & b[145])^(a[240] & b[146])^(a[239] & b[147])^(a[238] & b[148])^(a[237] & b[149])^(a[236] & b[150])^(a[235] & b[151])^(a[234] & b[152])^(a[233] & b[153])^(a[232] & b[154])^(a[231] & b[155])^(a[230] & b[156])^(a[229] & b[157])^(a[228] & b[158])^(a[227] & b[159])^(a[226] & b[160])^(a[225] & b[161])^(a[224] & b[162])^(a[223] & b[163])^(a[222] & b[164])^(a[221] & b[165])^(a[220] & b[166])^(a[219] & b[167])^(a[218] & b[168])^(a[217] & b[169])^(a[216] & b[170])^(a[215] & b[171])^(a[214] & b[172])^(a[213] & b[173])^(a[212] & b[174])^(a[211] & b[175])^(a[210] & b[176])^(a[209] & b[177])^(a[208] & b[178])^(a[207] & b[179])^(a[206] & b[180])^(a[205] & b[181])^(a[204] & b[182])^(a[203] & b[183])^(a[202] & b[184])^(a[201] & b[185])^(a[200] & b[186])^(a[199] & b[187])^(a[198] & b[188])^(a[197] & b[189])^(a[196] & b[190])^(a[195] & b[191])^(a[194] & b[192])^(a[193] & b[193])^(a[192] & b[194])^(a[191] & b[195])^(a[190] & b[196])^(a[189] & b[197])^(a[188] & b[198])^(a[187] & b[199])^(a[186] & b[200])^(a[185] & b[201])^(a[184] & b[202])^(a[183] & b[203])^(a[182] & b[204])^(a[181] & b[205])^(a[180] & b[206])^(a[179] & b[207])^(a[178] & b[208])^(a[177] & b[209])^(a[176] & b[210])^(a[175] & b[211])^(a[174] & b[212])^(a[173] & b[213])^(a[172] & b[214])^(a[171] & b[215])^(a[170] & b[216])^(a[169] & b[217])^(a[168] & b[218])^(a[167] & b[219])^(a[166] & b[220])^(a[165] & b[221])^(a[164] & b[222])^(a[163] & b[223])^(a[162] & b[224])^(a[161] & b[225])^(a[160] & b[226])^(a[159] & b[227])^(a[158] & b[228])^(a[157] & b[229])^(a[156] & b[230])^(a[155] & b[231])^(a[154] & b[232])^(a[153] & b[233])^(a[152] & b[234])^(a[151] & b[235])^(a[150] & b[236])^(a[149] & b[237])^(a[148] & b[238])^(a[147] & b[239])^(a[146] & b[240])^(a[145] & b[241])^(a[144] & b[242])^(a[143] & b[243])^(a[142] & b[244])^(a[141] & b[245])^(a[140] & b[246])^(a[139] & b[247])^(a[138] & b[248])^(a[137] & b[249])^(a[136] & b[250])^(a[135] & b[251])^(a[134] & b[252])^(a[133] & b[253])^(a[132] & b[254])^(a[131] & b[255])^(a[130] & b[256])^(a[129] & b[257])^(a[128] & b[258])^(a[127] & b[259])^(a[126] & b[260])^(a[125] & b[261])^(a[124] & b[262])^(a[123] & b[263])^(a[122] & b[264])^(a[121] & b[265])^(a[120] & b[266])^(a[119] & b[267])^(a[118] & b[268])^(a[117] & b[269])^(a[116] & b[270])^(a[115] & b[271])^(a[114] & b[272])^(a[113] & b[273])^(a[112] & b[274])^(a[111] & b[275])^(a[110] & b[276])^(a[109] & b[277])^(a[108] & b[278])^(a[107] & b[279])^(a[106] & b[280])^(a[105] & b[281])^(a[104] & b[282])^(a[103] & b[283])^(a[102] & b[284])^(a[101] & b[285])^(a[100] & b[286])^(a[99] & b[287])^(a[98] & b[288])^(a[97] & b[289])^(a[96] & b[290])^(a[95] & b[291])^(a[94] & b[292])^(a[93] & b[293])^(a[92] & b[294])^(a[91] & b[295])^(a[90] & b[296])^(a[89] & b[297])^(a[88] & b[298])^(a[87] & b[299])^(a[86] & b[300])^(a[85] & b[301])^(a[84] & b[302])^(a[83] & b[303])^(a[82] & b[304])^(a[81] & b[305])^(a[80] & b[306])^(a[79] & b[307])^(a[78] & b[308])^(a[77] & b[309])^(a[76] & b[310])^(a[75] & b[311])^(a[74] & b[312])^(a[73] & b[313])^(a[72] & b[314])^(a[71] & b[315])^(a[70] & b[316])^(a[69] & b[317])^(a[68] & b[318])^(a[67] & b[319])^(a[66] & b[320])^(a[65] & b[321])^(a[64] & b[322])^(a[63] & b[323])^(a[62] & b[324])^(a[61] & b[325])^(a[60] & b[326])^(a[59] & b[327])^(a[58] & b[328])^(a[57] & b[329])^(a[56] & b[330])^(a[55] & b[331])^(a[54] & b[332])^(a[53] & b[333])^(a[52] & b[334])^(a[51] & b[335])^(a[50] & b[336])^(a[49] & b[337])^(a[48] & b[338])^(a[47] & b[339])^(a[46] & b[340])^(a[45] & b[341])^(a[44] & b[342])^(a[43] & b[343])^(a[42] & b[344])^(a[41] & b[345])^(a[40] & b[346])^(a[39] & b[347])^(a[38] & b[348])^(a[37] & b[349])^(a[36] & b[350])^(a[35] & b[351])^(a[34] & b[352])^(a[33] & b[353])^(a[32] & b[354])^(a[31] & b[355])^(a[30] & b[356])^(a[29] & b[357])^(a[28] & b[358])^(a[27] & b[359])^(a[26] & b[360])^(a[25] & b[361])^(a[24] & b[362])^(a[23] & b[363])^(a[22] & b[364])^(a[21] & b[365])^(a[20] & b[366])^(a[19] & b[367])^(a[18] & b[368])^(a[17] & b[369])^(a[16] & b[370])^(a[15] & b[371])^(a[14] & b[372])^(a[13] & b[373])^(a[12] & b[374])^(a[11] & b[375])^(a[10] & b[376])^(a[9] & b[377])^(a[8] & b[378])^(a[7] & b[379])^(a[6] & b[380])^(a[5] & b[381])^(a[4] & b[382])^(a[3] & b[383])^(a[2] & b[384])^(a[1] & b[385])^(a[0] & b[386]);
assign y[387] = (a[387] & b[0])^(a[386] & b[1])^(a[385] & b[2])^(a[384] & b[3])^(a[383] & b[4])^(a[382] & b[5])^(a[381] & b[6])^(a[380] & b[7])^(a[379] & b[8])^(a[378] & b[9])^(a[377] & b[10])^(a[376] & b[11])^(a[375] & b[12])^(a[374] & b[13])^(a[373] & b[14])^(a[372] & b[15])^(a[371] & b[16])^(a[370] & b[17])^(a[369] & b[18])^(a[368] & b[19])^(a[367] & b[20])^(a[366] & b[21])^(a[365] & b[22])^(a[364] & b[23])^(a[363] & b[24])^(a[362] & b[25])^(a[361] & b[26])^(a[360] & b[27])^(a[359] & b[28])^(a[358] & b[29])^(a[357] & b[30])^(a[356] & b[31])^(a[355] & b[32])^(a[354] & b[33])^(a[353] & b[34])^(a[352] & b[35])^(a[351] & b[36])^(a[350] & b[37])^(a[349] & b[38])^(a[348] & b[39])^(a[347] & b[40])^(a[346] & b[41])^(a[345] & b[42])^(a[344] & b[43])^(a[343] & b[44])^(a[342] & b[45])^(a[341] & b[46])^(a[340] & b[47])^(a[339] & b[48])^(a[338] & b[49])^(a[337] & b[50])^(a[336] & b[51])^(a[335] & b[52])^(a[334] & b[53])^(a[333] & b[54])^(a[332] & b[55])^(a[331] & b[56])^(a[330] & b[57])^(a[329] & b[58])^(a[328] & b[59])^(a[327] & b[60])^(a[326] & b[61])^(a[325] & b[62])^(a[324] & b[63])^(a[323] & b[64])^(a[322] & b[65])^(a[321] & b[66])^(a[320] & b[67])^(a[319] & b[68])^(a[318] & b[69])^(a[317] & b[70])^(a[316] & b[71])^(a[315] & b[72])^(a[314] & b[73])^(a[313] & b[74])^(a[312] & b[75])^(a[311] & b[76])^(a[310] & b[77])^(a[309] & b[78])^(a[308] & b[79])^(a[307] & b[80])^(a[306] & b[81])^(a[305] & b[82])^(a[304] & b[83])^(a[303] & b[84])^(a[302] & b[85])^(a[301] & b[86])^(a[300] & b[87])^(a[299] & b[88])^(a[298] & b[89])^(a[297] & b[90])^(a[296] & b[91])^(a[295] & b[92])^(a[294] & b[93])^(a[293] & b[94])^(a[292] & b[95])^(a[291] & b[96])^(a[290] & b[97])^(a[289] & b[98])^(a[288] & b[99])^(a[287] & b[100])^(a[286] & b[101])^(a[285] & b[102])^(a[284] & b[103])^(a[283] & b[104])^(a[282] & b[105])^(a[281] & b[106])^(a[280] & b[107])^(a[279] & b[108])^(a[278] & b[109])^(a[277] & b[110])^(a[276] & b[111])^(a[275] & b[112])^(a[274] & b[113])^(a[273] & b[114])^(a[272] & b[115])^(a[271] & b[116])^(a[270] & b[117])^(a[269] & b[118])^(a[268] & b[119])^(a[267] & b[120])^(a[266] & b[121])^(a[265] & b[122])^(a[264] & b[123])^(a[263] & b[124])^(a[262] & b[125])^(a[261] & b[126])^(a[260] & b[127])^(a[259] & b[128])^(a[258] & b[129])^(a[257] & b[130])^(a[256] & b[131])^(a[255] & b[132])^(a[254] & b[133])^(a[253] & b[134])^(a[252] & b[135])^(a[251] & b[136])^(a[250] & b[137])^(a[249] & b[138])^(a[248] & b[139])^(a[247] & b[140])^(a[246] & b[141])^(a[245] & b[142])^(a[244] & b[143])^(a[243] & b[144])^(a[242] & b[145])^(a[241] & b[146])^(a[240] & b[147])^(a[239] & b[148])^(a[238] & b[149])^(a[237] & b[150])^(a[236] & b[151])^(a[235] & b[152])^(a[234] & b[153])^(a[233] & b[154])^(a[232] & b[155])^(a[231] & b[156])^(a[230] & b[157])^(a[229] & b[158])^(a[228] & b[159])^(a[227] & b[160])^(a[226] & b[161])^(a[225] & b[162])^(a[224] & b[163])^(a[223] & b[164])^(a[222] & b[165])^(a[221] & b[166])^(a[220] & b[167])^(a[219] & b[168])^(a[218] & b[169])^(a[217] & b[170])^(a[216] & b[171])^(a[215] & b[172])^(a[214] & b[173])^(a[213] & b[174])^(a[212] & b[175])^(a[211] & b[176])^(a[210] & b[177])^(a[209] & b[178])^(a[208] & b[179])^(a[207] & b[180])^(a[206] & b[181])^(a[205] & b[182])^(a[204] & b[183])^(a[203] & b[184])^(a[202] & b[185])^(a[201] & b[186])^(a[200] & b[187])^(a[199] & b[188])^(a[198] & b[189])^(a[197] & b[190])^(a[196] & b[191])^(a[195] & b[192])^(a[194] & b[193])^(a[193] & b[194])^(a[192] & b[195])^(a[191] & b[196])^(a[190] & b[197])^(a[189] & b[198])^(a[188] & b[199])^(a[187] & b[200])^(a[186] & b[201])^(a[185] & b[202])^(a[184] & b[203])^(a[183] & b[204])^(a[182] & b[205])^(a[181] & b[206])^(a[180] & b[207])^(a[179] & b[208])^(a[178] & b[209])^(a[177] & b[210])^(a[176] & b[211])^(a[175] & b[212])^(a[174] & b[213])^(a[173] & b[214])^(a[172] & b[215])^(a[171] & b[216])^(a[170] & b[217])^(a[169] & b[218])^(a[168] & b[219])^(a[167] & b[220])^(a[166] & b[221])^(a[165] & b[222])^(a[164] & b[223])^(a[163] & b[224])^(a[162] & b[225])^(a[161] & b[226])^(a[160] & b[227])^(a[159] & b[228])^(a[158] & b[229])^(a[157] & b[230])^(a[156] & b[231])^(a[155] & b[232])^(a[154] & b[233])^(a[153] & b[234])^(a[152] & b[235])^(a[151] & b[236])^(a[150] & b[237])^(a[149] & b[238])^(a[148] & b[239])^(a[147] & b[240])^(a[146] & b[241])^(a[145] & b[242])^(a[144] & b[243])^(a[143] & b[244])^(a[142] & b[245])^(a[141] & b[246])^(a[140] & b[247])^(a[139] & b[248])^(a[138] & b[249])^(a[137] & b[250])^(a[136] & b[251])^(a[135] & b[252])^(a[134] & b[253])^(a[133] & b[254])^(a[132] & b[255])^(a[131] & b[256])^(a[130] & b[257])^(a[129] & b[258])^(a[128] & b[259])^(a[127] & b[260])^(a[126] & b[261])^(a[125] & b[262])^(a[124] & b[263])^(a[123] & b[264])^(a[122] & b[265])^(a[121] & b[266])^(a[120] & b[267])^(a[119] & b[268])^(a[118] & b[269])^(a[117] & b[270])^(a[116] & b[271])^(a[115] & b[272])^(a[114] & b[273])^(a[113] & b[274])^(a[112] & b[275])^(a[111] & b[276])^(a[110] & b[277])^(a[109] & b[278])^(a[108] & b[279])^(a[107] & b[280])^(a[106] & b[281])^(a[105] & b[282])^(a[104] & b[283])^(a[103] & b[284])^(a[102] & b[285])^(a[101] & b[286])^(a[100] & b[287])^(a[99] & b[288])^(a[98] & b[289])^(a[97] & b[290])^(a[96] & b[291])^(a[95] & b[292])^(a[94] & b[293])^(a[93] & b[294])^(a[92] & b[295])^(a[91] & b[296])^(a[90] & b[297])^(a[89] & b[298])^(a[88] & b[299])^(a[87] & b[300])^(a[86] & b[301])^(a[85] & b[302])^(a[84] & b[303])^(a[83] & b[304])^(a[82] & b[305])^(a[81] & b[306])^(a[80] & b[307])^(a[79] & b[308])^(a[78] & b[309])^(a[77] & b[310])^(a[76] & b[311])^(a[75] & b[312])^(a[74] & b[313])^(a[73] & b[314])^(a[72] & b[315])^(a[71] & b[316])^(a[70] & b[317])^(a[69] & b[318])^(a[68] & b[319])^(a[67] & b[320])^(a[66] & b[321])^(a[65] & b[322])^(a[64] & b[323])^(a[63] & b[324])^(a[62] & b[325])^(a[61] & b[326])^(a[60] & b[327])^(a[59] & b[328])^(a[58] & b[329])^(a[57] & b[330])^(a[56] & b[331])^(a[55] & b[332])^(a[54] & b[333])^(a[53] & b[334])^(a[52] & b[335])^(a[51] & b[336])^(a[50] & b[337])^(a[49] & b[338])^(a[48] & b[339])^(a[47] & b[340])^(a[46] & b[341])^(a[45] & b[342])^(a[44] & b[343])^(a[43] & b[344])^(a[42] & b[345])^(a[41] & b[346])^(a[40] & b[347])^(a[39] & b[348])^(a[38] & b[349])^(a[37] & b[350])^(a[36] & b[351])^(a[35] & b[352])^(a[34] & b[353])^(a[33] & b[354])^(a[32] & b[355])^(a[31] & b[356])^(a[30] & b[357])^(a[29] & b[358])^(a[28] & b[359])^(a[27] & b[360])^(a[26] & b[361])^(a[25] & b[362])^(a[24] & b[363])^(a[23] & b[364])^(a[22] & b[365])^(a[21] & b[366])^(a[20] & b[367])^(a[19] & b[368])^(a[18] & b[369])^(a[17] & b[370])^(a[16] & b[371])^(a[15] & b[372])^(a[14] & b[373])^(a[13] & b[374])^(a[12] & b[375])^(a[11] & b[376])^(a[10] & b[377])^(a[9] & b[378])^(a[8] & b[379])^(a[7] & b[380])^(a[6] & b[381])^(a[5] & b[382])^(a[4] & b[383])^(a[3] & b[384])^(a[2] & b[385])^(a[1] & b[386])^(a[0] & b[387]);
assign y[388] = (a[388] & b[0])^(a[387] & b[1])^(a[386] & b[2])^(a[385] & b[3])^(a[384] & b[4])^(a[383] & b[5])^(a[382] & b[6])^(a[381] & b[7])^(a[380] & b[8])^(a[379] & b[9])^(a[378] & b[10])^(a[377] & b[11])^(a[376] & b[12])^(a[375] & b[13])^(a[374] & b[14])^(a[373] & b[15])^(a[372] & b[16])^(a[371] & b[17])^(a[370] & b[18])^(a[369] & b[19])^(a[368] & b[20])^(a[367] & b[21])^(a[366] & b[22])^(a[365] & b[23])^(a[364] & b[24])^(a[363] & b[25])^(a[362] & b[26])^(a[361] & b[27])^(a[360] & b[28])^(a[359] & b[29])^(a[358] & b[30])^(a[357] & b[31])^(a[356] & b[32])^(a[355] & b[33])^(a[354] & b[34])^(a[353] & b[35])^(a[352] & b[36])^(a[351] & b[37])^(a[350] & b[38])^(a[349] & b[39])^(a[348] & b[40])^(a[347] & b[41])^(a[346] & b[42])^(a[345] & b[43])^(a[344] & b[44])^(a[343] & b[45])^(a[342] & b[46])^(a[341] & b[47])^(a[340] & b[48])^(a[339] & b[49])^(a[338] & b[50])^(a[337] & b[51])^(a[336] & b[52])^(a[335] & b[53])^(a[334] & b[54])^(a[333] & b[55])^(a[332] & b[56])^(a[331] & b[57])^(a[330] & b[58])^(a[329] & b[59])^(a[328] & b[60])^(a[327] & b[61])^(a[326] & b[62])^(a[325] & b[63])^(a[324] & b[64])^(a[323] & b[65])^(a[322] & b[66])^(a[321] & b[67])^(a[320] & b[68])^(a[319] & b[69])^(a[318] & b[70])^(a[317] & b[71])^(a[316] & b[72])^(a[315] & b[73])^(a[314] & b[74])^(a[313] & b[75])^(a[312] & b[76])^(a[311] & b[77])^(a[310] & b[78])^(a[309] & b[79])^(a[308] & b[80])^(a[307] & b[81])^(a[306] & b[82])^(a[305] & b[83])^(a[304] & b[84])^(a[303] & b[85])^(a[302] & b[86])^(a[301] & b[87])^(a[300] & b[88])^(a[299] & b[89])^(a[298] & b[90])^(a[297] & b[91])^(a[296] & b[92])^(a[295] & b[93])^(a[294] & b[94])^(a[293] & b[95])^(a[292] & b[96])^(a[291] & b[97])^(a[290] & b[98])^(a[289] & b[99])^(a[288] & b[100])^(a[287] & b[101])^(a[286] & b[102])^(a[285] & b[103])^(a[284] & b[104])^(a[283] & b[105])^(a[282] & b[106])^(a[281] & b[107])^(a[280] & b[108])^(a[279] & b[109])^(a[278] & b[110])^(a[277] & b[111])^(a[276] & b[112])^(a[275] & b[113])^(a[274] & b[114])^(a[273] & b[115])^(a[272] & b[116])^(a[271] & b[117])^(a[270] & b[118])^(a[269] & b[119])^(a[268] & b[120])^(a[267] & b[121])^(a[266] & b[122])^(a[265] & b[123])^(a[264] & b[124])^(a[263] & b[125])^(a[262] & b[126])^(a[261] & b[127])^(a[260] & b[128])^(a[259] & b[129])^(a[258] & b[130])^(a[257] & b[131])^(a[256] & b[132])^(a[255] & b[133])^(a[254] & b[134])^(a[253] & b[135])^(a[252] & b[136])^(a[251] & b[137])^(a[250] & b[138])^(a[249] & b[139])^(a[248] & b[140])^(a[247] & b[141])^(a[246] & b[142])^(a[245] & b[143])^(a[244] & b[144])^(a[243] & b[145])^(a[242] & b[146])^(a[241] & b[147])^(a[240] & b[148])^(a[239] & b[149])^(a[238] & b[150])^(a[237] & b[151])^(a[236] & b[152])^(a[235] & b[153])^(a[234] & b[154])^(a[233] & b[155])^(a[232] & b[156])^(a[231] & b[157])^(a[230] & b[158])^(a[229] & b[159])^(a[228] & b[160])^(a[227] & b[161])^(a[226] & b[162])^(a[225] & b[163])^(a[224] & b[164])^(a[223] & b[165])^(a[222] & b[166])^(a[221] & b[167])^(a[220] & b[168])^(a[219] & b[169])^(a[218] & b[170])^(a[217] & b[171])^(a[216] & b[172])^(a[215] & b[173])^(a[214] & b[174])^(a[213] & b[175])^(a[212] & b[176])^(a[211] & b[177])^(a[210] & b[178])^(a[209] & b[179])^(a[208] & b[180])^(a[207] & b[181])^(a[206] & b[182])^(a[205] & b[183])^(a[204] & b[184])^(a[203] & b[185])^(a[202] & b[186])^(a[201] & b[187])^(a[200] & b[188])^(a[199] & b[189])^(a[198] & b[190])^(a[197] & b[191])^(a[196] & b[192])^(a[195] & b[193])^(a[194] & b[194])^(a[193] & b[195])^(a[192] & b[196])^(a[191] & b[197])^(a[190] & b[198])^(a[189] & b[199])^(a[188] & b[200])^(a[187] & b[201])^(a[186] & b[202])^(a[185] & b[203])^(a[184] & b[204])^(a[183] & b[205])^(a[182] & b[206])^(a[181] & b[207])^(a[180] & b[208])^(a[179] & b[209])^(a[178] & b[210])^(a[177] & b[211])^(a[176] & b[212])^(a[175] & b[213])^(a[174] & b[214])^(a[173] & b[215])^(a[172] & b[216])^(a[171] & b[217])^(a[170] & b[218])^(a[169] & b[219])^(a[168] & b[220])^(a[167] & b[221])^(a[166] & b[222])^(a[165] & b[223])^(a[164] & b[224])^(a[163] & b[225])^(a[162] & b[226])^(a[161] & b[227])^(a[160] & b[228])^(a[159] & b[229])^(a[158] & b[230])^(a[157] & b[231])^(a[156] & b[232])^(a[155] & b[233])^(a[154] & b[234])^(a[153] & b[235])^(a[152] & b[236])^(a[151] & b[237])^(a[150] & b[238])^(a[149] & b[239])^(a[148] & b[240])^(a[147] & b[241])^(a[146] & b[242])^(a[145] & b[243])^(a[144] & b[244])^(a[143] & b[245])^(a[142] & b[246])^(a[141] & b[247])^(a[140] & b[248])^(a[139] & b[249])^(a[138] & b[250])^(a[137] & b[251])^(a[136] & b[252])^(a[135] & b[253])^(a[134] & b[254])^(a[133] & b[255])^(a[132] & b[256])^(a[131] & b[257])^(a[130] & b[258])^(a[129] & b[259])^(a[128] & b[260])^(a[127] & b[261])^(a[126] & b[262])^(a[125] & b[263])^(a[124] & b[264])^(a[123] & b[265])^(a[122] & b[266])^(a[121] & b[267])^(a[120] & b[268])^(a[119] & b[269])^(a[118] & b[270])^(a[117] & b[271])^(a[116] & b[272])^(a[115] & b[273])^(a[114] & b[274])^(a[113] & b[275])^(a[112] & b[276])^(a[111] & b[277])^(a[110] & b[278])^(a[109] & b[279])^(a[108] & b[280])^(a[107] & b[281])^(a[106] & b[282])^(a[105] & b[283])^(a[104] & b[284])^(a[103] & b[285])^(a[102] & b[286])^(a[101] & b[287])^(a[100] & b[288])^(a[99] & b[289])^(a[98] & b[290])^(a[97] & b[291])^(a[96] & b[292])^(a[95] & b[293])^(a[94] & b[294])^(a[93] & b[295])^(a[92] & b[296])^(a[91] & b[297])^(a[90] & b[298])^(a[89] & b[299])^(a[88] & b[300])^(a[87] & b[301])^(a[86] & b[302])^(a[85] & b[303])^(a[84] & b[304])^(a[83] & b[305])^(a[82] & b[306])^(a[81] & b[307])^(a[80] & b[308])^(a[79] & b[309])^(a[78] & b[310])^(a[77] & b[311])^(a[76] & b[312])^(a[75] & b[313])^(a[74] & b[314])^(a[73] & b[315])^(a[72] & b[316])^(a[71] & b[317])^(a[70] & b[318])^(a[69] & b[319])^(a[68] & b[320])^(a[67] & b[321])^(a[66] & b[322])^(a[65] & b[323])^(a[64] & b[324])^(a[63] & b[325])^(a[62] & b[326])^(a[61] & b[327])^(a[60] & b[328])^(a[59] & b[329])^(a[58] & b[330])^(a[57] & b[331])^(a[56] & b[332])^(a[55] & b[333])^(a[54] & b[334])^(a[53] & b[335])^(a[52] & b[336])^(a[51] & b[337])^(a[50] & b[338])^(a[49] & b[339])^(a[48] & b[340])^(a[47] & b[341])^(a[46] & b[342])^(a[45] & b[343])^(a[44] & b[344])^(a[43] & b[345])^(a[42] & b[346])^(a[41] & b[347])^(a[40] & b[348])^(a[39] & b[349])^(a[38] & b[350])^(a[37] & b[351])^(a[36] & b[352])^(a[35] & b[353])^(a[34] & b[354])^(a[33] & b[355])^(a[32] & b[356])^(a[31] & b[357])^(a[30] & b[358])^(a[29] & b[359])^(a[28] & b[360])^(a[27] & b[361])^(a[26] & b[362])^(a[25] & b[363])^(a[24] & b[364])^(a[23] & b[365])^(a[22] & b[366])^(a[21] & b[367])^(a[20] & b[368])^(a[19] & b[369])^(a[18] & b[370])^(a[17] & b[371])^(a[16] & b[372])^(a[15] & b[373])^(a[14] & b[374])^(a[13] & b[375])^(a[12] & b[376])^(a[11] & b[377])^(a[10] & b[378])^(a[9] & b[379])^(a[8] & b[380])^(a[7] & b[381])^(a[6] & b[382])^(a[5] & b[383])^(a[4] & b[384])^(a[3] & b[385])^(a[2] & b[386])^(a[1] & b[387])^(a[0] & b[388]);
assign y[389] = (a[389] & b[0])^(a[388] & b[1])^(a[387] & b[2])^(a[386] & b[3])^(a[385] & b[4])^(a[384] & b[5])^(a[383] & b[6])^(a[382] & b[7])^(a[381] & b[8])^(a[380] & b[9])^(a[379] & b[10])^(a[378] & b[11])^(a[377] & b[12])^(a[376] & b[13])^(a[375] & b[14])^(a[374] & b[15])^(a[373] & b[16])^(a[372] & b[17])^(a[371] & b[18])^(a[370] & b[19])^(a[369] & b[20])^(a[368] & b[21])^(a[367] & b[22])^(a[366] & b[23])^(a[365] & b[24])^(a[364] & b[25])^(a[363] & b[26])^(a[362] & b[27])^(a[361] & b[28])^(a[360] & b[29])^(a[359] & b[30])^(a[358] & b[31])^(a[357] & b[32])^(a[356] & b[33])^(a[355] & b[34])^(a[354] & b[35])^(a[353] & b[36])^(a[352] & b[37])^(a[351] & b[38])^(a[350] & b[39])^(a[349] & b[40])^(a[348] & b[41])^(a[347] & b[42])^(a[346] & b[43])^(a[345] & b[44])^(a[344] & b[45])^(a[343] & b[46])^(a[342] & b[47])^(a[341] & b[48])^(a[340] & b[49])^(a[339] & b[50])^(a[338] & b[51])^(a[337] & b[52])^(a[336] & b[53])^(a[335] & b[54])^(a[334] & b[55])^(a[333] & b[56])^(a[332] & b[57])^(a[331] & b[58])^(a[330] & b[59])^(a[329] & b[60])^(a[328] & b[61])^(a[327] & b[62])^(a[326] & b[63])^(a[325] & b[64])^(a[324] & b[65])^(a[323] & b[66])^(a[322] & b[67])^(a[321] & b[68])^(a[320] & b[69])^(a[319] & b[70])^(a[318] & b[71])^(a[317] & b[72])^(a[316] & b[73])^(a[315] & b[74])^(a[314] & b[75])^(a[313] & b[76])^(a[312] & b[77])^(a[311] & b[78])^(a[310] & b[79])^(a[309] & b[80])^(a[308] & b[81])^(a[307] & b[82])^(a[306] & b[83])^(a[305] & b[84])^(a[304] & b[85])^(a[303] & b[86])^(a[302] & b[87])^(a[301] & b[88])^(a[300] & b[89])^(a[299] & b[90])^(a[298] & b[91])^(a[297] & b[92])^(a[296] & b[93])^(a[295] & b[94])^(a[294] & b[95])^(a[293] & b[96])^(a[292] & b[97])^(a[291] & b[98])^(a[290] & b[99])^(a[289] & b[100])^(a[288] & b[101])^(a[287] & b[102])^(a[286] & b[103])^(a[285] & b[104])^(a[284] & b[105])^(a[283] & b[106])^(a[282] & b[107])^(a[281] & b[108])^(a[280] & b[109])^(a[279] & b[110])^(a[278] & b[111])^(a[277] & b[112])^(a[276] & b[113])^(a[275] & b[114])^(a[274] & b[115])^(a[273] & b[116])^(a[272] & b[117])^(a[271] & b[118])^(a[270] & b[119])^(a[269] & b[120])^(a[268] & b[121])^(a[267] & b[122])^(a[266] & b[123])^(a[265] & b[124])^(a[264] & b[125])^(a[263] & b[126])^(a[262] & b[127])^(a[261] & b[128])^(a[260] & b[129])^(a[259] & b[130])^(a[258] & b[131])^(a[257] & b[132])^(a[256] & b[133])^(a[255] & b[134])^(a[254] & b[135])^(a[253] & b[136])^(a[252] & b[137])^(a[251] & b[138])^(a[250] & b[139])^(a[249] & b[140])^(a[248] & b[141])^(a[247] & b[142])^(a[246] & b[143])^(a[245] & b[144])^(a[244] & b[145])^(a[243] & b[146])^(a[242] & b[147])^(a[241] & b[148])^(a[240] & b[149])^(a[239] & b[150])^(a[238] & b[151])^(a[237] & b[152])^(a[236] & b[153])^(a[235] & b[154])^(a[234] & b[155])^(a[233] & b[156])^(a[232] & b[157])^(a[231] & b[158])^(a[230] & b[159])^(a[229] & b[160])^(a[228] & b[161])^(a[227] & b[162])^(a[226] & b[163])^(a[225] & b[164])^(a[224] & b[165])^(a[223] & b[166])^(a[222] & b[167])^(a[221] & b[168])^(a[220] & b[169])^(a[219] & b[170])^(a[218] & b[171])^(a[217] & b[172])^(a[216] & b[173])^(a[215] & b[174])^(a[214] & b[175])^(a[213] & b[176])^(a[212] & b[177])^(a[211] & b[178])^(a[210] & b[179])^(a[209] & b[180])^(a[208] & b[181])^(a[207] & b[182])^(a[206] & b[183])^(a[205] & b[184])^(a[204] & b[185])^(a[203] & b[186])^(a[202] & b[187])^(a[201] & b[188])^(a[200] & b[189])^(a[199] & b[190])^(a[198] & b[191])^(a[197] & b[192])^(a[196] & b[193])^(a[195] & b[194])^(a[194] & b[195])^(a[193] & b[196])^(a[192] & b[197])^(a[191] & b[198])^(a[190] & b[199])^(a[189] & b[200])^(a[188] & b[201])^(a[187] & b[202])^(a[186] & b[203])^(a[185] & b[204])^(a[184] & b[205])^(a[183] & b[206])^(a[182] & b[207])^(a[181] & b[208])^(a[180] & b[209])^(a[179] & b[210])^(a[178] & b[211])^(a[177] & b[212])^(a[176] & b[213])^(a[175] & b[214])^(a[174] & b[215])^(a[173] & b[216])^(a[172] & b[217])^(a[171] & b[218])^(a[170] & b[219])^(a[169] & b[220])^(a[168] & b[221])^(a[167] & b[222])^(a[166] & b[223])^(a[165] & b[224])^(a[164] & b[225])^(a[163] & b[226])^(a[162] & b[227])^(a[161] & b[228])^(a[160] & b[229])^(a[159] & b[230])^(a[158] & b[231])^(a[157] & b[232])^(a[156] & b[233])^(a[155] & b[234])^(a[154] & b[235])^(a[153] & b[236])^(a[152] & b[237])^(a[151] & b[238])^(a[150] & b[239])^(a[149] & b[240])^(a[148] & b[241])^(a[147] & b[242])^(a[146] & b[243])^(a[145] & b[244])^(a[144] & b[245])^(a[143] & b[246])^(a[142] & b[247])^(a[141] & b[248])^(a[140] & b[249])^(a[139] & b[250])^(a[138] & b[251])^(a[137] & b[252])^(a[136] & b[253])^(a[135] & b[254])^(a[134] & b[255])^(a[133] & b[256])^(a[132] & b[257])^(a[131] & b[258])^(a[130] & b[259])^(a[129] & b[260])^(a[128] & b[261])^(a[127] & b[262])^(a[126] & b[263])^(a[125] & b[264])^(a[124] & b[265])^(a[123] & b[266])^(a[122] & b[267])^(a[121] & b[268])^(a[120] & b[269])^(a[119] & b[270])^(a[118] & b[271])^(a[117] & b[272])^(a[116] & b[273])^(a[115] & b[274])^(a[114] & b[275])^(a[113] & b[276])^(a[112] & b[277])^(a[111] & b[278])^(a[110] & b[279])^(a[109] & b[280])^(a[108] & b[281])^(a[107] & b[282])^(a[106] & b[283])^(a[105] & b[284])^(a[104] & b[285])^(a[103] & b[286])^(a[102] & b[287])^(a[101] & b[288])^(a[100] & b[289])^(a[99] & b[290])^(a[98] & b[291])^(a[97] & b[292])^(a[96] & b[293])^(a[95] & b[294])^(a[94] & b[295])^(a[93] & b[296])^(a[92] & b[297])^(a[91] & b[298])^(a[90] & b[299])^(a[89] & b[300])^(a[88] & b[301])^(a[87] & b[302])^(a[86] & b[303])^(a[85] & b[304])^(a[84] & b[305])^(a[83] & b[306])^(a[82] & b[307])^(a[81] & b[308])^(a[80] & b[309])^(a[79] & b[310])^(a[78] & b[311])^(a[77] & b[312])^(a[76] & b[313])^(a[75] & b[314])^(a[74] & b[315])^(a[73] & b[316])^(a[72] & b[317])^(a[71] & b[318])^(a[70] & b[319])^(a[69] & b[320])^(a[68] & b[321])^(a[67] & b[322])^(a[66] & b[323])^(a[65] & b[324])^(a[64] & b[325])^(a[63] & b[326])^(a[62] & b[327])^(a[61] & b[328])^(a[60] & b[329])^(a[59] & b[330])^(a[58] & b[331])^(a[57] & b[332])^(a[56] & b[333])^(a[55] & b[334])^(a[54] & b[335])^(a[53] & b[336])^(a[52] & b[337])^(a[51] & b[338])^(a[50] & b[339])^(a[49] & b[340])^(a[48] & b[341])^(a[47] & b[342])^(a[46] & b[343])^(a[45] & b[344])^(a[44] & b[345])^(a[43] & b[346])^(a[42] & b[347])^(a[41] & b[348])^(a[40] & b[349])^(a[39] & b[350])^(a[38] & b[351])^(a[37] & b[352])^(a[36] & b[353])^(a[35] & b[354])^(a[34] & b[355])^(a[33] & b[356])^(a[32] & b[357])^(a[31] & b[358])^(a[30] & b[359])^(a[29] & b[360])^(a[28] & b[361])^(a[27] & b[362])^(a[26] & b[363])^(a[25] & b[364])^(a[24] & b[365])^(a[23] & b[366])^(a[22] & b[367])^(a[21] & b[368])^(a[20] & b[369])^(a[19] & b[370])^(a[18] & b[371])^(a[17] & b[372])^(a[16] & b[373])^(a[15] & b[374])^(a[14] & b[375])^(a[13] & b[376])^(a[12] & b[377])^(a[11] & b[378])^(a[10] & b[379])^(a[9] & b[380])^(a[8] & b[381])^(a[7] & b[382])^(a[6] & b[383])^(a[5] & b[384])^(a[4] & b[385])^(a[3] & b[386])^(a[2] & b[387])^(a[1] & b[388])^(a[0] & b[389]);
assign y[390] = (a[390] & b[0])^(a[389] & b[1])^(a[388] & b[2])^(a[387] & b[3])^(a[386] & b[4])^(a[385] & b[5])^(a[384] & b[6])^(a[383] & b[7])^(a[382] & b[8])^(a[381] & b[9])^(a[380] & b[10])^(a[379] & b[11])^(a[378] & b[12])^(a[377] & b[13])^(a[376] & b[14])^(a[375] & b[15])^(a[374] & b[16])^(a[373] & b[17])^(a[372] & b[18])^(a[371] & b[19])^(a[370] & b[20])^(a[369] & b[21])^(a[368] & b[22])^(a[367] & b[23])^(a[366] & b[24])^(a[365] & b[25])^(a[364] & b[26])^(a[363] & b[27])^(a[362] & b[28])^(a[361] & b[29])^(a[360] & b[30])^(a[359] & b[31])^(a[358] & b[32])^(a[357] & b[33])^(a[356] & b[34])^(a[355] & b[35])^(a[354] & b[36])^(a[353] & b[37])^(a[352] & b[38])^(a[351] & b[39])^(a[350] & b[40])^(a[349] & b[41])^(a[348] & b[42])^(a[347] & b[43])^(a[346] & b[44])^(a[345] & b[45])^(a[344] & b[46])^(a[343] & b[47])^(a[342] & b[48])^(a[341] & b[49])^(a[340] & b[50])^(a[339] & b[51])^(a[338] & b[52])^(a[337] & b[53])^(a[336] & b[54])^(a[335] & b[55])^(a[334] & b[56])^(a[333] & b[57])^(a[332] & b[58])^(a[331] & b[59])^(a[330] & b[60])^(a[329] & b[61])^(a[328] & b[62])^(a[327] & b[63])^(a[326] & b[64])^(a[325] & b[65])^(a[324] & b[66])^(a[323] & b[67])^(a[322] & b[68])^(a[321] & b[69])^(a[320] & b[70])^(a[319] & b[71])^(a[318] & b[72])^(a[317] & b[73])^(a[316] & b[74])^(a[315] & b[75])^(a[314] & b[76])^(a[313] & b[77])^(a[312] & b[78])^(a[311] & b[79])^(a[310] & b[80])^(a[309] & b[81])^(a[308] & b[82])^(a[307] & b[83])^(a[306] & b[84])^(a[305] & b[85])^(a[304] & b[86])^(a[303] & b[87])^(a[302] & b[88])^(a[301] & b[89])^(a[300] & b[90])^(a[299] & b[91])^(a[298] & b[92])^(a[297] & b[93])^(a[296] & b[94])^(a[295] & b[95])^(a[294] & b[96])^(a[293] & b[97])^(a[292] & b[98])^(a[291] & b[99])^(a[290] & b[100])^(a[289] & b[101])^(a[288] & b[102])^(a[287] & b[103])^(a[286] & b[104])^(a[285] & b[105])^(a[284] & b[106])^(a[283] & b[107])^(a[282] & b[108])^(a[281] & b[109])^(a[280] & b[110])^(a[279] & b[111])^(a[278] & b[112])^(a[277] & b[113])^(a[276] & b[114])^(a[275] & b[115])^(a[274] & b[116])^(a[273] & b[117])^(a[272] & b[118])^(a[271] & b[119])^(a[270] & b[120])^(a[269] & b[121])^(a[268] & b[122])^(a[267] & b[123])^(a[266] & b[124])^(a[265] & b[125])^(a[264] & b[126])^(a[263] & b[127])^(a[262] & b[128])^(a[261] & b[129])^(a[260] & b[130])^(a[259] & b[131])^(a[258] & b[132])^(a[257] & b[133])^(a[256] & b[134])^(a[255] & b[135])^(a[254] & b[136])^(a[253] & b[137])^(a[252] & b[138])^(a[251] & b[139])^(a[250] & b[140])^(a[249] & b[141])^(a[248] & b[142])^(a[247] & b[143])^(a[246] & b[144])^(a[245] & b[145])^(a[244] & b[146])^(a[243] & b[147])^(a[242] & b[148])^(a[241] & b[149])^(a[240] & b[150])^(a[239] & b[151])^(a[238] & b[152])^(a[237] & b[153])^(a[236] & b[154])^(a[235] & b[155])^(a[234] & b[156])^(a[233] & b[157])^(a[232] & b[158])^(a[231] & b[159])^(a[230] & b[160])^(a[229] & b[161])^(a[228] & b[162])^(a[227] & b[163])^(a[226] & b[164])^(a[225] & b[165])^(a[224] & b[166])^(a[223] & b[167])^(a[222] & b[168])^(a[221] & b[169])^(a[220] & b[170])^(a[219] & b[171])^(a[218] & b[172])^(a[217] & b[173])^(a[216] & b[174])^(a[215] & b[175])^(a[214] & b[176])^(a[213] & b[177])^(a[212] & b[178])^(a[211] & b[179])^(a[210] & b[180])^(a[209] & b[181])^(a[208] & b[182])^(a[207] & b[183])^(a[206] & b[184])^(a[205] & b[185])^(a[204] & b[186])^(a[203] & b[187])^(a[202] & b[188])^(a[201] & b[189])^(a[200] & b[190])^(a[199] & b[191])^(a[198] & b[192])^(a[197] & b[193])^(a[196] & b[194])^(a[195] & b[195])^(a[194] & b[196])^(a[193] & b[197])^(a[192] & b[198])^(a[191] & b[199])^(a[190] & b[200])^(a[189] & b[201])^(a[188] & b[202])^(a[187] & b[203])^(a[186] & b[204])^(a[185] & b[205])^(a[184] & b[206])^(a[183] & b[207])^(a[182] & b[208])^(a[181] & b[209])^(a[180] & b[210])^(a[179] & b[211])^(a[178] & b[212])^(a[177] & b[213])^(a[176] & b[214])^(a[175] & b[215])^(a[174] & b[216])^(a[173] & b[217])^(a[172] & b[218])^(a[171] & b[219])^(a[170] & b[220])^(a[169] & b[221])^(a[168] & b[222])^(a[167] & b[223])^(a[166] & b[224])^(a[165] & b[225])^(a[164] & b[226])^(a[163] & b[227])^(a[162] & b[228])^(a[161] & b[229])^(a[160] & b[230])^(a[159] & b[231])^(a[158] & b[232])^(a[157] & b[233])^(a[156] & b[234])^(a[155] & b[235])^(a[154] & b[236])^(a[153] & b[237])^(a[152] & b[238])^(a[151] & b[239])^(a[150] & b[240])^(a[149] & b[241])^(a[148] & b[242])^(a[147] & b[243])^(a[146] & b[244])^(a[145] & b[245])^(a[144] & b[246])^(a[143] & b[247])^(a[142] & b[248])^(a[141] & b[249])^(a[140] & b[250])^(a[139] & b[251])^(a[138] & b[252])^(a[137] & b[253])^(a[136] & b[254])^(a[135] & b[255])^(a[134] & b[256])^(a[133] & b[257])^(a[132] & b[258])^(a[131] & b[259])^(a[130] & b[260])^(a[129] & b[261])^(a[128] & b[262])^(a[127] & b[263])^(a[126] & b[264])^(a[125] & b[265])^(a[124] & b[266])^(a[123] & b[267])^(a[122] & b[268])^(a[121] & b[269])^(a[120] & b[270])^(a[119] & b[271])^(a[118] & b[272])^(a[117] & b[273])^(a[116] & b[274])^(a[115] & b[275])^(a[114] & b[276])^(a[113] & b[277])^(a[112] & b[278])^(a[111] & b[279])^(a[110] & b[280])^(a[109] & b[281])^(a[108] & b[282])^(a[107] & b[283])^(a[106] & b[284])^(a[105] & b[285])^(a[104] & b[286])^(a[103] & b[287])^(a[102] & b[288])^(a[101] & b[289])^(a[100] & b[290])^(a[99] & b[291])^(a[98] & b[292])^(a[97] & b[293])^(a[96] & b[294])^(a[95] & b[295])^(a[94] & b[296])^(a[93] & b[297])^(a[92] & b[298])^(a[91] & b[299])^(a[90] & b[300])^(a[89] & b[301])^(a[88] & b[302])^(a[87] & b[303])^(a[86] & b[304])^(a[85] & b[305])^(a[84] & b[306])^(a[83] & b[307])^(a[82] & b[308])^(a[81] & b[309])^(a[80] & b[310])^(a[79] & b[311])^(a[78] & b[312])^(a[77] & b[313])^(a[76] & b[314])^(a[75] & b[315])^(a[74] & b[316])^(a[73] & b[317])^(a[72] & b[318])^(a[71] & b[319])^(a[70] & b[320])^(a[69] & b[321])^(a[68] & b[322])^(a[67] & b[323])^(a[66] & b[324])^(a[65] & b[325])^(a[64] & b[326])^(a[63] & b[327])^(a[62] & b[328])^(a[61] & b[329])^(a[60] & b[330])^(a[59] & b[331])^(a[58] & b[332])^(a[57] & b[333])^(a[56] & b[334])^(a[55] & b[335])^(a[54] & b[336])^(a[53] & b[337])^(a[52] & b[338])^(a[51] & b[339])^(a[50] & b[340])^(a[49] & b[341])^(a[48] & b[342])^(a[47] & b[343])^(a[46] & b[344])^(a[45] & b[345])^(a[44] & b[346])^(a[43] & b[347])^(a[42] & b[348])^(a[41] & b[349])^(a[40] & b[350])^(a[39] & b[351])^(a[38] & b[352])^(a[37] & b[353])^(a[36] & b[354])^(a[35] & b[355])^(a[34] & b[356])^(a[33] & b[357])^(a[32] & b[358])^(a[31] & b[359])^(a[30] & b[360])^(a[29] & b[361])^(a[28] & b[362])^(a[27] & b[363])^(a[26] & b[364])^(a[25] & b[365])^(a[24] & b[366])^(a[23] & b[367])^(a[22] & b[368])^(a[21] & b[369])^(a[20] & b[370])^(a[19] & b[371])^(a[18] & b[372])^(a[17] & b[373])^(a[16] & b[374])^(a[15] & b[375])^(a[14] & b[376])^(a[13] & b[377])^(a[12] & b[378])^(a[11] & b[379])^(a[10] & b[380])^(a[9] & b[381])^(a[8] & b[382])^(a[7] & b[383])^(a[6] & b[384])^(a[5] & b[385])^(a[4] & b[386])^(a[3] & b[387])^(a[2] & b[388])^(a[1] & b[389])^(a[0] & b[390]);
assign y[391] = (a[391] & b[0])^(a[390] & b[1])^(a[389] & b[2])^(a[388] & b[3])^(a[387] & b[4])^(a[386] & b[5])^(a[385] & b[6])^(a[384] & b[7])^(a[383] & b[8])^(a[382] & b[9])^(a[381] & b[10])^(a[380] & b[11])^(a[379] & b[12])^(a[378] & b[13])^(a[377] & b[14])^(a[376] & b[15])^(a[375] & b[16])^(a[374] & b[17])^(a[373] & b[18])^(a[372] & b[19])^(a[371] & b[20])^(a[370] & b[21])^(a[369] & b[22])^(a[368] & b[23])^(a[367] & b[24])^(a[366] & b[25])^(a[365] & b[26])^(a[364] & b[27])^(a[363] & b[28])^(a[362] & b[29])^(a[361] & b[30])^(a[360] & b[31])^(a[359] & b[32])^(a[358] & b[33])^(a[357] & b[34])^(a[356] & b[35])^(a[355] & b[36])^(a[354] & b[37])^(a[353] & b[38])^(a[352] & b[39])^(a[351] & b[40])^(a[350] & b[41])^(a[349] & b[42])^(a[348] & b[43])^(a[347] & b[44])^(a[346] & b[45])^(a[345] & b[46])^(a[344] & b[47])^(a[343] & b[48])^(a[342] & b[49])^(a[341] & b[50])^(a[340] & b[51])^(a[339] & b[52])^(a[338] & b[53])^(a[337] & b[54])^(a[336] & b[55])^(a[335] & b[56])^(a[334] & b[57])^(a[333] & b[58])^(a[332] & b[59])^(a[331] & b[60])^(a[330] & b[61])^(a[329] & b[62])^(a[328] & b[63])^(a[327] & b[64])^(a[326] & b[65])^(a[325] & b[66])^(a[324] & b[67])^(a[323] & b[68])^(a[322] & b[69])^(a[321] & b[70])^(a[320] & b[71])^(a[319] & b[72])^(a[318] & b[73])^(a[317] & b[74])^(a[316] & b[75])^(a[315] & b[76])^(a[314] & b[77])^(a[313] & b[78])^(a[312] & b[79])^(a[311] & b[80])^(a[310] & b[81])^(a[309] & b[82])^(a[308] & b[83])^(a[307] & b[84])^(a[306] & b[85])^(a[305] & b[86])^(a[304] & b[87])^(a[303] & b[88])^(a[302] & b[89])^(a[301] & b[90])^(a[300] & b[91])^(a[299] & b[92])^(a[298] & b[93])^(a[297] & b[94])^(a[296] & b[95])^(a[295] & b[96])^(a[294] & b[97])^(a[293] & b[98])^(a[292] & b[99])^(a[291] & b[100])^(a[290] & b[101])^(a[289] & b[102])^(a[288] & b[103])^(a[287] & b[104])^(a[286] & b[105])^(a[285] & b[106])^(a[284] & b[107])^(a[283] & b[108])^(a[282] & b[109])^(a[281] & b[110])^(a[280] & b[111])^(a[279] & b[112])^(a[278] & b[113])^(a[277] & b[114])^(a[276] & b[115])^(a[275] & b[116])^(a[274] & b[117])^(a[273] & b[118])^(a[272] & b[119])^(a[271] & b[120])^(a[270] & b[121])^(a[269] & b[122])^(a[268] & b[123])^(a[267] & b[124])^(a[266] & b[125])^(a[265] & b[126])^(a[264] & b[127])^(a[263] & b[128])^(a[262] & b[129])^(a[261] & b[130])^(a[260] & b[131])^(a[259] & b[132])^(a[258] & b[133])^(a[257] & b[134])^(a[256] & b[135])^(a[255] & b[136])^(a[254] & b[137])^(a[253] & b[138])^(a[252] & b[139])^(a[251] & b[140])^(a[250] & b[141])^(a[249] & b[142])^(a[248] & b[143])^(a[247] & b[144])^(a[246] & b[145])^(a[245] & b[146])^(a[244] & b[147])^(a[243] & b[148])^(a[242] & b[149])^(a[241] & b[150])^(a[240] & b[151])^(a[239] & b[152])^(a[238] & b[153])^(a[237] & b[154])^(a[236] & b[155])^(a[235] & b[156])^(a[234] & b[157])^(a[233] & b[158])^(a[232] & b[159])^(a[231] & b[160])^(a[230] & b[161])^(a[229] & b[162])^(a[228] & b[163])^(a[227] & b[164])^(a[226] & b[165])^(a[225] & b[166])^(a[224] & b[167])^(a[223] & b[168])^(a[222] & b[169])^(a[221] & b[170])^(a[220] & b[171])^(a[219] & b[172])^(a[218] & b[173])^(a[217] & b[174])^(a[216] & b[175])^(a[215] & b[176])^(a[214] & b[177])^(a[213] & b[178])^(a[212] & b[179])^(a[211] & b[180])^(a[210] & b[181])^(a[209] & b[182])^(a[208] & b[183])^(a[207] & b[184])^(a[206] & b[185])^(a[205] & b[186])^(a[204] & b[187])^(a[203] & b[188])^(a[202] & b[189])^(a[201] & b[190])^(a[200] & b[191])^(a[199] & b[192])^(a[198] & b[193])^(a[197] & b[194])^(a[196] & b[195])^(a[195] & b[196])^(a[194] & b[197])^(a[193] & b[198])^(a[192] & b[199])^(a[191] & b[200])^(a[190] & b[201])^(a[189] & b[202])^(a[188] & b[203])^(a[187] & b[204])^(a[186] & b[205])^(a[185] & b[206])^(a[184] & b[207])^(a[183] & b[208])^(a[182] & b[209])^(a[181] & b[210])^(a[180] & b[211])^(a[179] & b[212])^(a[178] & b[213])^(a[177] & b[214])^(a[176] & b[215])^(a[175] & b[216])^(a[174] & b[217])^(a[173] & b[218])^(a[172] & b[219])^(a[171] & b[220])^(a[170] & b[221])^(a[169] & b[222])^(a[168] & b[223])^(a[167] & b[224])^(a[166] & b[225])^(a[165] & b[226])^(a[164] & b[227])^(a[163] & b[228])^(a[162] & b[229])^(a[161] & b[230])^(a[160] & b[231])^(a[159] & b[232])^(a[158] & b[233])^(a[157] & b[234])^(a[156] & b[235])^(a[155] & b[236])^(a[154] & b[237])^(a[153] & b[238])^(a[152] & b[239])^(a[151] & b[240])^(a[150] & b[241])^(a[149] & b[242])^(a[148] & b[243])^(a[147] & b[244])^(a[146] & b[245])^(a[145] & b[246])^(a[144] & b[247])^(a[143] & b[248])^(a[142] & b[249])^(a[141] & b[250])^(a[140] & b[251])^(a[139] & b[252])^(a[138] & b[253])^(a[137] & b[254])^(a[136] & b[255])^(a[135] & b[256])^(a[134] & b[257])^(a[133] & b[258])^(a[132] & b[259])^(a[131] & b[260])^(a[130] & b[261])^(a[129] & b[262])^(a[128] & b[263])^(a[127] & b[264])^(a[126] & b[265])^(a[125] & b[266])^(a[124] & b[267])^(a[123] & b[268])^(a[122] & b[269])^(a[121] & b[270])^(a[120] & b[271])^(a[119] & b[272])^(a[118] & b[273])^(a[117] & b[274])^(a[116] & b[275])^(a[115] & b[276])^(a[114] & b[277])^(a[113] & b[278])^(a[112] & b[279])^(a[111] & b[280])^(a[110] & b[281])^(a[109] & b[282])^(a[108] & b[283])^(a[107] & b[284])^(a[106] & b[285])^(a[105] & b[286])^(a[104] & b[287])^(a[103] & b[288])^(a[102] & b[289])^(a[101] & b[290])^(a[100] & b[291])^(a[99] & b[292])^(a[98] & b[293])^(a[97] & b[294])^(a[96] & b[295])^(a[95] & b[296])^(a[94] & b[297])^(a[93] & b[298])^(a[92] & b[299])^(a[91] & b[300])^(a[90] & b[301])^(a[89] & b[302])^(a[88] & b[303])^(a[87] & b[304])^(a[86] & b[305])^(a[85] & b[306])^(a[84] & b[307])^(a[83] & b[308])^(a[82] & b[309])^(a[81] & b[310])^(a[80] & b[311])^(a[79] & b[312])^(a[78] & b[313])^(a[77] & b[314])^(a[76] & b[315])^(a[75] & b[316])^(a[74] & b[317])^(a[73] & b[318])^(a[72] & b[319])^(a[71] & b[320])^(a[70] & b[321])^(a[69] & b[322])^(a[68] & b[323])^(a[67] & b[324])^(a[66] & b[325])^(a[65] & b[326])^(a[64] & b[327])^(a[63] & b[328])^(a[62] & b[329])^(a[61] & b[330])^(a[60] & b[331])^(a[59] & b[332])^(a[58] & b[333])^(a[57] & b[334])^(a[56] & b[335])^(a[55] & b[336])^(a[54] & b[337])^(a[53] & b[338])^(a[52] & b[339])^(a[51] & b[340])^(a[50] & b[341])^(a[49] & b[342])^(a[48] & b[343])^(a[47] & b[344])^(a[46] & b[345])^(a[45] & b[346])^(a[44] & b[347])^(a[43] & b[348])^(a[42] & b[349])^(a[41] & b[350])^(a[40] & b[351])^(a[39] & b[352])^(a[38] & b[353])^(a[37] & b[354])^(a[36] & b[355])^(a[35] & b[356])^(a[34] & b[357])^(a[33] & b[358])^(a[32] & b[359])^(a[31] & b[360])^(a[30] & b[361])^(a[29] & b[362])^(a[28] & b[363])^(a[27] & b[364])^(a[26] & b[365])^(a[25] & b[366])^(a[24] & b[367])^(a[23] & b[368])^(a[22] & b[369])^(a[21] & b[370])^(a[20] & b[371])^(a[19] & b[372])^(a[18] & b[373])^(a[17] & b[374])^(a[16] & b[375])^(a[15] & b[376])^(a[14] & b[377])^(a[13] & b[378])^(a[12] & b[379])^(a[11] & b[380])^(a[10] & b[381])^(a[9] & b[382])^(a[8] & b[383])^(a[7] & b[384])^(a[6] & b[385])^(a[5] & b[386])^(a[4] & b[387])^(a[3] & b[388])^(a[2] & b[389])^(a[1] & b[390])^(a[0] & b[391]);
assign y[392] = (a[392] & b[0])^(a[391] & b[1])^(a[390] & b[2])^(a[389] & b[3])^(a[388] & b[4])^(a[387] & b[5])^(a[386] & b[6])^(a[385] & b[7])^(a[384] & b[8])^(a[383] & b[9])^(a[382] & b[10])^(a[381] & b[11])^(a[380] & b[12])^(a[379] & b[13])^(a[378] & b[14])^(a[377] & b[15])^(a[376] & b[16])^(a[375] & b[17])^(a[374] & b[18])^(a[373] & b[19])^(a[372] & b[20])^(a[371] & b[21])^(a[370] & b[22])^(a[369] & b[23])^(a[368] & b[24])^(a[367] & b[25])^(a[366] & b[26])^(a[365] & b[27])^(a[364] & b[28])^(a[363] & b[29])^(a[362] & b[30])^(a[361] & b[31])^(a[360] & b[32])^(a[359] & b[33])^(a[358] & b[34])^(a[357] & b[35])^(a[356] & b[36])^(a[355] & b[37])^(a[354] & b[38])^(a[353] & b[39])^(a[352] & b[40])^(a[351] & b[41])^(a[350] & b[42])^(a[349] & b[43])^(a[348] & b[44])^(a[347] & b[45])^(a[346] & b[46])^(a[345] & b[47])^(a[344] & b[48])^(a[343] & b[49])^(a[342] & b[50])^(a[341] & b[51])^(a[340] & b[52])^(a[339] & b[53])^(a[338] & b[54])^(a[337] & b[55])^(a[336] & b[56])^(a[335] & b[57])^(a[334] & b[58])^(a[333] & b[59])^(a[332] & b[60])^(a[331] & b[61])^(a[330] & b[62])^(a[329] & b[63])^(a[328] & b[64])^(a[327] & b[65])^(a[326] & b[66])^(a[325] & b[67])^(a[324] & b[68])^(a[323] & b[69])^(a[322] & b[70])^(a[321] & b[71])^(a[320] & b[72])^(a[319] & b[73])^(a[318] & b[74])^(a[317] & b[75])^(a[316] & b[76])^(a[315] & b[77])^(a[314] & b[78])^(a[313] & b[79])^(a[312] & b[80])^(a[311] & b[81])^(a[310] & b[82])^(a[309] & b[83])^(a[308] & b[84])^(a[307] & b[85])^(a[306] & b[86])^(a[305] & b[87])^(a[304] & b[88])^(a[303] & b[89])^(a[302] & b[90])^(a[301] & b[91])^(a[300] & b[92])^(a[299] & b[93])^(a[298] & b[94])^(a[297] & b[95])^(a[296] & b[96])^(a[295] & b[97])^(a[294] & b[98])^(a[293] & b[99])^(a[292] & b[100])^(a[291] & b[101])^(a[290] & b[102])^(a[289] & b[103])^(a[288] & b[104])^(a[287] & b[105])^(a[286] & b[106])^(a[285] & b[107])^(a[284] & b[108])^(a[283] & b[109])^(a[282] & b[110])^(a[281] & b[111])^(a[280] & b[112])^(a[279] & b[113])^(a[278] & b[114])^(a[277] & b[115])^(a[276] & b[116])^(a[275] & b[117])^(a[274] & b[118])^(a[273] & b[119])^(a[272] & b[120])^(a[271] & b[121])^(a[270] & b[122])^(a[269] & b[123])^(a[268] & b[124])^(a[267] & b[125])^(a[266] & b[126])^(a[265] & b[127])^(a[264] & b[128])^(a[263] & b[129])^(a[262] & b[130])^(a[261] & b[131])^(a[260] & b[132])^(a[259] & b[133])^(a[258] & b[134])^(a[257] & b[135])^(a[256] & b[136])^(a[255] & b[137])^(a[254] & b[138])^(a[253] & b[139])^(a[252] & b[140])^(a[251] & b[141])^(a[250] & b[142])^(a[249] & b[143])^(a[248] & b[144])^(a[247] & b[145])^(a[246] & b[146])^(a[245] & b[147])^(a[244] & b[148])^(a[243] & b[149])^(a[242] & b[150])^(a[241] & b[151])^(a[240] & b[152])^(a[239] & b[153])^(a[238] & b[154])^(a[237] & b[155])^(a[236] & b[156])^(a[235] & b[157])^(a[234] & b[158])^(a[233] & b[159])^(a[232] & b[160])^(a[231] & b[161])^(a[230] & b[162])^(a[229] & b[163])^(a[228] & b[164])^(a[227] & b[165])^(a[226] & b[166])^(a[225] & b[167])^(a[224] & b[168])^(a[223] & b[169])^(a[222] & b[170])^(a[221] & b[171])^(a[220] & b[172])^(a[219] & b[173])^(a[218] & b[174])^(a[217] & b[175])^(a[216] & b[176])^(a[215] & b[177])^(a[214] & b[178])^(a[213] & b[179])^(a[212] & b[180])^(a[211] & b[181])^(a[210] & b[182])^(a[209] & b[183])^(a[208] & b[184])^(a[207] & b[185])^(a[206] & b[186])^(a[205] & b[187])^(a[204] & b[188])^(a[203] & b[189])^(a[202] & b[190])^(a[201] & b[191])^(a[200] & b[192])^(a[199] & b[193])^(a[198] & b[194])^(a[197] & b[195])^(a[196] & b[196])^(a[195] & b[197])^(a[194] & b[198])^(a[193] & b[199])^(a[192] & b[200])^(a[191] & b[201])^(a[190] & b[202])^(a[189] & b[203])^(a[188] & b[204])^(a[187] & b[205])^(a[186] & b[206])^(a[185] & b[207])^(a[184] & b[208])^(a[183] & b[209])^(a[182] & b[210])^(a[181] & b[211])^(a[180] & b[212])^(a[179] & b[213])^(a[178] & b[214])^(a[177] & b[215])^(a[176] & b[216])^(a[175] & b[217])^(a[174] & b[218])^(a[173] & b[219])^(a[172] & b[220])^(a[171] & b[221])^(a[170] & b[222])^(a[169] & b[223])^(a[168] & b[224])^(a[167] & b[225])^(a[166] & b[226])^(a[165] & b[227])^(a[164] & b[228])^(a[163] & b[229])^(a[162] & b[230])^(a[161] & b[231])^(a[160] & b[232])^(a[159] & b[233])^(a[158] & b[234])^(a[157] & b[235])^(a[156] & b[236])^(a[155] & b[237])^(a[154] & b[238])^(a[153] & b[239])^(a[152] & b[240])^(a[151] & b[241])^(a[150] & b[242])^(a[149] & b[243])^(a[148] & b[244])^(a[147] & b[245])^(a[146] & b[246])^(a[145] & b[247])^(a[144] & b[248])^(a[143] & b[249])^(a[142] & b[250])^(a[141] & b[251])^(a[140] & b[252])^(a[139] & b[253])^(a[138] & b[254])^(a[137] & b[255])^(a[136] & b[256])^(a[135] & b[257])^(a[134] & b[258])^(a[133] & b[259])^(a[132] & b[260])^(a[131] & b[261])^(a[130] & b[262])^(a[129] & b[263])^(a[128] & b[264])^(a[127] & b[265])^(a[126] & b[266])^(a[125] & b[267])^(a[124] & b[268])^(a[123] & b[269])^(a[122] & b[270])^(a[121] & b[271])^(a[120] & b[272])^(a[119] & b[273])^(a[118] & b[274])^(a[117] & b[275])^(a[116] & b[276])^(a[115] & b[277])^(a[114] & b[278])^(a[113] & b[279])^(a[112] & b[280])^(a[111] & b[281])^(a[110] & b[282])^(a[109] & b[283])^(a[108] & b[284])^(a[107] & b[285])^(a[106] & b[286])^(a[105] & b[287])^(a[104] & b[288])^(a[103] & b[289])^(a[102] & b[290])^(a[101] & b[291])^(a[100] & b[292])^(a[99] & b[293])^(a[98] & b[294])^(a[97] & b[295])^(a[96] & b[296])^(a[95] & b[297])^(a[94] & b[298])^(a[93] & b[299])^(a[92] & b[300])^(a[91] & b[301])^(a[90] & b[302])^(a[89] & b[303])^(a[88] & b[304])^(a[87] & b[305])^(a[86] & b[306])^(a[85] & b[307])^(a[84] & b[308])^(a[83] & b[309])^(a[82] & b[310])^(a[81] & b[311])^(a[80] & b[312])^(a[79] & b[313])^(a[78] & b[314])^(a[77] & b[315])^(a[76] & b[316])^(a[75] & b[317])^(a[74] & b[318])^(a[73] & b[319])^(a[72] & b[320])^(a[71] & b[321])^(a[70] & b[322])^(a[69] & b[323])^(a[68] & b[324])^(a[67] & b[325])^(a[66] & b[326])^(a[65] & b[327])^(a[64] & b[328])^(a[63] & b[329])^(a[62] & b[330])^(a[61] & b[331])^(a[60] & b[332])^(a[59] & b[333])^(a[58] & b[334])^(a[57] & b[335])^(a[56] & b[336])^(a[55] & b[337])^(a[54] & b[338])^(a[53] & b[339])^(a[52] & b[340])^(a[51] & b[341])^(a[50] & b[342])^(a[49] & b[343])^(a[48] & b[344])^(a[47] & b[345])^(a[46] & b[346])^(a[45] & b[347])^(a[44] & b[348])^(a[43] & b[349])^(a[42] & b[350])^(a[41] & b[351])^(a[40] & b[352])^(a[39] & b[353])^(a[38] & b[354])^(a[37] & b[355])^(a[36] & b[356])^(a[35] & b[357])^(a[34] & b[358])^(a[33] & b[359])^(a[32] & b[360])^(a[31] & b[361])^(a[30] & b[362])^(a[29] & b[363])^(a[28] & b[364])^(a[27] & b[365])^(a[26] & b[366])^(a[25] & b[367])^(a[24] & b[368])^(a[23] & b[369])^(a[22] & b[370])^(a[21] & b[371])^(a[20] & b[372])^(a[19] & b[373])^(a[18] & b[374])^(a[17] & b[375])^(a[16] & b[376])^(a[15] & b[377])^(a[14] & b[378])^(a[13] & b[379])^(a[12] & b[380])^(a[11] & b[381])^(a[10] & b[382])^(a[9] & b[383])^(a[8] & b[384])^(a[7] & b[385])^(a[6] & b[386])^(a[5] & b[387])^(a[4] & b[388])^(a[3] & b[389])^(a[2] & b[390])^(a[1] & b[391])^(a[0] & b[392]);
assign y[393] = (a[393] & b[0])^(a[392] & b[1])^(a[391] & b[2])^(a[390] & b[3])^(a[389] & b[4])^(a[388] & b[5])^(a[387] & b[6])^(a[386] & b[7])^(a[385] & b[8])^(a[384] & b[9])^(a[383] & b[10])^(a[382] & b[11])^(a[381] & b[12])^(a[380] & b[13])^(a[379] & b[14])^(a[378] & b[15])^(a[377] & b[16])^(a[376] & b[17])^(a[375] & b[18])^(a[374] & b[19])^(a[373] & b[20])^(a[372] & b[21])^(a[371] & b[22])^(a[370] & b[23])^(a[369] & b[24])^(a[368] & b[25])^(a[367] & b[26])^(a[366] & b[27])^(a[365] & b[28])^(a[364] & b[29])^(a[363] & b[30])^(a[362] & b[31])^(a[361] & b[32])^(a[360] & b[33])^(a[359] & b[34])^(a[358] & b[35])^(a[357] & b[36])^(a[356] & b[37])^(a[355] & b[38])^(a[354] & b[39])^(a[353] & b[40])^(a[352] & b[41])^(a[351] & b[42])^(a[350] & b[43])^(a[349] & b[44])^(a[348] & b[45])^(a[347] & b[46])^(a[346] & b[47])^(a[345] & b[48])^(a[344] & b[49])^(a[343] & b[50])^(a[342] & b[51])^(a[341] & b[52])^(a[340] & b[53])^(a[339] & b[54])^(a[338] & b[55])^(a[337] & b[56])^(a[336] & b[57])^(a[335] & b[58])^(a[334] & b[59])^(a[333] & b[60])^(a[332] & b[61])^(a[331] & b[62])^(a[330] & b[63])^(a[329] & b[64])^(a[328] & b[65])^(a[327] & b[66])^(a[326] & b[67])^(a[325] & b[68])^(a[324] & b[69])^(a[323] & b[70])^(a[322] & b[71])^(a[321] & b[72])^(a[320] & b[73])^(a[319] & b[74])^(a[318] & b[75])^(a[317] & b[76])^(a[316] & b[77])^(a[315] & b[78])^(a[314] & b[79])^(a[313] & b[80])^(a[312] & b[81])^(a[311] & b[82])^(a[310] & b[83])^(a[309] & b[84])^(a[308] & b[85])^(a[307] & b[86])^(a[306] & b[87])^(a[305] & b[88])^(a[304] & b[89])^(a[303] & b[90])^(a[302] & b[91])^(a[301] & b[92])^(a[300] & b[93])^(a[299] & b[94])^(a[298] & b[95])^(a[297] & b[96])^(a[296] & b[97])^(a[295] & b[98])^(a[294] & b[99])^(a[293] & b[100])^(a[292] & b[101])^(a[291] & b[102])^(a[290] & b[103])^(a[289] & b[104])^(a[288] & b[105])^(a[287] & b[106])^(a[286] & b[107])^(a[285] & b[108])^(a[284] & b[109])^(a[283] & b[110])^(a[282] & b[111])^(a[281] & b[112])^(a[280] & b[113])^(a[279] & b[114])^(a[278] & b[115])^(a[277] & b[116])^(a[276] & b[117])^(a[275] & b[118])^(a[274] & b[119])^(a[273] & b[120])^(a[272] & b[121])^(a[271] & b[122])^(a[270] & b[123])^(a[269] & b[124])^(a[268] & b[125])^(a[267] & b[126])^(a[266] & b[127])^(a[265] & b[128])^(a[264] & b[129])^(a[263] & b[130])^(a[262] & b[131])^(a[261] & b[132])^(a[260] & b[133])^(a[259] & b[134])^(a[258] & b[135])^(a[257] & b[136])^(a[256] & b[137])^(a[255] & b[138])^(a[254] & b[139])^(a[253] & b[140])^(a[252] & b[141])^(a[251] & b[142])^(a[250] & b[143])^(a[249] & b[144])^(a[248] & b[145])^(a[247] & b[146])^(a[246] & b[147])^(a[245] & b[148])^(a[244] & b[149])^(a[243] & b[150])^(a[242] & b[151])^(a[241] & b[152])^(a[240] & b[153])^(a[239] & b[154])^(a[238] & b[155])^(a[237] & b[156])^(a[236] & b[157])^(a[235] & b[158])^(a[234] & b[159])^(a[233] & b[160])^(a[232] & b[161])^(a[231] & b[162])^(a[230] & b[163])^(a[229] & b[164])^(a[228] & b[165])^(a[227] & b[166])^(a[226] & b[167])^(a[225] & b[168])^(a[224] & b[169])^(a[223] & b[170])^(a[222] & b[171])^(a[221] & b[172])^(a[220] & b[173])^(a[219] & b[174])^(a[218] & b[175])^(a[217] & b[176])^(a[216] & b[177])^(a[215] & b[178])^(a[214] & b[179])^(a[213] & b[180])^(a[212] & b[181])^(a[211] & b[182])^(a[210] & b[183])^(a[209] & b[184])^(a[208] & b[185])^(a[207] & b[186])^(a[206] & b[187])^(a[205] & b[188])^(a[204] & b[189])^(a[203] & b[190])^(a[202] & b[191])^(a[201] & b[192])^(a[200] & b[193])^(a[199] & b[194])^(a[198] & b[195])^(a[197] & b[196])^(a[196] & b[197])^(a[195] & b[198])^(a[194] & b[199])^(a[193] & b[200])^(a[192] & b[201])^(a[191] & b[202])^(a[190] & b[203])^(a[189] & b[204])^(a[188] & b[205])^(a[187] & b[206])^(a[186] & b[207])^(a[185] & b[208])^(a[184] & b[209])^(a[183] & b[210])^(a[182] & b[211])^(a[181] & b[212])^(a[180] & b[213])^(a[179] & b[214])^(a[178] & b[215])^(a[177] & b[216])^(a[176] & b[217])^(a[175] & b[218])^(a[174] & b[219])^(a[173] & b[220])^(a[172] & b[221])^(a[171] & b[222])^(a[170] & b[223])^(a[169] & b[224])^(a[168] & b[225])^(a[167] & b[226])^(a[166] & b[227])^(a[165] & b[228])^(a[164] & b[229])^(a[163] & b[230])^(a[162] & b[231])^(a[161] & b[232])^(a[160] & b[233])^(a[159] & b[234])^(a[158] & b[235])^(a[157] & b[236])^(a[156] & b[237])^(a[155] & b[238])^(a[154] & b[239])^(a[153] & b[240])^(a[152] & b[241])^(a[151] & b[242])^(a[150] & b[243])^(a[149] & b[244])^(a[148] & b[245])^(a[147] & b[246])^(a[146] & b[247])^(a[145] & b[248])^(a[144] & b[249])^(a[143] & b[250])^(a[142] & b[251])^(a[141] & b[252])^(a[140] & b[253])^(a[139] & b[254])^(a[138] & b[255])^(a[137] & b[256])^(a[136] & b[257])^(a[135] & b[258])^(a[134] & b[259])^(a[133] & b[260])^(a[132] & b[261])^(a[131] & b[262])^(a[130] & b[263])^(a[129] & b[264])^(a[128] & b[265])^(a[127] & b[266])^(a[126] & b[267])^(a[125] & b[268])^(a[124] & b[269])^(a[123] & b[270])^(a[122] & b[271])^(a[121] & b[272])^(a[120] & b[273])^(a[119] & b[274])^(a[118] & b[275])^(a[117] & b[276])^(a[116] & b[277])^(a[115] & b[278])^(a[114] & b[279])^(a[113] & b[280])^(a[112] & b[281])^(a[111] & b[282])^(a[110] & b[283])^(a[109] & b[284])^(a[108] & b[285])^(a[107] & b[286])^(a[106] & b[287])^(a[105] & b[288])^(a[104] & b[289])^(a[103] & b[290])^(a[102] & b[291])^(a[101] & b[292])^(a[100] & b[293])^(a[99] & b[294])^(a[98] & b[295])^(a[97] & b[296])^(a[96] & b[297])^(a[95] & b[298])^(a[94] & b[299])^(a[93] & b[300])^(a[92] & b[301])^(a[91] & b[302])^(a[90] & b[303])^(a[89] & b[304])^(a[88] & b[305])^(a[87] & b[306])^(a[86] & b[307])^(a[85] & b[308])^(a[84] & b[309])^(a[83] & b[310])^(a[82] & b[311])^(a[81] & b[312])^(a[80] & b[313])^(a[79] & b[314])^(a[78] & b[315])^(a[77] & b[316])^(a[76] & b[317])^(a[75] & b[318])^(a[74] & b[319])^(a[73] & b[320])^(a[72] & b[321])^(a[71] & b[322])^(a[70] & b[323])^(a[69] & b[324])^(a[68] & b[325])^(a[67] & b[326])^(a[66] & b[327])^(a[65] & b[328])^(a[64] & b[329])^(a[63] & b[330])^(a[62] & b[331])^(a[61] & b[332])^(a[60] & b[333])^(a[59] & b[334])^(a[58] & b[335])^(a[57] & b[336])^(a[56] & b[337])^(a[55] & b[338])^(a[54] & b[339])^(a[53] & b[340])^(a[52] & b[341])^(a[51] & b[342])^(a[50] & b[343])^(a[49] & b[344])^(a[48] & b[345])^(a[47] & b[346])^(a[46] & b[347])^(a[45] & b[348])^(a[44] & b[349])^(a[43] & b[350])^(a[42] & b[351])^(a[41] & b[352])^(a[40] & b[353])^(a[39] & b[354])^(a[38] & b[355])^(a[37] & b[356])^(a[36] & b[357])^(a[35] & b[358])^(a[34] & b[359])^(a[33] & b[360])^(a[32] & b[361])^(a[31] & b[362])^(a[30] & b[363])^(a[29] & b[364])^(a[28] & b[365])^(a[27] & b[366])^(a[26] & b[367])^(a[25] & b[368])^(a[24] & b[369])^(a[23] & b[370])^(a[22] & b[371])^(a[21] & b[372])^(a[20] & b[373])^(a[19] & b[374])^(a[18] & b[375])^(a[17] & b[376])^(a[16] & b[377])^(a[15] & b[378])^(a[14] & b[379])^(a[13] & b[380])^(a[12] & b[381])^(a[11] & b[382])^(a[10] & b[383])^(a[9] & b[384])^(a[8] & b[385])^(a[7] & b[386])^(a[6] & b[387])^(a[5] & b[388])^(a[4] & b[389])^(a[3] & b[390])^(a[2] & b[391])^(a[1] & b[392])^(a[0] & b[393]);
assign y[394] = (a[394] & b[0])^(a[393] & b[1])^(a[392] & b[2])^(a[391] & b[3])^(a[390] & b[4])^(a[389] & b[5])^(a[388] & b[6])^(a[387] & b[7])^(a[386] & b[8])^(a[385] & b[9])^(a[384] & b[10])^(a[383] & b[11])^(a[382] & b[12])^(a[381] & b[13])^(a[380] & b[14])^(a[379] & b[15])^(a[378] & b[16])^(a[377] & b[17])^(a[376] & b[18])^(a[375] & b[19])^(a[374] & b[20])^(a[373] & b[21])^(a[372] & b[22])^(a[371] & b[23])^(a[370] & b[24])^(a[369] & b[25])^(a[368] & b[26])^(a[367] & b[27])^(a[366] & b[28])^(a[365] & b[29])^(a[364] & b[30])^(a[363] & b[31])^(a[362] & b[32])^(a[361] & b[33])^(a[360] & b[34])^(a[359] & b[35])^(a[358] & b[36])^(a[357] & b[37])^(a[356] & b[38])^(a[355] & b[39])^(a[354] & b[40])^(a[353] & b[41])^(a[352] & b[42])^(a[351] & b[43])^(a[350] & b[44])^(a[349] & b[45])^(a[348] & b[46])^(a[347] & b[47])^(a[346] & b[48])^(a[345] & b[49])^(a[344] & b[50])^(a[343] & b[51])^(a[342] & b[52])^(a[341] & b[53])^(a[340] & b[54])^(a[339] & b[55])^(a[338] & b[56])^(a[337] & b[57])^(a[336] & b[58])^(a[335] & b[59])^(a[334] & b[60])^(a[333] & b[61])^(a[332] & b[62])^(a[331] & b[63])^(a[330] & b[64])^(a[329] & b[65])^(a[328] & b[66])^(a[327] & b[67])^(a[326] & b[68])^(a[325] & b[69])^(a[324] & b[70])^(a[323] & b[71])^(a[322] & b[72])^(a[321] & b[73])^(a[320] & b[74])^(a[319] & b[75])^(a[318] & b[76])^(a[317] & b[77])^(a[316] & b[78])^(a[315] & b[79])^(a[314] & b[80])^(a[313] & b[81])^(a[312] & b[82])^(a[311] & b[83])^(a[310] & b[84])^(a[309] & b[85])^(a[308] & b[86])^(a[307] & b[87])^(a[306] & b[88])^(a[305] & b[89])^(a[304] & b[90])^(a[303] & b[91])^(a[302] & b[92])^(a[301] & b[93])^(a[300] & b[94])^(a[299] & b[95])^(a[298] & b[96])^(a[297] & b[97])^(a[296] & b[98])^(a[295] & b[99])^(a[294] & b[100])^(a[293] & b[101])^(a[292] & b[102])^(a[291] & b[103])^(a[290] & b[104])^(a[289] & b[105])^(a[288] & b[106])^(a[287] & b[107])^(a[286] & b[108])^(a[285] & b[109])^(a[284] & b[110])^(a[283] & b[111])^(a[282] & b[112])^(a[281] & b[113])^(a[280] & b[114])^(a[279] & b[115])^(a[278] & b[116])^(a[277] & b[117])^(a[276] & b[118])^(a[275] & b[119])^(a[274] & b[120])^(a[273] & b[121])^(a[272] & b[122])^(a[271] & b[123])^(a[270] & b[124])^(a[269] & b[125])^(a[268] & b[126])^(a[267] & b[127])^(a[266] & b[128])^(a[265] & b[129])^(a[264] & b[130])^(a[263] & b[131])^(a[262] & b[132])^(a[261] & b[133])^(a[260] & b[134])^(a[259] & b[135])^(a[258] & b[136])^(a[257] & b[137])^(a[256] & b[138])^(a[255] & b[139])^(a[254] & b[140])^(a[253] & b[141])^(a[252] & b[142])^(a[251] & b[143])^(a[250] & b[144])^(a[249] & b[145])^(a[248] & b[146])^(a[247] & b[147])^(a[246] & b[148])^(a[245] & b[149])^(a[244] & b[150])^(a[243] & b[151])^(a[242] & b[152])^(a[241] & b[153])^(a[240] & b[154])^(a[239] & b[155])^(a[238] & b[156])^(a[237] & b[157])^(a[236] & b[158])^(a[235] & b[159])^(a[234] & b[160])^(a[233] & b[161])^(a[232] & b[162])^(a[231] & b[163])^(a[230] & b[164])^(a[229] & b[165])^(a[228] & b[166])^(a[227] & b[167])^(a[226] & b[168])^(a[225] & b[169])^(a[224] & b[170])^(a[223] & b[171])^(a[222] & b[172])^(a[221] & b[173])^(a[220] & b[174])^(a[219] & b[175])^(a[218] & b[176])^(a[217] & b[177])^(a[216] & b[178])^(a[215] & b[179])^(a[214] & b[180])^(a[213] & b[181])^(a[212] & b[182])^(a[211] & b[183])^(a[210] & b[184])^(a[209] & b[185])^(a[208] & b[186])^(a[207] & b[187])^(a[206] & b[188])^(a[205] & b[189])^(a[204] & b[190])^(a[203] & b[191])^(a[202] & b[192])^(a[201] & b[193])^(a[200] & b[194])^(a[199] & b[195])^(a[198] & b[196])^(a[197] & b[197])^(a[196] & b[198])^(a[195] & b[199])^(a[194] & b[200])^(a[193] & b[201])^(a[192] & b[202])^(a[191] & b[203])^(a[190] & b[204])^(a[189] & b[205])^(a[188] & b[206])^(a[187] & b[207])^(a[186] & b[208])^(a[185] & b[209])^(a[184] & b[210])^(a[183] & b[211])^(a[182] & b[212])^(a[181] & b[213])^(a[180] & b[214])^(a[179] & b[215])^(a[178] & b[216])^(a[177] & b[217])^(a[176] & b[218])^(a[175] & b[219])^(a[174] & b[220])^(a[173] & b[221])^(a[172] & b[222])^(a[171] & b[223])^(a[170] & b[224])^(a[169] & b[225])^(a[168] & b[226])^(a[167] & b[227])^(a[166] & b[228])^(a[165] & b[229])^(a[164] & b[230])^(a[163] & b[231])^(a[162] & b[232])^(a[161] & b[233])^(a[160] & b[234])^(a[159] & b[235])^(a[158] & b[236])^(a[157] & b[237])^(a[156] & b[238])^(a[155] & b[239])^(a[154] & b[240])^(a[153] & b[241])^(a[152] & b[242])^(a[151] & b[243])^(a[150] & b[244])^(a[149] & b[245])^(a[148] & b[246])^(a[147] & b[247])^(a[146] & b[248])^(a[145] & b[249])^(a[144] & b[250])^(a[143] & b[251])^(a[142] & b[252])^(a[141] & b[253])^(a[140] & b[254])^(a[139] & b[255])^(a[138] & b[256])^(a[137] & b[257])^(a[136] & b[258])^(a[135] & b[259])^(a[134] & b[260])^(a[133] & b[261])^(a[132] & b[262])^(a[131] & b[263])^(a[130] & b[264])^(a[129] & b[265])^(a[128] & b[266])^(a[127] & b[267])^(a[126] & b[268])^(a[125] & b[269])^(a[124] & b[270])^(a[123] & b[271])^(a[122] & b[272])^(a[121] & b[273])^(a[120] & b[274])^(a[119] & b[275])^(a[118] & b[276])^(a[117] & b[277])^(a[116] & b[278])^(a[115] & b[279])^(a[114] & b[280])^(a[113] & b[281])^(a[112] & b[282])^(a[111] & b[283])^(a[110] & b[284])^(a[109] & b[285])^(a[108] & b[286])^(a[107] & b[287])^(a[106] & b[288])^(a[105] & b[289])^(a[104] & b[290])^(a[103] & b[291])^(a[102] & b[292])^(a[101] & b[293])^(a[100] & b[294])^(a[99] & b[295])^(a[98] & b[296])^(a[97] & b[297])^(a[96] & b[298])^(a[95] & b[299])^(a[94] & b[300])^(a[93] & b[301])^(a[92] & b[302])^(a[91] & b[303])^(a[90] & b[304])^(a[89] & b[305])^(a[88] & b[306])^(a[87] & b[307])^(a[86] & b[308])^(a[85] & b[309])^(a[84] & b[310])^(a[83] & b[311])^(a[82] & b[312])^(a[81] & b[313])^(a[80] & b[314])^(a[79] & b[315])^(a[78] & b[316])^(a[77] & b[317])^(a[76] & b[318])^(a[75] & b[319])^(a[74] & b[320])^(a[73] & b[321])^(a[72] & b[322])^(a[71] & b[323])^(a[70] & b[324])^(a[69] & b[325])^(a[68] & b[326])^(a[67] & b[327])^(a[66] & b[328])^(a[65] & b[329])^(a[64] & b[330])^(a[63] & b[331])^(a[62] & b[332])^(a[61] & b[333])^(a[60] & b[334])^(a[59] & b[335])^(a[58] & b[336])^(a[57] & b[337])^(a[56] & b[338])^(a[55] & b[339])^(a[54] & b[340])^(a[53] & b[341])^(a[52] & b[342])^(a[51] & b[343])^(a[50] & b[344])^(a[49] & b[345])^(a[48] & b[346])^(a[47] & b[347])^(a[46] & b[348])^(a[45] & b[349])^(a[44] & b[350])^(a[43] & b[351])^(a[42] & b[352])^(a[41] & b[353])^(a[40] & b[354])^(a[39] & b[355])^(a[38] & b[356])^(a[37] & b[357])^(a[36] & b[358])^(a[35] & b[359])^(a[34] & b[360])^(a[33] & b[361])^(a[32] & b[362])^(a[31] & b[363])^(a[30] & b[364])^(a[29] & b[365])^(a[28] & b[366])^(a[27] & b[367])^(a[26] & b[368])^(a[25] & b[369])^(a[24] & b[370])^(a[23] & b[371])^(a[22] & b[372])^(a[21] & b[373])^(a[20] & b[374])^(a[19] & b[375])^(a[18] & b[376])^(a[17] & b[377])^(a[16] & b[378])^(a[15] & b[379])^(a[14] & b[380])^(a[13] & b[381])^(a[12] & b[382])^(a[11] & b[383])^(a[10] & b[384])^(a[9] & b[385])^(a[8] & b[386])^(a[7] & b[387])^(a[6] & b[388])^(a[5] & b[389])^(a[4] & b[390])^(a[3] & b[391])^(a[2] & b[392])^(a[1] & b[393])^(a[0] & b[394]);
assign y[395] = (a[395] & b[0])^(a[394] & b[1])^(a[393] & b[2])^(a[392] & b[3])^(a[391] & b[4])^(a[390] & b[5])^(a[389] & b[6])^(a[388] & b[7])^(a[387] & b[8])^(a[386] & b[9])^(a[385] & b[10])^(a[384] & b[11])^(a[383] & b[12])^(a[382] & b[13])^(a[381] & b[14])^(a[380] & b[15])^(a[379] & b[16])^(a[378] & b[17])^(a[377] & b[18])^(a[376] & b[19])^(a[375] & b[20])^(a[374] & b[21])^(a[373] & b[22])^(a[372] & b[23])^(a[371] & b[24])^(a[370] & b[25])^(a[369] & b[26])^(a[368] & b[27])^(a[367] & b[28])^(a[366] & b[29])^(a[365] & b[30])^(a[364] & b[31])^(a[363] & b[32])^(a[362] & b[33])^(a[361] & b[34])^(a[360] & b[35])^(a[359] & b[36])^(a[358] & b[37])^(a[357] & b[38])^(a[356] & b[39])^(a[355] & b[40])^(a[354] & b[41])^(a[353] & b[42])^(a[352] & b[43])^(a[351] & b[44])^(a[350] & b[45])^(a[349] & b[46])^(a[348] & b[47])^(a[347] & b[48])^(a[346] & b[49])^(a[345] & b[50])^(a[344] & b[51])^(a[343] & b[52])^(a[342] & b[53])^(a[341] & b[54])^(a[340] & b[55])^(a[339] & b[56])^(a[338] & b[57])^(a[337] & b[58])^(a[336] & b[59])^(a[335] & b[60])^(a[334] & b[61])^(a[333] & b[62])^(a[332] & b[63])^(a[331] & b[64])^(a[330] & b[65])^(a[329] & b[66])^(a[328] & b[67])^(a[327] & b[68])^(a[326] & b[69])^(a[325] & b[70])^(a[324] & b[71])^(a[323] & b[72])^(a[322] & b[73])^(a[321] & b[74])^(a[320] & b[75])^(a[319] & b[76])^(a[318] & b[77])^(a[317] & b[78])^(a[316] & b[79])^(a[315] & b[80])^(a[314] & b[81])^(a[313] & b[82])^(a[312] & b[83])^(a[311] & b[84])^(a[310] & b[85])^(a[309] & b[86])^(a[308] & b[87])^(a[307] & b[88])^(a[306] & b[89])^(a[305] & b[90])^(a[304] & b[91])^(a[303] & b[92])^(a[302] & b[93])^(a[301] & b[94])^(a[300] & b[95])^(a[299] & b[96])^(a[298] & b[97])^(a[297] & b[98])^(a[296] & b[99])^(a[295] & b[100])^(a[294] & b[101])^(a[293] & b[102])^(a[292] & b[103])^(a[291] & b[104])^(a[290] & b[105])^(a[289] & b[106])^(a[288] & b[107])^(a[287] & b[108])^(a[286] & b[109])^(a[285] & b[110])^(a[284] & b[111])^(a[283] & b[112])^(a[282] & b[113])^(a[281] & b[114])^(a[280] & b[115])^(a[279] & b[116])^(a[278] & b[117])^(a[277] & b[118])^(a[276] & b[119])^(a[275] & b[120])^(a[274] & b[121])^(a[273] & b[122])^(a[272] & b[123])^(a[271] & b[124])^(a[270] & b[125])^(a[269] & b[126])^(a[268] & b[127])^(a[267] & b[128])^(a[266] & b[129])^(a[265] & b[130])^(a[264] & b[131])^(a[263] & b[132])^(a[262] & b[133])^(a[261] & b[134])^(a[260] & b[135])^(a[259] & b[136])^(a[258] & b[137])^(a[257] & b[138])^(a[256] & b[139])^(a[255] & b[140])^(a[254] & b[141])^(a[253] & b[142])^(a[252] & b[143])^(a[251] & b[144])^(a[250] & b[145])^(a[249] & b[146])^(a[248] & b[147])^(a[247] & b[148])^(a[246] & b[149])^(a[245] & b[150])^(a[244] & b[151])^(a[243] & b[152])^(a[242] & b[153])^(a[241] & b[154])^(a[240] & b[155])^(a[239] & b[156])^(a[238] & b[157])^(a[237] & b[158])^(a[236] & b[159])^(a[235] & b[160])^(a[234] & b[161])^(a[233] & b[162])^(a[232] & b[163])^(a[231] & b[164])^(a[230] & b[165])^(a[229] & b[166])^(a[228] & b[167])^(a[227] & b[168])^(a[226] & b[169])^(a[225] & b[170])^(a[224] & b[171])^(a[223] & b[172])^(a[222] & b[173])^(a[221] & b[174])^(a[220] & b[175])^(a[219] & b[176])^(a[218] & b[177])^(a[217] & b[178])^(a[216] & b[179])^(a[215] & b[180])^(a[214] & b[181])^(a[213] & b[182])^(a[212] & b[183])^(a[211] & b[184])^(a[210] & b[185])^(a[209] & b[186])^(a[208] & b[187])^(a[207] & b[188])^(a[206] & b[189])^(a[205] & b[190])^(a[204] & b[191])^(a[203] & b[192])^(a[202] & b[193])^(a[201] & b[194])^(a[200] & b[195])^(a[199] & b[196])^(a[198] & b[197])^(a[197] & b[198])^(a[196] & b[199])^(a[195] & b[200])^(a[194] & b[201])^(a[193] & b[202])^(a[192] & b[203])^(a[191] & b[204])^(a[190] & b[205])^(a[189] & b[206])^(a[188] & b[207])^(a[187] & b[208])^(a[186] & b[209])^(a[185] & b[210])^(a[184] & b[211])^(a[183] & b[212])^(a[182] & b[213])^(a[181] & b[214])^(a[180] & b[215])^(a[179] & b[216])^(a[178] & b[217])^(a[177] & b[218])^(a[176] & b[219])^(a[175] & b[220])^(a[174] & b[221])^(a[173] & b[222])^(a[172] & b[223])^(a[171] & b[224])^(a[170] & b[225])^(a[169] & b[226])^(a[168] & b[227])^(a[167] & b[228])^(a[166] & b[229])^(a[165] & b[230])^(a[164] & b[231])^(a[163] & b[232])^(a[162] & b[233])^(a[161] & b[234])^(a[160] & b[235])^(a[159] & b[236])^(a[158] & b[237])^(a[157] & b[238])^(a[156] & b[239])^(a[155] & b[240])^(a[154] & b[241])^(a[153] & b[242])^(a[152] & b[243])^(a[151] & b[244])^(a[150] & b[245])^(a[149] & b[246])^(a[148] & b[247])^(a[147] & b[248])^(a[146] & b[249])^(a[145] & b[250])^(a[144] & b[251])^(a[143] & b[252])^(a[142] & b[253])^(a[141] & b[254])^(a[140] & b[255])^(a[139] & b[256])^(a[138] & b[257])^(a[137] & b[258])^(a[136] & b[259])^(a[135] & b[260])^(a[134] & b[261])^(a[133] & b[262])^(a[132] & b[263])^(a[131] & b[264])^(a[130] & b[265])^(a[129] & b[266])^(a[128] & b[267])^(a[127] & b[268])^(a[126] & b[269])^(a[125] & b[270])^(a[124] & b[271])^(a[123] & b[272])^(a[122] & b[273])^(a[121] & b[274])^(a[120] & b[275])^(a[119] & b[276])^(a[118] & b[277])^(a[117] & b[278])^(a[116] & b[279])^(a[115] & b[280])^(a[114] & b[281])^(a[113] & b[282])^(a[112] & b[283])^(a[111] & b[284])^(a[110] & b[285])^(a[109] & b[286])^(a[108] & b[287])^(a[107] & b[288])^(a[106] & b[289])^(a[105] & b[290])^(a[104] & b[291])^(a[103] & b[292])^(a[102] & b[293])^(a[101] & b[294])^(a[100] & b[295])^(a[99] & b[296])^(a[98] & b[297])^(a[97] & b[298])^(a[96] & b[299])^(a[95] & b[300])^(a[94] & b[301])^(a[93] & b[302])^(a[92] & b[303])^(a[91] & b[304])^(a[90] & b[305])^(a[89] & b[306])^(a[88] & b[307])^(a[87] & b[308])^(a[86] & b[309])^(a[85] & b[310])^(a[84] & b[311])^(a[83] & b[312])^(a[82] & b[313])^(a[81] & b[314])^(a[80] & b[315])^(a[79] & b[316])^(a[78] & b[317])^(a[77] & b[318])^(a[76] & b[319])^(a[75] & b[320])^(a[74] & b[321])^(a[73] & b[322])^(a[72] & b[323])^(a[71] & b[324])^(a[70] & b[325])^(a[69] & b[326])^(a[68] & b[327])^(a[67] & b[328])^(a[66] & b[329])^(a[65] & b[330])^(a[64] & b[331])^(a[63] & b[332])^(a[62] & b[333])^(a[61] & b[334])^(a[60] & b[335])^(a[59] & b[336])^(a[58] & b[337])^(a[57] & b[338])^(a[56] & b[339])^(a[55] & b[340])^(a[54] & b[341])^(a[53] & b[342])^(a[52] & b[343])^(a[51] & b[344])^(a[50] & b[345])^(a[49] & b[346])^(a[48] & b[347])^(a[47] & b[348])^(a[46] & b[349])^(a[45] & b[350])^(a[44] & b[351])^(a[43] & b[352])^(a[42] & b[353])^(a[41] & b[354])^(a[40] & b[355])^(a[39] & b[356])^(a[38] & b[357])^(a[37] & b[358])^(a[36] & b[359])^(a[35] & b[360])^(a[34] & b[361])^(a[33] & b[362])^(a[32] & b[363])^(a[31] & b[364])^(a[30] & b[365])^(a[29] & b[366])^(a[28] & b[367])^(a[27] & b[368])^(a[26] & b[369])^(a[25] & b[370])^(a[24] & b[371])^(a[23] & b[372])^(a[22] & b[373])^(a[21] & b[374])^(a[20] & b[375])^(a[19] & b[376])^(a[18] & b[377])^(a[17] & b[378])^(a[16] & b[379])^(a[15] & b[380])^(a[14] & b[381])^(a[13] & b[382])^(a[12] & b[383])^(a[11] & b[384])^(a[10] & b[385])^(a[9] & b[386])^(a[8] & b[387])^(a[7] & b[388])^(a[6] & b[389])^(a[5] & b[390])^(a[4] & b[391])^(a[3] & b[392])^(a[2] & b[393])^(a[1] & b[394])^(a[0] & b[395]);
assign y[396] = (a[396] & b[0])^(a[395] & b[1])^(a[394] & b[2])^(a[393] & b[3])^(a[392] & b[4])^(a[391] & b[5])^(a[390] & b[6])^(a[389] & b[7])^(a[388] & b[8])^(a[387] & b[9])^(a[386] & b[10])^(a[385] & b[11])^(a[384] & b[12])^(a[383] & b[13])^(a[382] & b[14])^(a[381] & b[15])^(a[380] & b[16])^(a[379] & b[17])^(a[378] & b[18])^(a[377] & b[19])^(a[376] & b[20])^(a[375] & b[21])^(a[374] & b[22])^(a[373] & b[23])^(a[372] & b[24])^(a[371] & b[25])^(a[370] & b[26])^(a[369] & b[27])^(a[368] & b[28])^(a[367] & b[29])^(a[366] & b[30])^(a[365] & b[31])^(a[364] & b[32])^(a[363] & b[33])^(a[362] & b[34])^(a[361] & b[35])^(a[360] & b[36])^(a[359] & b[37])^(a[358] & b[38])^(a[357] & b[39])^(a[356] & b[40])^(a[355] & b[41])^(a[354] & b[42])^(a[353] & b[43])^(a[352] & b[44])^(a[351] & b[45])^(a[350] & b[46])^(a[349] & b[47])^(a[348] & b[48])^(a[347] & b[49])^(a[346] & b[50])^(a[345] & b[51])^(a[344] & b[52])^(a[343] & b[53])^(a[342] & b[54])^(a[341] & b[55])^(a[340] & b[56])^(a[339] & b[57])^(a[338] & b[58])^(a[337] & b[59])^(a[336] & b[60])^(a[335] & b[61])^(a[334] & b[62])^(a[333] & b[63])^(a[332] & b[64])^(a[331] & b[65])^(a[330] & b[66])^(a[329] & b[67])^(a[328] & b[68])^(a[327] & b[69])^(a[326] & b[70])^(a[325] & b[71])^(a[324] & b[72])^(a[323] & b[73])^(a[322] & b[74])^(a[321] & b[75])^(a[320] & b[76])^(a[319] & b[77])^(a[318] & b[78])^(a[317] & b[79])^(a[316] & b[80])^(a[315] & b[81])^(a[314] & b[82])^(a[313] & b[83])^(a[312] & b[84])^(a[311] & b[85])^(a[310] & b[86])^(a[309] & b[87])^(a[308] & b[88])^(a[307] & b[89])^(a[306] & b[90])^(a[305] & b[91])^(a[304] & b[92])^(a[303] & b[93])^(a[302] & b[94])^(a[301] & b[95])^(a[300] & b[96])^(a[299] & b[97])^(a[298] & b[98])^(a[297] & b[99])^(a[296] & b[100])^(a[295] & b[101])^(a[294] & b[102])^(a[293] & b[103])^(a[292] & b[104])^(a[291] & b[105])^(a[290] & b[106])^(a[289] & b[107])^(a[288] & b[108])^(a[287] & b[109])^(a[286] & b[110])^(a[285] & b[111])^(a[284] & b[112])^(a[283] & b[113])^(a[282] & b[114])^(a[281] & b[115])^(a[280] & b[116])^(a[279] & b[117])^(a[278] & b[118])^(a[277] & b[119])^(a[276] & b[120])^(a[275] & b[121])^(a[274] & b[122])^(a[273] & b[123])^(a[272] & b[124])^(a[271] & b[125])^(a[270] & b[126])^(a[269] & b[127])^(a[268] & b[128])^(a[267] & b[129])^(a[266] & b[130])^(a[265] & b[131])^(a[264] & b[132])^(a[263] & b[133])^(a[262] & b[134])^(a[261] & b[135])^(a[260] & b[136])^(a[259] & b[137])^(a[258] & b[138])^(a[257] & b[139])^(a[256] & b[140])^(a[255] & b[141])^(a[254] & b[142])^(a[253] & b[143])^(a[252] & b[144])^(a[251] & b[145])^(a[250] & b[146])^(a[249] & b[147])^(a[248] & b[148])^(a[247] & b[149])^(a[246] & b[150])^(a[245] & b[151])^(a[244] & b[152])^(a[243] & b[153])^(a[242] & b[154])^(a[241] & b[155])^(a[240] & b[156])^(a[239] & b[157])^(a[238] & b[158])^(a[237] & b[159])^(a[236] & b[160])^(a[235] & b[161])^(a[234] & b[162])^(a[233] & b[163])^(a[232] & b[164])^(a[231] & b[165])^(a[230] & b[166])^(a[229] & b[167])^(a[228] & b[168])^(a[227] & b[169])^(a[226] & b[170])^(a[225] & b[171])^(a[224] & b[172])^(a[223] & b[173])^(a[222] & b[174])^(a[221] & b[175])^(a[220] & b[176])^(a[219] & b[177])^(a[218] & b[178])^(a[217] & b[179])^(a[216] & b[180])^(a[215] & b[181])^(a[214] & b[182])^(a[213] & b[183])^(a[212] & b[184])^(a[211] & b[185])^(a[210] & b[186])^(a[209] & b[187])^(a[208] & b[188])^(a[207] & b[189])^(a[206] & b[190])^(a[205] & b[191])^(a[204] & b[192])^(a[203] & b[193])^(a[202] & b[194])^(a[201] & b[195])^(a[200] & b[196])^(a[199] & b[197])^(a[198] & b[198])^(a[197] & b[199])^(a[196] & b[200])^(a[195] & b[201])^(a[194] & b[202])^(a[193] & b[203])^(a[192] & b[204])^(a[191] & b[205])^(a[190] & b[206])^(a[189] & b[207])^(a[188] & b[208])^(a[187] & b[209])^(a[186] & b[210])^(a[185] & b[211])^(a[184] & b[212])^(a[183] & b[213])^(a[182] & b[214])^(a[181] & b[215])^(a[180] & b[216])^(a[179] & b[217])^(a[178] & b[218])^(a[177] & b[219])^(a[176] & b[220])^(a[175] & b[221])^(a[174] & b[222])^(a[173] & b[223])^(a[172] & b[224])^(a[171] & b[225])^(a[170] & b[226])^(a[169] & b[227])^(a[168] & b[228])^(a[167] & b[229])^(a[166] & b[230])^(a[165] & b[231])^(a[164] & b[232])^(a[163] & b[233])^(a[162] & b[234])^(a[161] & b[235])^(a[160] & b[236])^(a[159] & b[237])^(a[158] & b[238])^(a[157] & b[239])^(a[156] & b[240])^(a[155] & b[241])^(a[154] & b[242])^(a[153] & b[243])^(a[152] & b[244])^(a[151] & b[245])^(a[150] & b[246])^(a[149] & b[247])^(a[148] & b[248])^(a[147] & b[249])^(a[146] & b[250])^(a[145] & b[251])^(a[144] & b[252])^(a[143] & b[253])^(a[142] & b[254])^(a[141] & b[255])^(a[140] & b[256])^(a[139] & b[257])^(a[138] & b[258])^(a[137] & b[259])^(a[136] & b[260])^(a[135] & b[261])^(a[134] & b[262])^(a[133] & b[263])^(a[132] & b[264])^(a[131] & b[265])^(a[130] & b[266])^(a[129] & b[267])^(a[128] & b[268])^(a[127] & b[269])^(a[126] & b[270])^(a[125] & b[271])^(a[124] & b[272])^(a[123] & b[273])^(a[122] & b[274])^(a[121] & b[275])^(a[120] & b[276])^(a[119] & b[277])^(a[118] & b[278])^(a[117] & b[279])^(a[116] & b[280])^(a[115] & b[281])^(a[114] & b[282])^(a[113] & b[283])^(a[112] & b[284])^(a[111] & b[285])^(a[110] & b[286])^(a[109] & b[287])^(a[108] & b[288])^(a[107] & b[289])^(a[106] & b[290])^(a[105] & b[291])^(a[104] & b[292])^(a[103] & b[293])^(a[102] & b[294])^(a[101] & b[295])^(a[100] & b[296])^(a[99] & b[297])^(a[98] & b[298])^(a[97] & b[299])^(a[96] & b[300])^(a[95] & b[301])^(a[94] & b[302])^(a[93] & b[303])^(a[92] & b[304])^(a[91] & b[305])^(a[90] & b[306])^(a[89] & b[307])^(a[88] & b[308])^(a[87] & b[309])^(a[86] & b[310])^(a[85] & b[311])^(a[84] & b[312])^(a[83] & b[313])^(a[82] & b[314])^(a[81] & b[315])^(a[80] & b[316])^(a[79] & b[317])^(a[78] & b[318])^(a[77] & b[319])^(a[76] & b[320])^(a[75] & b[321])^(a[74] & b[322])^(a[73] & b[323])^(a[72] & b[324])^(a[71] & b[325])^(a[70] & b[326])^(a[69] & b[327])^(a[68] & b[328])^(a[67] & b[329])^(a[66] & b[330])^(a[65] & b[331])^(a[64] & b[332])^(a[63] & b[333])^(a[62] & b[334])^(a[61] & b[335])^(a[60] & b[336])^(a[59] & b[337])^(a[58] & b[338])^(a[57] & b[339])^(a[56] & b[340])^(a[55] & b[341])^(a[54] & b[342])^(a[53] & b[343])^(a[52] & b[344])^(a[51] & b[345])^(a[50] & b[346])^(a[49] & b[347])^(a[48] & b[348])^(a[47] & b[349])^(a[46] & b[350])^(a[45] & b[351])^(a[44] & b[352])^(a[43] & b[353])^(a[42] & b[354])^(a[41] & b[355])^(a[40] & b[356])^(a[39] & b[357])^(a[38] & b[358])^(a[37] & b[359])^(a[36] & b[360])^(a[35] & b[361])^(a[34] & b[362])^(a[33] & b[363])^(a[32] & b[364])^(a[31] & b[365])^(a[30] & b[366])^(a[29] & b[367])^(a[28] & b[368])^(a[27] & b[369])^(a[26] & b[370])^(a[25] & b[371])^(a[24] & b[372])^(a[23] & b[373])^(a[22] & b[374])^(a[21] & b[375])^(a[20] & b[376])^(a[19] & b[377])^(a[18] & b[378])^(a[17] & b[379])^(a[16] & b[380])^(a[15] & b[381])^(a[14] & b[382])^(a[13] & b[383])^(a[12] & b[384])^(a[11] & b[385])^(a[10] & b[386])^(a[9] & b[387])^(a[8] & b[388])^(a[7] & b[389])^(a[6] & b[390])^(a[5] & b[391])^(a[4] & b[392])^(a[3] & b[393])^(a[2] & b[394])^(a[1] & b[395])^(a[0] & b[396]);
assign y[397] = (a[397] & b[0])^(a[396] & b[1])^(a[395] & b[2])^(a[394] & b[3])^(a[393] & b[4])^(a[392] & b[5])^(a[391] & b[6])^(a[390] & b[7])^(a[389] & b[8])^(a[388] & b[9])^(a[387] & b[10])^(a[386] & b[11])^(a[385] & b[12])^(a[384] & b[13])^(a[383] & b[14])^(a[382] & b[15])^(a[381] & b[16])^(a[380] & b[17])^(a[379] & b[18])^(a[378] & b[19])^(a[377] & b[20])^(a[376] & b[21])^(a[375] & b[22])^(a[374] & b[23])^(a[373] & b[24])^(a[372] & b[25])^(a[371] & b[26])^(a[370] & b[27])^(a[369] & b[28])^(a[368] & b[29])^(a[367] & b[30])^(a[366] & b[31])^(a[365] & b[32])^(a[364] & b[33])^(a[363] & b[34])^(a[362] & b[35])^(a[361] & b[36])^(a[360] & b[37])^(a[359] & b[38])^(a[358] & b[39])^(a[357] & b[40])^(a[356] & b[41])^(a[355] & b[42])^(a[354] & b[43])^(a[353] & b[44])^(a[352] & b[45])^(a[351] & b[46])^(a[350] & b[47])^(a[349] & b[48])^(a[348] & b[49])^(a[347] & b[50])^(a[346] & b[51])^(a[345] & b[52])^(a[344] & b[53])^(a[343] & b[54])^(a[342] & b[55])^(a[341] & b[56])^(a[340] & b[57])^(a[339] & b[58])^(a[338] & b[59])^(a[337] & b[60])^(a[336] & b[61])^(a[335] & b[62])^(a[334] & b[63])^(a[333] & b[64])^(a[332] & b[65])^(a[331] & b[66])^(a[330] & b[67])^(a[329] & b[68])^(a[328] & b[69])^(a[327] & b[70])^(a[326] & b[71])^(a[325] & b[72])^(a[324] & b[73])^(a[323] & b[74])^(a[322] & b[75])^(a[321] & b[76])^(a[320] & b[77])^(a[319] & b[78])^(a[318] & b[79])^(a[317] & b[80])^(a[316] & b[81])^(a[315] & b[82])^(a[314] & b[83])^(a[313] & b[84])^(a[312] & b[85])^(a[311] & b[86])^(a[310] & b[87])^(a[309] & b[88])^(a[308] & b[89])^(a[307] & b[90])^(a[306] & b[91])^(a[305] & b[92])^(a[304] & b[93])^(a[303] & b[94])^(a[302] & b[95])^(a[301] & b[96])^(a[300] & b[97])^(a[299] & b[98])^(a[298] & b[99])^(a[297] & b[100])^(a[296] & b[101])^(a[295] & b[102])^(a[294] & b[103])^(a[293] & b[104])^(a[292] & b[105])^(a[291] & b[106])^(a[290] & b[107])^(a[289] & b[108])^(a[288] & b[109])^(a[287] & b[110])^(a[286] & b[111])^(a[285] & b[112])^(a[284] & b[113])^(a[283] & b[114])^(a[282] & b[115])^(a[281] & b[116])^(a[280] & b[117])^(a[279] & b[118])^(a[278] & b[119])^(a[277] & b[120])^(a[276] & b[121])^(a[275] & b[122])^(a[274] & b[123])^(a[273] & b[124])^(a[272] & b[125])^(a[271] & b[126])^(a[270] & b[127])^(a[269] & b[128])^(a[268] & b[129])^(a[267] & b[130])^(a[266] & b[131])^(a[265] & b[132])^(a[264] & b[133])^(a[263] & b[134])^(a[262] & b[135])^(a[261] & b[136])^(a[260] & b[137])^(a[259] & b[138])^(a[258] & b[139])^(a[257] & b[140])^(a[256] & b[141])^(a[255] & b[142])^(a[254] & b[143])^(a[253] & b[144])^(a[252] & b[145])^(a[251] & b[146])^(a[250] & b[147])^(a[249] & b[148])^(a[248] & b[149])^(a[247] & b[150])^(a[246] & b[151])^(a[245] & b[152])^(a[244] & b[153])^(a[243] & b[154])^(a[242] & b[155])^(a[241] & b[156])^(a[240] & b[157])^(a[239] & b[158])^(a[238] & b[159])^(a[237] & b[160])^(a[236] & b[161])^(a[235] & b[162])^(a[234] & b[163])^(a[233] & b[164])^(a[232] & b[165])^(a[231] & b[166])^(a[230] & b[167])^(a[229] & b[168])^(a[228] & b[169])^(a[227] & b[170])^(a[226] & b[171])^(a[225] & b[172])^(a[224] & b[173])^(a[223] & b[174])^(a[222] & b[175])^(a[221] & b[176])^(a[220] & b[177])^(a[219] & b[178])^(a[218] & b[179])^(a[217] & b[180])^(a[216] & b[181])^(a[215] & b[182])^(a[214] & b[183])^(a[213] & b[184])^(a[212] & b[185])^(a[211] & b[186])^(a[210] & b[187])^(a[209] & b[188])^(a[208] & b[189])^(a[207] & b[190])^(a[206] & b[191])^(a[205] & b[192])^(a[204] & b[193])^(a[203] & b[194])^(a[202] & b[195])^(a[201] & b[196])^(a[200] & b[197])^(a[199] & b[198])^(a[198] & b[199])^(a[197] & b[200])^(a[196] & b[201])^(a[195] & b[202])^(a[194] & b[203])^(a[193] & b[204])^(a[192] & b[205])^(a[191] & b[206])^(a[190] & b[207])^(a[189] & b[208])^(a[188] & b[209])^(a[187] & b[210])^(a[186] & b[211])^(a[185] & b[212])^(a[184] & b[213])^(a[183] & b[214])^(a[182] & b[215])^(a[181] & b[216])^(a[180] & b[217])^(a[179] & b[218])^(a[178] & b[219])^(a[177] & b[220])^(a[176] & b[221])^(a[175] & b[222])^(a[174] & b[223])^(a[173] & b[224])^(a[172] & b[225])^(a[171] & b[226])^(a[170] & b[227])^(a[169] & b[228])^(a[168] & b[229])^(a[167] & b[230])^(a[166] & b[231])^(a[165] & b[232])^(a[164] & b[233])^(a[163] & b[234])^(a[162] & b[235])^(a[161] & b[236])^(a[160] & b[237])^(a[159] & b[238])^(a[158] & b[239])^(a[157] & b[240])^(a[156] & b[241])^(a[155] & b[242])^(a[154] & b[243])^(a[153] & b[244])^(a[152] & b[245])^(a[151] & b[246])^(a[150] & b[247])^(a[149] & b[248])^(a[148] & b[249])^(a[147] & b[250])^(a[146] & b[251])^(a[145] & b[252])^(a[144] & b[253])^(a[143] & b[254])^(a[142] & b[255])^(a[141] & b[256])^(a[140] & b[257])^(a[139] & b[258])^(a[138] & b[259])^(a[137] & b[260])^(a[136] & b[261])^(a[135] & b[262])^(a[134] & b[263])^(a[133] & b[264])^(a[132] & b[265])^(a[131] & b[266])^(a[130] & b[267])^(a[129] & b[268])^(a[128] & b[269])^(a[127] & b[270])^(a[126] & b[271])^(a[125] & b[272])^(a[124] & b[273])^(a[123] & b[274])^(a[122] & b[275])^(a[121] & b[276])^(a[120] & b[277])^(a[119] & b[278])^(a[118] & b[279])^(a[117] & b[280])^(a[116] & b[281])^(a[115] & b[282])^(a[114] & b[283])^(a[113] & b[284])^(a[112] & b[285])^(a[111] & b[286])^(a[110] & b[287])^(a[109] & b[288])^(a[108] & b[289])^(a[107] & b[290])^(a[106] & b[291])^(a[105] & b[292])^(a[104] & b[293])^(a[103] & b[294])^(a[102] & b[295])^(a[101] & b[296])^(a[100] & b[297])^(a[99] & b[298])^(a[98] & b[299])^(a[97] & b[300])^(a[96] & b[301])^(a[95] & b[302])^(a[94] & b[303])^(a[93] & b[304])^(a[92] & b[305])^(a[91] & b[306])^(a[90] & b[307])^(a[89] & b[308])^(a[88] & b[309])^(a[87] & b[310])^(a[86] & b[311])^(a[85] & b[312])^(a[84] & b[313])^(a[83] & b[314])^(a[82] & b[315])^(a[81] & b[316])^(a[80] & b[317])^(a[79] & b[318])^(a[78] & b[319])^(a[77] & b[320])^(a[76] & b[321])^(a[75] & b[322])^(a[74] & b[323])^(a[73] & b[324])^(a[72] & b[325])^(a[71] & b[326])^(a[70] & b[327])^(a[69] & b[328])^(a[68] & b[329])^(a[67] & b[330])^(a[66] & b[331])^(a[65] & b[332])^(a[64] & b[333])^(a[63] & b[334])^(a[62] & b[335])^(a[61] & b[336])^(a[60] & b[337])^(a[59] & b[338])^(a[58] & b[339])^(a[57] & b[340])^(a[56] & b[341])^(a[55] & b[342])^(a[54] & b[343])^(a[53] & b[344])^(a[52] & b[345])^(a[51] & b[346])^(a[50] & b[347])^(a[49] & b[348])^(a[48] & b[349])^(a[47] & b[350])^(a[46] & b[351])^(a[45] & b[352])^(a[44] & b[353])^(a[43] & b[354])^(a[42] & b[355])^(a[41] & b[356])^(a[40] & b[357])^(a[39] & b[358])^(a[38] & b[359])^(a[37] & b[360])^(a[36] & b[361])^(a[35] & b[362])^(a[34] & b[363])^(a[33] & b[364])^(a[32] & b[365])^(a[31] & b[366])^(a[30] & b[367])^(a[29] & b[368])^(a[28] & b[369])^(a[27] & b[370])^(a[26] & b[371])^(a[25] & b[372])^(a[24] & b[373])^(a[23] & b[374])^(a[22] & b[375])^(a[21] & b[376])^(a[20] & b[377])^(a[19] & b[378])^(a[18] & b[379])^(a[17] & b[380])^(a[16] & b[381])^(a[15] & b[382])^(a[14] & b[383])^(a[13] & b[384])^(a[12] & b[385])^(a[11] & b[386])^(a[10] & b[387])^(a[9] & b[388])^(a[8] & b[389])^(a[7] & b[390])^(a[6] & b[391])^(a[5] & b[392])^(a[4] & b[393])^(a[3] & b[394])^(a[2] & b[395])^(a[1] & b[396])^(a[0] & b[397]);
assign y[398] = (a[398] & b[0])^(a[397] & b[1])^(a[396] & b[2])^(a[395] & b[3])^(a[394] & b[4])^(a[393] & b[5])^(a[392] & b[6])^(a[391] & b[7])^(a[390] & b[8])^(a[389] & b[9])^(a[388] & b[10])^(a[387] & b[11])^(a[386] & b[12])^(a[385] & b[13])^(a[384] & b[14])^(a[383] & b[15])^(a[382] & b[16])^(a[381] & b[17])^(a[380] & b[18])^(a[379] & b[19])^(a[378] & b[20])^(a[377] & b[21])^(a[376] & b[22])^(a[375] & b[23])^(a[374] & b[24])^(a[373] & b[25])^(a[372] & b[26])^(a[371] & b[27])^(a[370] & b[28])^(a[369] & b[29])^(a[368] & b[30])^(a[367] & b[31])^(a[366] & b[32])^(a[365] & b[33])^(a[364] & b[34])^(a[363] & b[35])^(a[362] & b[36])^(a[361] & b[37])^(a[360] & b[38])^(a[359] & b[39])^(a[358] & b[40])^(a[357] & b[41])^(a[356] & b[42])^(a[355] & b[43])^(a[354] & b[44])^(a[353] & b[45])^(a[352] & b[46])^(a[351] & b[47])^(a[350] & b[48])^(a[349] & b[49])^(a[348] & b[50])^(a[347] & b[51])^(a[346] & b[52])^(a[345] & b[53])^(a[344] & b[54])^(a[343] & b[55])^(a[342] & b[56])^(a[341] & b[57])^(a[340] & b[58])^(a[339] & b[59])^(a[338] & b[60])^(a[337] & b[61])^(a[336] & b[62])^(a[335] & b[63])^(a[334] & b[64])^(a[333] & b[65])^(a[332] & b[66])^(a[331] & b[67])^(a[330] & b[68])^(a[329] & b[69])^(a[328] & b[70])^(a[327] & b[71])^(a[326] & b[72])^(a[325] & b[73])^(a[324] & b[74])^(a[323] & b[75])^(a[322] & b[76])^(a[321] & b[77])^(a[320] & b[78])^(a[319] & b[79])^(a[318] & b[80])^(a[317] & b[81])^(a[316] & b[82])^(a[315] & b[83])^(a[314] & b[84])^(a[313] & b[85])^(a[312] & b[86])^(a[311] & b[87])^(a[310] & b[88])^(a[309] & b[89])^(a[308] & b[90])^(a[307] & b[91])^(a[306] & b[92])^(a[305] & b[93])^(a[304] & b[94])^(a[303] & b[95])^(a[302] & b[96])^(a[301] & b[97])^(a[300] & b[98])^(a[299] & b[99])^(a[298] & b[100])^(a[297] & b[101])^(a[296] & b[102])^(a[295] & b[103])^(a[294] & b[104])^(a[293] & b[105])^(a[292] & b[106])^(a[291] & b[107])^(a[290] & b[108])^(a[289] & b[109])^(a[288] & b[110])^(a[287] & b[111])^(a[286] & b[112])^(a[285] & b[113])^(a[284] & b[114])^(a[283] & b[115])^(a[282] & b[116])^(a[281] & b[117])^(a[280] & b[118])^(a[279] & b[119])^(a[278] & b[120])^(a[277] & b[121])^(a[276] & b[122])^(a[275] & b[123])^(a[274] & b[124])^(a[273] & b[125])^(a[272] & b[126])^(a[271] & b[127])^(a[270] & b[128])^(a[269] & b[129])^(a[268] & b[130])^(a[267] & b[131])^(a[266] & b[132])^(a[265] & b[133])^(a[264] & b[134])^(a[263] & b[135])^(a[262] & b[136])^(a[261] & b[137])^(a[260] & b[138])^(a[259] & b[139])^(a[258] & b[140])^(a[257] & b[141])^(a[256] & b[142])^(a[255] & b[143])^(a[254] & b[144])^(a[253] & b[145])^(a[252] & b[146])^(a[251] & b[147])^(a[250] & b[148])^(a[249] & b[149])^(a[248] & b[150])^(a[247] & b[151])^(a[246] & b[152])^(a[245] & b[153])^(a[244] & b[154])^(a[243] & b[155])^(a[242] & b[156])^(a[241] & b[157])^(a[240] & b[158])^(a[239] & b[159])^(a[238] & b[160])^(a[237] & b[161])^(a[236] & b[162])^(a[235] & b[163])^(a[234] & b[164])^(a[233] & b[165])^(a[232] & b[166])^(a[231] & b[167])^(a[230] & b[168])^(a[229] & b[169])^(a[228] & b[170])^(a[227] & b[171])^(a[226] & b[172])^(a[225] & b[173])^(a[224] & b[174])^(a[223] & b[175])^(a[222] & b[176])^(a[221] & b[177])^(a[220] & b[178])^(a[219] & b[179])^(a[218] & b[180])^(a[217] & b[181])^(a[216] & b[182])^(a[215] & b[183])^(a[214] & b[184])^(a[213] & b[185])^(a[212] & b[186])^(a[211] & b[187])^(a[210] & b[188])^(a[209] & b[189])^(a[208] & b[190])^(a[207] & b[191])^(a[206] & b[192])^(a[205] & b[193])^(a[204] & b[194])^(a[203] & b[195])^(a[202] & b[196])^(a[201] & b[197])^(a[200] & b[198])^(a[199] & b[199])^(a[198] & b[200])^(a[197] & b[201])^(a[196] & b[202])^(a[195] & b[203])^(a[194] & b[204])^(a[193] & b[205])^(a[192] & b[206])^(a[191] & b[207])^(a[190] & b[208])^(a[189] & b[209])^(a[188] & b[210])^(a[187] & b[211])^(a[186] & b[212])^(a[185] & b[213])^(a[184] & b[214])^(a[183] & b[215])^(a[182] & b[216])^(a[181] & b[217])^(a[180] & b[218])^(a[179] & b[219])^(a[178] & b[220])^(a[177] & b[221])^(a[176] & b[222])^(a[175] & b[223])^(a[174] & b[224])^(a[173] & b[225])^(a[172] & b[226])^(a[171] & b[227])^(a[170] & b[228])^(a[169] & b[229])^(a[168] & b[230])^(a[167] & b[231])^(a[166] & b[232])^(a[165] & b[233])^(a[164] & b[234])^(a[163] & b[235])^(a[162] & b[236])^(a[161] & b[237])^(a[160] & b[238])^(a[159] & b[239])^(a[158] & b[240])^(a[157] & b[241])^(a[156] & b[242])^(a[155] & b[243])^(a[154] & b[244])^(a[153] & b[245])^(a[152] & b[246])^(a[151] & b[247])^(a[150] & b[248])^(a[149] & b[249])^(a[148] & b[250])^(a[147] & b[251])^(a[146] & b[252])^(a[145] & b[253])^(a[144] & b[254])^(a[143] & b[255])^(a[142] & b[256])^(a[141] & b[257])^(a[140] & b[258])^(a[139] & b[259])^(a[138] & b[260])^(a[137] & b[261])^(a[136] & b[262])^(a[135] & b[263])^(a[134] & b[264])^(a[133] & b[265])^(a[132] & b[266])^(a[131] & b[267])^(a[130] & b[268])^(a[129] & b[269])^(a[128] & b[270])^(a[127] & b[271])^(a[126] & b[272])^(a[125] & b[273])^(a[124] & b[274])^(a[123] & b[275])^(a[122] & b[276])^(a[121] & b[277])^(a[120] & b[278])^(a[119] & b[279])^(a[118] & b[280])^(a[117] & b[281])^(a[116] & b[282])^(a[115] & b[283])^(a[114] & b[284])^(a[113] & b[285])^(a[112] & b[286])^(a[111] & b[287])^(a[110] & b[288])^(a[109] & b[289])^(a[108] & b[290])^(a[107] & b[291])^(a[106] & b[292])^(a[105] & b[293])^(a[104] & b[294])^(a[103] & b[295])^(a[102] & b[296])^(a[101] & b[297])^(a[100] & b[298])^(a[99] & b[299])^(a[98] & b[300])^(a[97] & b[301])^(a[96] & b[302])^(a[95] & b[303])^(a[94] & b[304])^(a[93] & b[305])^(a[92] & b[306])^(a[91] & b[307])^(a[90] & b[308])^(a[89] & b[309])^(a[88] & b[310])^(a[87] & b[311])^(a[86] & b[312])^(a[85] & b[313])^(a[84] & b[314])^(a[83] & b[315])^(a[82] & b[316])^(a[81] & b[317])^(a[80] & b[318])^(a[79] & b[319])^(a[78] & b[320])^(a[77] & b[321])^(a[76] & b[322])^(a[75] & b[323])^(a[74] & b[324])^(a[73] & b[325])^(a[72] & b[326])^(a[71] & b[327])^(a[70] & b[328])^(a[69] & b[329])^(a[68] & b[330])^(a[67] & b[331])^(a[66] & b[332])^(a[65] & b[333])^(a[64] & b[334])^(a[63] & b[335])^(a[62] & b[336])^(a[61] & b[337])^(a[60] & b[338])^(a[59] & b[339])^(a[58] & b[340])^(a[57] & b[341])^(a[56] & b[342])^(a[55] & b[343])^(a[54] & b[344])^(a[53] & b[345])^(a[52] & b[346])^(a[51] & b[347])^(a[50] & b[348])^(a[49] & b[349])^(a[48] & b[350])^(a[47] & b[351])^(a[46] & b[352])^(a[45] & b[353])^(a[44] & b[354])^(a[43] & b[355])^(a[42] & b[356])^(a[41] & b[357])^(a[40] & b[358])^(a[39] & b[359])^(a[38] & b[360])^(a[37] & b[361])^(a[36] & b[362])^(a[35] & b[363])^(a[34] & b[364])^(a[33] & b[365])^(a[32] & b[366])^(a[31] & b[367])^(a[30] & b[368])^(a[29] & b[369])^(a[28] & b[370])^(a[27] & b[371])^(a[26] & b[372])^(a[25] & b[373])^(a[24] & b[374])^(a[23] & b[375])^(a[22] & b[376])^(a[21] & b[377])^(a[20] & b[378])^(a[19] & b[379])^(a[18] & b[380])^(a[17] & b[381])^(a[16] & b[382])^(a[15] & b[383])^(a[14] & b[384])^(a[13] & b[385])^(a[12] & b[386])^(a[11] & b[387])^(a[10] & b[388])^(a[9] & b[389])^(a[8] & b[390])^(a[7] & b[391])^(a[6] & b[392])^(a[5] & b[393])^(a[4] & b[394])^(a[3] & b[395])^(a[2] & b[396])^(a[1] & b[397])^(a[0] & b[398]);
assign y[399] = (a[399] & b[0])^(a[398] & b[1])^(a[397] & b[2])^(a[396] & b[3])^(a[395] & b[4])^(a[394] & b[5])^(a[393] & b[6])^(a[392] & b[7])^(a[391] & b[8])^(a[390] & b[9])^(a[389] & b[10])^(a[388] & b[11])^(a[387] & b[12])^(a[386] & b[13])^(a[385] & b[14])^(a[384] & b[15])^(a[383] & b[16])^(a[382] & b[17])^(a[381] & b[18])^(a[380] & b[19])^(a[379] & b[20])^(a[378] & b[21])^(a[377] & b[22])^(a[376] & b[23])^(a[375] & b[24])^(a[374] & b[25])^(a[373] & b[26])^(a[372] & b[27])^(a[371] & b[28])^(a[370] & b[29])^(a[369] & b[30])^(a[368] & b[31])^(a[367] & b[32])^(a[366] & b[33])^(a[365] & b[34])^(a[364] & b[35])^(a[363] & b[36])^(a[362] & b[37])^(a[361] & b[38])^(a[360] & b[39])^(a[359] & b[40])^(a[358] & b[41])^(a[357] & b[42])^(a[356] & b[43])^(a[355] & b[44])^(a[354] & b[45])^(a[353] & b[46])^(a[352] & b[47])^(a[351] & b[48])^(a[350] & b[49])^(a[349] & b[50])^(a[348] & b[51])^(a[347] & b[52])^(a[346] & b[53])^(a[345] & b[54])^(a[344] & b[55])^(a[343] & b[56])^(a[342] & b[57])^(a[341] & b[58])^(a[340] & b[59])^(a[339] & b[60])^(a[338] & b[61])^(a[337] & b[62])^(a[336] & b[63])^(a[335] & b[64])^(a[334] & b[65])^(a[333] & b[66])^(a[332] & b[67])^(a[331] & b[68])^(a[330] & b[69])^(a[329] & b[70])^(a[328] & b[71])^(a[327] & b[72])^(a[326] & b[73])^(a[325] & b[74])^(a[324] & b[75])^(a[323] & b[76])^(a[322] & b[77])^(a[321] & b[78])^(a[320] & b[79])^(a[319] & b[80])^(a[318] & b[81])^(a[317] & b[82])^(a[316] & b[83])^(a[315] & b[84])^(a[314] & b[85])^(a[313] & b[86])^(a[312] & b[87])^(a[311] & b[88])^(a[310] & b[89])^(a[309] & b[90])^(a[308] & b[91])^(a[307] & b[92])^(a[306] & b[93])^(a[305] & b[94])^(a[304] & b[95])^(a[303] & b[96])^(a[302] & b[97])^(a[301] & b[98])^(a[300] & b[99])^(a[299] & b[100])^(a[298] & b[101])^(a[297] & b[102])^(a[296] & b[103])^(a[295] & b[104])^(a[294] & b[105])^(a[293] & b[106])^(a[292] & b[107])^(a[291] & b[108])^(a[290] & b[109])^(a[289] & b[110])^(a[288] & b[111])^(a[287] & b[112])^(a[286] & b[113])^(a[285] & b[114])^(a[284] & b[115])^(a[283] & b[116])^(a[282] & b[117])^(a[281] & b[118])^(a[280] & b[119])^(a[279] & b[120])^(a[278] & b[121])^(a[277] & b[122])^(a[276] & b[123])^(a[275] & b[124])^(a[274] & b[125])^(a[273] & b[126])^(a[272] & b[127])^(a[271] & b[128])^(a[270] & b[129])^(a[269] & b[130])^(a[268] & b[131])^(a[267] & b[132])^(a[266] & b[133])^(a[265] & b[134])^(a[264] & b[135])^(a[263] & b[136])^(a[262] & b[137])^(a[261] & b[138])^(a[260] & b[139])^(a[259] & b[140])^(a[258] & b[141])^(a[257] & b[142])^(a[256] & b[143])^(a[255] & b[144])^(a[254] & b[145])^(a[253] & b[146])^(a[252] & b[147])^(a[251] & b[148])^(a[250] & b[149])^(a[249] & b[150])^(a[248] & b[151])^(a[247] & b[152])^(a[246] & b[153])^(a[245] & b[154])^(a[244] & b[155])^(a[243] & b[156])^(a[242] & b[157])^(a[241] & b[158])^(a[240] & b[159])^(a[239] & b[160])^(a[238] & b[161])^(a[237] & b[162])^(a[236] & b[163])^(a[235] & b[164])^(a[234] & b[165])^(a[233] & b[166])^(a[232] & b[167])^(a[231] & b[168])^(a[230] & b[169])^(a[229] & b[170])^(a[228] & b[171])^(a[227] & b[172])^(a[226] & b[173])^(a[225] & b[174])^(a[224] & b[175])^(a[223] & b[176])^(a[222] & b[177])^(a[221] & b[178])^(a[220] & b[179])^(a[219] & b[180])^(a[218] & b[181])^(a[217] & b[182])^(a[216] & b[183])^(a[215] & b[184])^(a[214] & b[185])^(a[213] & b[186])^(a[212] & b[187])^(a[211] & b[188])^(a[210] & b[189])^(a[209] & b[190])^(a[208] & b[191])^(a[207] & b[192])^(a[206] & b[193])^(a[205] & b[194])^(a[204] & b[195])^(a[203] & b[196])^(a[202] & b[197])^(a[201] & b[198])^(a[200] & b[199])^(a[199] & b[200])^(a[198] & b[201])^(a[197] & b[202])^(a[196] & b[203])^(a[195] & b[204])^(a[194] & b[205])^(a[193] & b[206])^(a[192] & b[207])^(a[191] & b[208])^(a[190] & b[209])^(a[189] & b[210])^(a[188] & b[211])^(a[187] & b[212])^(a[186] & b[213])^(a[185] & b[214])^(a[184] & b[215])^(a[183] & b[216])^(a[182] & b[217])^(a[181] & b[218])^(a[180] & b[219])^(a[179] & b[220])^(a[178] & b[221])^(a[177] & b[222])^(a[176] & b[223])^(a[175] & b[224])^(a[174] & b[225])^(a[173] & b[226])^(a[172] & b[227])^(a[171] & b[228])^(a[170] & b[229])^(a[169] & b[230])^(a[168] & b[231])^(a[167] & b[232])^(a[166] & b[233])^(a[165] & b[234])^(a[164] & b[235])^(a[163] & b[236])^(a[162] & b[237])^(a[161] & b[238])^(a[160] & b[239])^(a[159] & b[240])^(a[158] & b[241])^(a[157] & b[242])^(a[156] & b[243])^(a[155] & b[244])^(a[154] & b[245])^(a[153] & b[246])^(a[152] & b[247])^(a[151] & b[248])^(a[150] & b[249])^(a[149] & b[250])^(a[148] & b[251])^(a[147] & b[252])^(a[146] & b[253])^(a[145] & b[254])^(a[144] & b[255])^(a[143] & b[256])^(a[142] & b[257])^(a[141] & b[258])^(a[140] & b[259])^(a[139] & b[260])^(a[138] & b[261])^(a[137] & b[262])^(a[136] & b[263])^(a[135] & b[264])^(a[134] & b[265])^(a[133] & b[266])^(a[132] & b[267])^(a[131] & b[268])^(a[130] & b[269])^(a[129] & b[270])^(a[128] & b[271])^(a[127] & b[272])^(a[126] & b[273])^(a[125] & b[274])^(a[124] & b[275])^(a[123] & b[276])^(a[122] & b[277])^(a[121] & b[278])^(a[120] & b[279])^(a[119] & b[280])^(a[118] & b[281])^(a[117] & b[282])^(a[116] & b[283])^(a[115] & b[284])^(a[114] & b[285])^(a[113] & b[286])^(a[112] & b[287])^(a[111] & b[288])^(a[110] & b[289])^(a[109] & b[290])^(a[108] & b[291])^(a[107] & b[292])^(a[106] & b[293])^(a[105] & b[294])^(a[104] & b[295])^(a[103] & b[296])^(a[102] & b[297])^(a[101] & b[298])^(a[100] & b[299])^(a[99] & b[300])^(a[98] & b[301])^(a[97] & b[302])^(a[96] & b[303])^(a[95] & b[304])^(a[94] & b[305])^(a[93] & b[306])^(a[92] & b[307])^(a[91] & b[308])^(a[90] & b[309])^(a[89] & b[310])^(a[88] & b[311])^(a[87] & b[312])^(a[86] & b[313])^(a[85] & b[314])^(a[84] & b[315])^(a[83] & b[316])^(a[82] & b[317])^(a[81] & b[318])^(a[80] & b[319])^(a[79] & b[320])^(a[78] & b[321])^(a[77] & b[322])^(a[76] & b[323])^(a[75] & b[324])^(a[74] & b[325])^(a[73] & b[326])^(a[72] & b[327])^(a[71] & b[328])^(a[70] & b[329])^(a[69] & b[330])^(a[68] & b[331])^(a[67] & b[332])^(a[66] & b[333])^(a[65] & b[334])^(a[64] & b[335])^(a[63] & b[336])^(a[62] & b[337])^(a[61] & b[338])^(a[60] & b[339])^(a[59] & b[340])^(a[58] & b[341])^(a[57] & b[342])^(a[56] & b[343])^(a[55] & b[344])^(a[54] & b[345])^(a[53] & b[346])^(a[52] & b[347])^(a[51] & b[348])^(a[50] & b[349])^(a[49] & b[350])^(a[48] & b[351])^(a[47] & b[352])^(a[46] & b[353])^(a[45] & b[354])^(a[44] & b[355])^(a[43] & b[356])^(a[42] & b[357])^(a[41] & b[358])^(a[40] & b[359])^(a[39] & b[360])^(a[38] & b[361])^(a[37] & b[362])^(a[36] & b[363])^(a[35] & b[364])^(a[34] & b[365])^(a[33] & b[366])^(a[32] & b[367])^(a[31] & b[368])^(a[30] & b[369])^(a[29] & b[370])^(a[28] & b[371])^(a[27] & b[372])^(a[26] & b[373])^(a[25] & b[374])^(a[24] & b[375])^(a[23] & b[376])^(a[22] & b[377])^(a[21] & b[378])^(a[20] & b[379])^(a[19] & b[380])^(a[18] & b[381])^(a[17] & b[382])^(a[16] & b[383])^(a[15] & b[384])^(a[14] & b[385])^(a[13] & b[386])^(a[12] & b[387])^(a[11] & b[388])^(a[10] & b[389])^(a[9] & b[390])^(a[8] & b[391])^(a[7] & b[392])^(a[6] & b[393])^(a[5] & b[394])^(a[4] & b[395])^(a[3] & b[396])^(a[2] & b[397])^(a[1] & b[398])^(a[0] & b[399]);
assign y[400] = (a[400] & b[0])^(a[399] & b[1])^(a[398] & b[2])^(a[397] & b[3])^(a[396] & b[4])^(a[395] & b[5])^(a[394] & b[6])^(a[393] & b[7])^(a[392] & b[8])^(a[391] & b[9])^(a[390] & b[10])^(a[389] & b[11])^(a[388] & b[12])^(a[387] & b[13])^(a[386] & b[14])^(a[385] & b[15])^(a[384] & b[16])^(a[383] & b[17])^(a[382] & b[18])^(a[381] & b[19])^(a[380] & b[20])^(a[379] & b[21])^(a[378] & b[22])^(a[377] & b[23])^(a[376] & b[24])^(a[375] & b[25])^(a[374] & b[26])^(a[373] & b[27])^(a[372] & b[28])^(a[371] & b[29])^(a[370] & b[30])^(a[369] & b[31])^(a[368] & b[32])^(a[367] & b[33])^(a[366] & b[34])^(a[365] & b[35])^(a[364] & b[36])^(a[363] & b[37])^(a[362] & b[38])^(a[361] & b[39])^(a[360] & b[40])^(a[359] & b[41])^(a[358] & b[42])^(a[357] & b[43])^(a[356] & b[44])^(a[355] & b[45])^(a[354] & b[46])^(a[353] & b[47])^(a[352] & b[48])^(a[351] & b[49])^(a[350] & b[50])^(a[349] & b[51])^(a[348] & b[52])^(a[347] & b[53])^(a[346] & b[54])^(a[345] & b[55])^(a[344] & b[56])^(a[343] & b[57])^(a[342] & b[58])^(a[341] & b[59])^(a[340] & b[60])^(a[339] & b[61])^(a[338] & b[62])^(a[337] & b[63])^(a[336] & b[64])^(a[335] & b[65])^(a[334] & b[66])^(a[333] & b[67])^(a[332] & b[68])^(a[331] & b[69])^(a[330] & b[70])^(a[329] & b[71])^(a[328] & b[72])^(a[327] & b[73])^(a[326] & b[74])^(a[325] & b[75])^(a[324] & b[76])^(a[323] & b[77])^(a[322] & b[78])^(a[321] & b[79])^(a[320] & b[80])^(a[319] & b[81])^(a[318] & b[82])^(a[317] & b[83])^(a[316] & b[84])^(a[315] & b[85])^(a[314] & b[86])^(a[313] & b[87])^(a[312] & b[88])^(a[311] & b[89])^(a[310] & b[90])^(a[309] & b[91])^(a[308] & b[92])^(a[307] & b[93])^(a[306] & b[94])^(a[305] & b[95])^(a[304] & b[96])^(a[303] & b[97])^(a[302] & b[98])^(a[301] & b[99])^(a[300] & b[100])^(a[299] & b[101])^(a[298] & b[102])^(a[297] & b[103])^(a[296] & b[104])^(a[295] & b[105])^(a[294] & b[106])^(a[293] & b[107])^(a[292] & b[108])^(a[291] & b[109])^(a[290] & b[110])^(a[289] & b[111])^(a[288] & b[112])^(a[287] & b[113])^(a[286] & b[114])^(a[285] & b[115])^(a[284] & b[116])^(a[283] & b[117])^(a[282] & b[118])^(a[281] & b[119])^(a[280] & b[120])^(a[279] & b[121])^(a[278] & b[122])^(a[277] & b[123])^(a[276] & b[124])^(a[275] & b[125])^(a[274] & b[126])^(a[273] & b[127])^(a[272] & b[128])^(a[271] & b[129])^(a[270] & b[130])^(a[269] & b[131])^(a[268] & b[132])^(a[267] & b[133])^(a[266] & b[134])^(a[265] & b[135])^(a[264] & b[136])^(a[263] & b[137])^(a[262] & b[138])^(a[261] & b[139])^(a[260] & b[140])^(a[259] & b[141])^(a[258] & b[142])^(a[257] & b[143])^(a[256] & b[144])^(a[255] & b[145])^(a[254] & b[146])^(a[253] & b[147])^(a[252] & b[148])^(a[251] & b[149])^(a[250] & b[150])^(a[249] & b[151])^(a[248] & b[152])^(a[247] & b[153])^(a[246] & b[154])^(a[245] & b[155])^(a[244] & b[156])^(a[243] & b[157])^(a[242] & b[158])^(a[241] & b[159])^(a[240] & b[160])^(a[239] & b[161])^(a[238] & b[162])^(a[237] & b[163])^(a[236] & b[164])^(a[235] & b[165])^(a[234] & b[166])^(a[233] & b[167])^(a[232] & b[168])^(a[231] & b[169])^(a[230] & b[170])^(a[229] & b[171])^(a[228] & b[172])^(a[227] & b[173])^(a[226] & b[174])^(a[225] & b[175])^(a[224] & b[176])^(a[223] & b[177])^(a[222] & b[178])^(a[221] & b[179])^(a[220] & b[180])^(a[219] & b[181])^(a[218] & b[182])^(a[217] & b[183])^(a[216] & b[184])^(a[215] & b[185])^(a[214] & b[186])^(a[213] & b[187])^(a[212] & b[188])^(a[211] & b[189])^(a[210] & b[190])^(a[209] & b[191])^(a[208] & b[192])^(a[207] & b[193])^(a[206] & b[194])^(a[205] & b[195])^(a[204] & b[196])^(a[203] & b[197])^(a[202] & b[198])^(a[201] & b[199])^(a[200] & b[200])^(a[199] & b[201])^(a[198] & b[202])^(a[197] & b[203])^(a[196] & b[204])^(a[195] & b[205])^(a[194] & b[206])^(a[193] & b[207])^(a[192] & b[208])^(a[191] & b[209])^(a[190] & b[210])^(a[189] & b[211])^(a[188] & b[212])^(a[187] & b[213])^(a[186] & b[214])^(a[185] & b[215])^(a[184] & b[216])^(a[183] & b[217])^(a[182] & b[218])^(a[181] & b[219])^(a[180] & b[220])^(a[179] & b[221])^(a[178] & b[222])^(a[177] & b[223])^(a[176] & b[224])^(a[175] & b[225])^(a[174] & b[226])^(a[173] & b[227])^(a[172] & b[228])^(a[171] & b[229])^(a[170] & b[230])^(a[169] & b[231])^(a[168] & b[232])^(a[167] & b[233])^(a[166] & b[234])^(a[165] & b[235])^(a[164] & b[236])^(a[163] & b[237])^(a[162] & b[238])^(a[161] & b[239])^(a[160] & b[240])^(a[159] & b[241])^(a[158] & b[242])^(a[157] & b[243])^(a[156] & b[244])^(a[155] & b[245])^(a[154] & b[246])^(a[153] & b[247])^(a[152] & b[248])^(a[151] & b[249])^(a[150] & b[250])^(a[149] & b[251])^(a[148] & b[252])^(a[147] & b[253])^(a[146] & b[254])^(a[145] & b[255])^(a[144] & b[256])^(a[143] & b[257])^(a[142] & b[258])^(a[141] & b[259])^(a[140] & b[260])^(a[139] & b[261])^(a[138] & b[262])^(a[137] & b[263])^(a[136] & b[264])^(a[135] & b[265])^(a[134] & b[266])^(a[133] & b[267])^(a[132] & b[268])^(a[131] & b[269])^(a[130] & b[270])^(a[129] & b[271])^(a[128] & b[272])^(a[127] & b[273])^(a[126] & b[274])^(a[125] & b[275])^(a[124] & b[276])^(a[123] & b[277])^(a[122] & b[278])^(a[121] & b[279])^(a[120] & b[280])^(a[119] & b[281])^(a[118] & b[282])^(a[117] & b[283])^(a[116] & b[284])^(a[115] & b[285])^(a[114] & b[286])^(a[113] & b[287])^(a[112] & b[288])^(a[111] & b[289])^(a[110] & b[290])^(a[109] & b[291])^(a[108] & b[292])^(a[107] & b[293])^(a[106] & b[294])^(a[105] & b[295])^(a[104] & b[296])^(a[103] & b[297])^(a[102] & b[298])^(a[101] & b[299])^(a[100] & b[300])^(a[99] & b[301])^(a[98] & b[302])^(a[97] & b[303])^(a[96] & b[304])^(a[95] & b[305])^(a[94] & b[306])^(a[93] & b[307])^(a[92] & b[308])^(a[91] & b[309])^(a[90] & b[310])^(a[89] & b[311])^(a[88] & b[312])^(a[87] & b[313])^(a[86] & b[314])^(a[85] & b[315])^(a[84] & b[316])^(a[83] & b[317])^(a[82] & b[318])^(a[81] & b[319])^(a[80] & b[320])^(a[79] & b[321])^(a[78] & b[322])^(a[77] & b[323])^(a[76] & b[324])^(a[75] & b[325])^(a[74] & b[326])^(a[73] & b[327])^(a[72] & b[328])^(a[71] & b[329])^(a[70] & b[330])^(a[69] & b[331])^(a[68] & b[332])^(a[67] & b[333])^(a[66] & b[334])^(a[65] & b[335])^(a[64] & b[336])^(a[63] & b[337])^(a[62] & b[338])^(a[61] & b[339])^(a[60] & b[340])^(a[59] & b[341])^(a[58] & b[342])^(a[57] & b[343])^(a[56] & b[344])^(a[55] & b[345])^(a[54] & b[346])^(a[53] & b[347])^(a[52] & b[348])^(a[51] & b[349])^(a[50] & b[350])^(a[49] & b[351])^(a[48] & b[352])^(a[47] & b[353])^(a[46] & b[354])^(a[45] & b[355])^(a[44] & b[356])^(a[43] & b[357])^(a[42] & b[358])^(a[41] & b[359])^(a[40] & b[360])^(a[39] & b[361])^(a[38] & b[362])^(a[37] & b[363])^(a[36] & b[364])^(a[35] & b[365])^(a[34] & b[366])^(a[33] & b[367])^(a[32] & b[368])^(a[31] & b[369])^(a[30] & b[370])^(a[29] & b[371])^(a[28] & b[372])^(a[27] & b[373])^(a[26] & b[374])^(a[25] & b[375])^(a[24] & b[376])^(a[23] & b[377])^(a[22] & b[378])^(a[21] & b[379])^(a[20] & b[380])^(a[19] & b[381])^(a[18] & b[382])^(a[17] & b[383])^(a[16] & b[384])^(a[15] & b[385])^(a[14] & b[386])^(a[13] & b[387])^(a[12] & b[388])^(a[11] & b[389])^(a[10] & b[390])^(a[9] & b[391])^(a[8] & b[392])^(a[7] & b[393])^(a[6] & b[394])^(a[5] & b[395])^(a[4] & b[396])^(a[3] & b[397])^(a[2] & b[398])^(a[1] & b[399])^(a[0] & b[400]);
assign y[401] = (a[401] & b[0])^(a[400] & b[1])^(a[399] & b[2])^(a[398] & b[3])^(a[397] & b[4])^(a[396] & b[5])^(a[395] & b[6])^(a[394] & b[7])^(a[393] & b[8])^(a[392] & b[9])^(a[391] & b[10])^(a[390] & b[11])^(a[389] & b[12])^(a[388] & b[13])^(a[387] & b[14])^(a[386] & b[15])^(a[385] & b[16])^(a[384] & b[17])^(a[383] & b[18])^(a[382] & b[19])^(a[381] & b[20])^(a[380] & b[21])^(a[379] & b[22])^(a[378] & b[23])^(a[377] & b[24])^(a[376] & b[25])^(a[375] & b[26])^(a[374] & b[27])^(a[373] & b[28])^(a[372] & b[29])^(a[371] & b[30])^(a[370] & b[31])^(a[369] & b[32])^(a[368] & b[33])^(a[367] & b[34])^(a[366] & b[35])^(a[365] & b[36])^(a[364] & b[37])^(a[363] & b[38])^(a[362] & b[39])^(a[361] & b[40])^(a[360] & b[41])^(a[359] & b[42])^(a[358] & b[43])^(a[357] & b[44])^(a[356] & b[45])^(a[355] & b[46])^(a[354] & b[47])^(a[353] & b[48])^(a[352] & b[49])^(a[351] & b[50])^(a[350] & b[51])^(a[349] & b[52])^(a[348] & b[53])^(a[347] & b[54])^(a[346] & b[55])^(a[345] & b[56])^(a[344] & b[57])^(a[343] & b[58])^(a[342] & b[59])^(a[341] & b[60])^(a[340] & b[61])^(a[339] & b[62])^(a[338] & b[63])^(a[337] & b[64])^(a[336] & b[65])^(a[335] & b[66])^(a[334] & b[67])^(a[333] & b[68])^(a[332] & b[69])^(a[331] & b[70])^(a[330] & b[71])^(a[329] & b[72])^(a[328] & b[73])^(a[327] & b[74])^(a[326] & b[75])^(a[325] & b[76])^(a[324] & b[77])^(a[323] & b[78])^(a[322] & b[79])^(a[321] & b[80])^(a[320] & b[81])^(a[319] & b[82])^(a[318] & b[83])^(a[317] & b[84])^(a[316] & b[85])^(a[315] & b[86])^(a[314] & b[87])^(a[313] & b[88])^(a[312] & b[89])^(a[311] & b[90])^(a[310] & b[91])^(a[309] & b[92])^(a[308] & b[93])^(a[307] & b[94])^(a[306] & b[95])^(a[305] & b[96])^(a[304] & b[97])^(a[303] & b[98])^(a[302] & b[99])^(a[301] & b[100])^(a[300] & b[101])^(a[299] & b[102])^(a[298] & b[103])^(a[297] & b[104])^(a[296] & b[105])^(a[295] & b[106])^(a[294] & b[107])^(a[293] & b[108])^(a[292] & b[109])^(a[291] & b[110])^(a[290] & b[111])^(a[289] & b[112])^(a[288] & b[113])^(a[287] & b[114])^(a[286] & b[115])^(a[285] & b[116])^(a[284] & b[117])^(a[283] & b[118])^(a[282] & b[119])^(a[281] & b[120])^(a[280] & b[121])^(a[279] & b[122])^(a[278] & b[123])^(a[277] & b[124])^(a[276] & b[125])^(a[275] & b[126])^(a[274] & b[127])^(a[273] & b[128])^(a[272] & b[129])^(a[271] & b[130])^(a[270] & b[131])^(a[269] & b[132])^(a[268] & b[133])^(a[267] & b[134])^(a[266] & b[135])^(a[265] & b[136])^(a[264] & b[137])^(a[263] & b[138])^(a[262] & b[139])^(a[261] & b[140])^(a[260] & b[141])^(a[259] & b[142])^(a[258] & b[143])^(a[257] & b[144])^(a[256] & b[145])^(a[255] & b[146])^(a[254] & b[147])^(a[253] & b[148])^(a[252] & b[149])^(a[251] & b[150])^(a[250] & b[151])^(a[249] & b[152])^(a[248] & b[153])^(a[247] & b[154])^(a[246] & b[155])^(a[245] & b[156])^(a[244] & b[157])^(a[243] & b[158])^(a[242] & b[159])^(a[241] & b[160])^(a[240] & b[161])^(a[239] & b[162])^(a[238] & b[163])^(a[237] & b[164])^(a[236] & b[165])^(a[235] & b[166])^(a[234] & b[167])^(a[233] & b[168])^(a[232] & b[169])^(a[231] & b[170])^(a[230] & b[171])^(a[229] & b[172])^(a[228] & b[173])^(a[227] & b[174])^(a[226] & b[175])^(a[225] & b[176])^(a[224] & b[177])^(a[223] & b[178])^(a[222] & b[179])^(a[221] & b[180])^(a[220] & b[181])^(a[219] & b[182])^(a[218] & b[183])^(a[217] & b[184])^(a[216] & b[185])^(a[215] & b[186])^(a[214] & b[187])^(a[213] & b[188])^(a[212] & b[189])^(a[211] & b[190])^(a[210] & b[191])^(a[209] & b[192])^(a[208] & b[193])^(a[207] & b[194])^(a[206] & b[195])^(a[205] & b[196])^(a[204] & b[197])^(a[203] & b[198])^(a[202] & b[199])^(a[201] & b[200])^(a[200] & b[201])^(a[199] & b[202])^(a[198] & b[203])^(a[197] & b[204])^(a[196] & b[205])^(a[195] & b[206])^(a[194] & b[207])^(a[193] & b[208])^(a[192] & b[209])^(a[191] & b[210])^(a[190] & b[211])^(a[189] & b[212])^(a[188] & b[213])^(a[187] & b[214])^(a[186] & b[215])^(a[185] & b[216])^(a[184] & b[217])^(a[183] & b[218])^(a[182] & b[219])^(a[181] & b[220])^(a[180] & b[221])^(a[179] & b[222])^(a[178] & b[223])^(a[177] & b[224])^(a[176] & b[225])^(a[175] & b[226])^(a[174] & b[227])^(a[173] & b[228])^(a[172] & b[229])^(a[171] & b[230])^(a[170] & b[231])^(a[169] & b[232])^(a[168] & b[233])^(a[167] & b[234])^(a[166] & b[235])^(a[165] & b[236])^(a[164] & b[237])^(a[163] & b[238])^(a[162] & b[239])^(a[161] & b[240])^(a[160] & b[241])^(a[159] & b[242])^(a[158] & b[243])^(a[157] & b[244])^(a[156] & b[245])^(a[155] & b[246])^(a[154] & b[247])^(a[153] & b[248])^(a[152] & b[249])^(a[151] & b[250])^(a[150] & b[251])^(a[149] & b[252])^(a[148] & b[253])^(a[147] & b[254])^(a[146] & b[255])^(a[145] & b[256])^(a[144] & b[257])^(a[143] & b[258])^(a[142] & b[259])^(a[141] & b[260])^(a[140] & b[261])^(a[139] & b[262])^(a[138] & b[263])^(a[137] & b[264])^(a[136] & b[265])^(a[135] & b[266])^(a[134] & b[267])^(a[133] & b[268])^(a[132] & b[269])^(a[131] & b[270])^(a[130] & b[271])^(a[129] & b[272])^(a[128] & b[273])^(a[127] & b[274])^(a[126] & b[275])^(a[125] & b[276])^(a[124] & b[277])^(a[123] & b[278])^(a[122] & b[279])^(a[121] & b[280])^(a[120] & b[281])^(a[119] & b[282])^(a[118] & b[283])^(a[117] & b[284])^(a[116] & b[285])^(a[115] & b[286])^(a[114] & b[287])^(a[113] & b[288])^(a[112] & b[289])^(a[111] & b[290])^(a[110] & b[291])^(a[109] & b[292])^(a[108] & b[293])^(a[107] & b[294])^(a[106] & b[295])^(a[105] & b[296])^(a[104] & b[297])^(a[103] & b[298])^(a[102] & b[299])^(a[101] & b[300])^(a[100] & b[301])^(a[99] & b[302])^(a[98] & b[303])^(a[97] & b[304])^(a[96] & b[305])^(a[95] & b[306])^(a[94] & b[307])^(a[93] & b[308])^(a[92] & b[309])^(a[91] & b[310])^(a[90] & b[311])^(a[89] & b[312])^(a[88] & b[313])^(a[87] & b[314])^(a[86] & b[315])^(a[85] & b[316])^(a[84] & b[317])^(a[83] & b[318])^(a[82] & b[319])^(a[81] & b[320])^(a[80] & b[321])^(a[79] & b[322])^(a[78] & b[323])^(a[77] & b[324])^(a[76] & b[325])^(a[75] & b[326])^(a[74] & b[327])^(a[73] & b[328])^(a[72] & b[329])^(a[71] & b[330])^(a[70] & b[331])^(a[69] & b[332])^(a[68] & b[333])^(a[67] & b[334])^(a[66] & b[335])^(a[65] & b[336])^(a[64] & b[337])^(a[63] & b[338])^(a[62] & b[339])^(a[61] & b[340])^(a[60] & b[341])^(a[59] & b[342])^(a[58] & b[343])^(a[57] & b[344])^(a[56] & b[345])^(a[55] & b[346])^(a[54] & b[347])^(a[53] & b[348])^(a[52] & b[349])^(a[51] & b[350])^(a[50] & b[351])^(a[49] & b[352])^(a[48] & b[353])^(a[47] & b[354])^(a[46] & b[355])^(a[45] & b[356])^(a[44] & b[357])^(a[43] & b[358])^(a[42] & b[359])^(a[41] & b[360])^(a[40] & b[361])^(a[39] & b[362])^(a[38] & b[363])^(a[37] & b[364])^(a[36] & b[365])^(a[35] & b[366])^(a[34] & b[367])^(a[33] & b[368])^(a[32] & b[369])^(a[31] & b[370])^(a[30] & b[371])^(a[29] & b[372])^(a[28] & b[373])^(a[27] & b[374])^(a[26] & b[375])^(a[25] & b[376])^(a[24] & b[377])^(a[23] & b[378])^(a[22] & b[379])^(a[21] & b[380])^(a[20] & b[381])^(a[19] & b[382])^(a[18] & b[383])^(a[17] & b[384])^(a[16] & b[385])^(a[15] & b[386])^(a[14] & b[387])^(a[13] & b[388])^(a[12] & b[389])^(a[11] & b[390])^(a[10] & b[391])^(a[9] & b[392])^(a[8] & b[393])^(a[7] & b[394])^(a[6] & b[395])^(a[5] & b[396])^(a[4] & b[397])^(a[3] & b[398])^(a[2] & b[399])^(a[1] & b[400])^(a[0] & b[401]);
assign y[402] = (a[402] & b[0])^(a[401] & b[1])^(a[400] & b[2])^(a[399] & b[3])^(a[398] & b[4])^(a[397] & b[5])^(a[396] & b[6])^(a[395] & b[7])^(a[394] & b[8])^(a[393] & b[9])^(a[392] & b[10])^(a[391] & b[11])^(a[390] & b[12])^(a[389] & b[13])^(a[388] & b[14])^(a[387] & b[15])^(a[386] & b[16])^(a[385] & b[17])^(a[384] & b[18])^(a[383] & b[19])^(a[382] & b[20])^(a[381] & b[21])^(a[380] & b[22])^(a[379] & b[23])^(a[378] & b[24])^(a[377] & b[25])^(a[376] & b[26])^(a[375] & b[27])^(a[374] & b[28])^(a[373] & b[29])^(a[372] & b[30])^(a[371] & b[31])^(a[370] & b[32])^(a[369] & b[33])^(a[368] & b[34])^(a[367] & b[35])^(a[366] & b[36])^(a[365] & b[37])^(a[364] & b[38])^(a[363] & b[39])^(a[362] & b[40])^(a[361] & b[41])^(a[360] & b[42])^(a[359] & b[43])^(a[358] & b[44])^(a[357] & b[45])^(a[356] & b[46])^(a[355] & b[47])^(a[354] & b[48])^(a[353] & b[49])^(a[352] & b[50])^(a[351] & b[51])^(a[350] & b[52])^(a[349] & b[53])^(a[348] & b[54])^(a[347] & b[55])^(a[346] & b[56])^(a[345] & b[57])^(a[344] & b[58])^(a[343] & b[59])^(a[342] & b[60])^(a[341] & b[61])^(a[340] & b[62])^(a[339] & b[63])^(a[338] & b[64])^(a[337] & b[65])^(a[336] & b[66])^(a[335] & b[67])^(a[334] & b[68])^(a[333] & b[69])^(a[332] & b[70])^(a[331] & b[71])^(a[330] & b[72])^(a[329] & b[73])^(a[328] & b[74])^(a[327] & b[75])^(a[326] & b[76])^(a[325] & b[77])^(a[324] & b[78])^(a[323] & b[79])^(a[322] & b[80])^(a[321] & b[81])^(a[320] & b[82])^(a[319] & b[83])^(a[318] & b[84])^(a[317] & b[85])^(a[316] & b[86])^(a[315] & b[87])^(a[314] & b[88])^(a[313] & b[89])^(a[312] & b[90])^(a[311] & b[91])^(a[310] & b[92])^(a[309] & b[93])^(a[308] & b[94])^(a[307] & b[95])^(a[306] & b[96])^(a[305] & b[97])^(a[304] & b[98])^(a[303] & b[99])^(a[302] & b[100])^(a[301] & b[101])^(a[300] & b[102])^(a[299] & b[103])^(a[298] & b[104])^(a[297] & b[105])^(a[296] & b[106])^(a[295] & b[107])^(a[294] & b[108])^(a[293] & b[109])^(a[292] & b[110])^(a[291] & b[111])^(a[290] & b[112])^(a[289] & b[113])^(a[288] & b[114])^(a[287] & b[115])^(a[286] & b[116])^(a[285] & b[117])^(a[284] & b[118])^(a[283] & b[119])^(a[282] & b[120])^(a[281] & b[121])^(a[280] & b[122])^(a[279] & b[123])^(a[278] & b[124])^(a[277] & b[125])^(a[276] & b[126])^(a[275] & b[127])^(a[274] & b[128])^(a[273] & b[129])^(a[272] & b[130])^(a[271] & b[131])^(a[270] & b[132])^(a[269] & b[133])^(a[268] & b[134])^(a[267] & b[135])^(a[266] & b[136])^(a[265] & b[137])^(a[264] & b[138])^(a[263] & b[139])^(a[262] & b[140])^(a[261] & b[141])^(a[260] & b[142])^(a[259] & b[143])^(a[258] & b[144])^(a[257] & b[145])^(a[256] & b[146])^(a[255] & b[147])^(a[254] & b[148])^(a[253] & b[149])^(a[252] & b[150])^(a[251] & b[151])^(a[250] & b[152])^(a[249] & b[153])^(a[248] & b[154])^(a[247] & b[155])^(a[246] & b[156])^(a[245] & b[157])^(a[244] & b[158])^(a[243] & b[159])^(a[242] & b[160])^(a[241] & b[161])^(a[240] & b[162])^(a[239] & b[163])^(a[238] & b[164])^(a[237] & b[165])^(a[236] & b[166])^(a[235] & b[167])^(a[234] & b[168])^(a[233] & b[169])^(a[232] & b[170])^(a[231] & b[171])^(a[230] & b[172])^(a[229] & b[173])^(a[228] & b[174])^(a[227] & b[175])^(a[226] & b[176])^(a[225] & b[177])^(a[224] & b[178])^(a[223] & b[179])^(a[222] & b[180])^(a[221] & b[181])^(a[220] & b[182])^(a[219] & b[183])^(a[218] & b[184])^(a[217] & b[185])^(a[216] & b[186])^(a[215] & b[187])^(a[214] & b[188])^(a[213] & b[189])^(a[212] & b[190])^(a[211] & b[191])^(a[210] & b[192])^(a[209] & b[193])^(a[208] & b[194])^(a[207] & b[195])^(a[206] & b[196])^(a[205] & b[197])^(a[204] & b[198])^(a[203] & b[199])^(a[202] & b[200])^(a[201] & b[201])^(a[200] & b[202])^(a[199] & b[203])^(a[198] & b[204])^(a[197] & b[205])^(a[196] & b[206])^(a[195] & b[207])^(a[194] & b[208])^(a[193] & b[209])^(a[192] & b[210])^(a[191] & b[211])^(a[190] & b[212])^(a[189] & b[213])^(a[188] & b[214])^(a[187] & b[215])^(a[186] & b[216])^(a[185] & b[217])^(a[184] & b[218])^(a[183] & b[219])^(a[182] & b[220])^(a[181] & b[221])^(a[180] & b[222])^(a[179] & b[223])^(a[178] & b[224])^(a[177] & b[225])^(a[176] & b[226])^(a[175] & b[227])^(a[174] & b[228])^(a[173] & b[229])^(a[172] & b[230])^(a[171] & b[231])^(a[170] & b[232])^(a[169] & b[233])^(a[168] & b[234])^(a[167] & b[235])^(a[166] & b[236])^(a[165] & b[237])^(a[164] & b[238])^(a[163] & b[239])^(a[162] & b[240])^(a[161] & b[241])^(a[160] & b[242])^(a[159] & b[243])^(a[158] & b[244])^(a[157] & b[245])^(a[156] & b[246])^(a[155] & b[247])^(a[154] & b[248])^(a[153] & b[249])^(a[152] & b[250])^(a[151] & b[251])^(a[150] & b[252])^(a[149] & b[253])^(a[148] & b[254])^(a[147] & b[255])^(a[146] & b[256])^(a[145] & b[257])^(a[144] & b[258])^(a[143] & b[259])^(a[142] & b[260])^(a[141] & b[261])^(a[140] & b[262])^(a[139] & b[263])^(a[138] & b[264])^(a[137] & b[265])^(a[136] & b[266])^(a[135] & b[267])^(a[134] & b[268])^(a[133] & b[269])^(a[132] & b[270])^(a[131] & b[271])^(a[130] & b[272])^(a[129] & b[273])^(a[128] & b[274])^(a[127] & b[275])^(a[126] & b[276])^(a[125] & b[277])^(a[124] & b[278])^(a[123] & b[279])^(a[122] & b[280])^(a[121] & b[281])^(a[120] & b[282])^(a[119] & b[283])^(a[118] & b[284])^(a[117] & b[285])^(a[116] & b[286])^(a[115] & b[287])^(a[114] & b[288])^(a[113] & b[289])^(a[112] & b[290])^(a[111] & b[291])^(a[110] & b[292])^(a[109] & b[293])^(a[108] & b[294])^(a[107] & b[295])^(a[106] & b[296])^(a[105] & b[297])^(a[104] & b[298])^(a[103] & b[299])^(a[102] & b[300])^(a[101] & b[301])^(a[100] & b[302])^(a[99] & b[303])^(a[98] & b[304])^(a[97] & b[305])^(a[96] & b[306])^(a[95] & b[307])^(a[94] & b[308])^(a[93] & b[309])^(a[92] & b[310])^(a[91] & b[311])^(a[90] & b[312])^(a[89] & b[313])^(a[88] & b[314])^(a[87] & b[315])^(a[86] & b[316])^(a[85] & b[317])^(a[84] & b[318])^(a[83] & b[319])^(a[82] & b[320])^(a[81] & b[321])^(a[80] & b[322])^(a[79] & b[323])^(a[78] & b[324])^(a[77] & b[325])^(a[76] & b[326])^(a[75] & b[327])^(a[74] & b[328])^(a[73] & b[329])^(a[72] & b[330])^(a[71] & b[331])^(a[70] & b[332])^(a[69] & b[333])^(a[68] & b[334])^(a[67] & b[335])^(a[66] & b[336])^(a[65] & b[337])^(a[64] & b[338])^(a[63] & b[339])^(a[62] & b[340])^(a[61] & b[341])^(a[60] & b[342])^(a[59] & b[343])^(a[58] & b[344])^(a[57] & b[345])^(a[56] & b[346])^(a[55] & b[347])^(a[54] & b[348])^(a[53] & b[349])^(a[52] & b[350])^(a[51] & b[351])^(a[50] & b[352])^(a[49] & b[353])^(a[48] & b[354])^(a[47] & b[355])^(a[46] & b[356])^(a[45] & b[357])^(a[44] & b[358])^(a[43] & b[359])^(a[42] & b[360])^(a[41] & b[361])^(a[40] & b[362])^(a[39] & b[363])^(a[38] & b[364])^(a[37] & b[365])^(a[36] & b[366])^(a[35] & b[367])^(a[34] & b[368])^(a[33] & b[369])^(a[32] & b[370])^(a[31] & b[371])^(a[30] & b[372])^(a[29] & b[373])^(a[28] & b[374])^(a[27] & b[375])^(a[26] & b[376])^(a[25] & b[377])^(a[24] & b[378])^(a[23] & b[379])^(a[22] & b[380])^(a[21] & b[381])^(a[20] & b[382])^(a[19] & b[383])^(a[18] & b[384])^(a[17] & b[385])^(a[16] & b[386])^(a[15] & b[387])^(a[14] & b[388])^(a[13] & b[389])^(a[12] & b[390])^(a[11] & b[391])^(a[10] & b[392])^(a[9] & b[393])^(a[8] & b[394])^(a[7] & b[395])^(a[6] & b[396])^(a[5] & b[397])^(a[4] & b[398])^(a[3] & b[399])^(a[2] & b[400])^(a[1] & b[401])^(a[0] & b[402]);
assign y[403] = (a[403] & b[0])^(a[402] & b[1])^(a[401] & b[2])^(a[400] & b[3])^(a[399] & b[4])^(a[398] & b[5])^(a[397] & b[6])^(a[396] & b[7])^(a[395] & b[8])^(a[394] & b[9])^(a[393] & b[10])^(a[392] & b[11])^(a[391] & b[12])^(a[390] & b[13])^(a[389] & b[14])^(a[388] & b[15])^(a[387] & b[16])^(a[386] & b[17])^(a[385] & b[18])^(a[384] & b[19])^(a[383] & b[20])^(a[382] & b[21])^(a[381] & b[22])^(a[380] & b[23])^(a[379] & b[24])^(a[378] & b[25])^(a[377] & b[26])^(a[376] & b[27])^(a[375] & b[28])^(a[374] & b[29])^(a[373] & b[30])^(a[372] & b[31])^(a[371] & b[32])^(a[370] & b[33])^(a[369] & b[34])^(a[368] & b[35])^(a[367] & b[36])^(a[366] & b[37])^(a[365] & b[38])^(a[364] & b[39])^(a[363] & b[40])^(a[362] & b[41])^(a[361] & b[42])^(a[360] & b[43])^(a[359] & b[44])^(a[358] & b[45])^(a[357] & b[46])^(a[356] & b[47])^(a[355] & b[48])^(a[354] & b[49])^(a[353] & b[50])^(a[352] & b[51])^(a[351] & b[52])^(a[350] & b[53])^(a[349] & b[54])^(a[348] & b[55])^(a[347] & b[56])^(a[346] & b[57])^(a[345] & b[58])^(a[344] & b[59])^(a[343] & b[60])^(a[342] & b[61])^(a[341] & b[62])^(a[340] & b[63])^(a[339] & b[64])^(a[338] & b[65])^(a[337] & b[66])^(a[336] & b[67])^(a[335] & b[68])^(a[334] & b[69])^(a[333] & b[70])^(a[332] & b[71])^(a[331] & b[72])^(a[330] & b[73])^(a[329] & b[74])^(a[328] & b[75])^(a[327] & b[76])^(a[326] & b[77])^(a[325] & b[78])^(a[324] & b[79])^(a[323] & b[80])^(a[322] & b[81])^(a[321] & b[82])^(a[320] & b[83])^(a[319] & b[84])^(a[318] & b[85])^(a[317] & b[86])^(a[316] & b[87])^(a[315] & b[88])^(a[314] & b[89])^(a[313] & b[90])^(a[312] & b[91])^(a[311] & b[92])^(a[310] & b[93])^(a[309] & b[94])^(a[308] & b[95])^(a[307] & b[96])^(a[306] & b[97])^(a[305] & b[98])^(a[304] & b[99])^(a[303] & b[100])^(a[302] & b[101])^(a[301] & b[102])^(a[300] & b[103])^(a[299] & b[104])^(a[298] & b[105])^(a[297] & b[106])^(a[296] & b[107])^(a[295] & b[108])^(a[294] & b[109])^(a[293] & b[110])^(a[292] & b[111])^(a[291] & b[112])^(a[290] & b[113])^(a[289] & b[114])^(a[288] & b[115])^(a[287] & b[116])^(a[286] & b[117])^(a[285] & b[118])^(a[284] & b[119])^(a[283] & b[120])^(a[282] & b[121])^(a[281] & b[122])^(a[280] & b[123])^(a[279] & b[124])^(a[278] & b[125])^(a[277] & b[126])^(a[276] & b[127])^(a[275] & b[128])^(a[274] & b[129])^(a[273] & b[130])^(a[272] & b[131])^(a[271] & b[132])^(a[270] & b[133])^(a[269] & b[134])^(a[268] & b[135])^(a[267] & b[136])^(a[266] & b[137])^(a[265] & b[138])^(a[264] & b[139])^(a[263] & b[140])^(a[262] & b[141])^(a[261] & b[142])^(a[260] & b[143])^(a[259] & b[144])^(a[258] & b[145])^(a[257] & b[146])^(a[256] & b[147])^(a[255] & b[148])^(a[254] & b[149])^(a[253] & b[150])^(a[252] & b[151])^(a[251] & b[152])^(a[250] & b[153])^(a[249] & b[154])^(a[248] & b[155])^(a[247] & b[156])^(a[246] & b[157])^(a[245] & b[158])^(a[244] & b[159])^(a[243] & b[160])^(a[242] & b[161])^(a[241] & b[162])^(a[240] & b[163])^(a[239] & b[164])^(a[238] & b[165])^(a[237] & b[166])^(a[236] & b[167])^(a[235] & b[168])^(a[234] & b[169])^(a[233] & b[170])^(a[232] & b[171])^(a[231] & b[172])^(a[230] & b[173])^(a[229] & b[174])^(a[228] & b[175])^(a[227] & b[176])^(a[226] & b[177])^(a[225] & b[178])^(a[224] & b[179])^(a[223] & b[180])^(a[222] & b[181])^(a[221] & b[182])^(a[220] & b[183])^(a[219] & b[184])^(a[218] & b[185])^(a[217] & b[186])^(a[216] & b[187])^(a[215] & b[188])^(a[214] & b[189])^(a[213] & b[190])^(a[212] & b[191])^(a[211] & b[192])^(a[210] & b[193])^(a[209] & b[194])^(a[208] & b[195])^(a[207] & b[196])^(a[206] & b[197])^(a[205] & b[198])^(a[204] & b[199])^(a[203] & b[200])^(a[202] & b[201])^(a[201] & b[202])^(a[200] & b[203])^(a[199] & b[204])^(a[198] & b[205])^(a[197] & b[206])^(a[196] & b[207])^(a[195] & b[208])^(a[194] & b[209])^(a[193] & b[210])^(a[192] & b[211])^(a[191] & b[212])^(a[190] & b[213])^(a[189] & b[214])^(a[188] & b[215])^(a[187] & b[216])^(a[186] & b[217])^(a[185] & b[218])^(a[184] & b[219])^(a[183] & b[220])^(a[182] & b[221])^(a[181] & b[222])^(a[180] & b[223])^(a[179] & b[224])^(a[178] & b[225])^(a[177] & b[226])^(a[176] & b[227])^(a[175] & b[228])^(a[174] & b[229])^(a[173] & b[230])^(a[172] & b[231])^(a[171] & b[232])^(a[170] & b[233])^(a[169] & b[234])^(a[168] & b[235])^(a[167] & b[236])^(a[166] & b[237])^(a[165] & b[238])^(a[164] & b[239])^(a[163] & b[240])^(a[162] & b[241])^(a[161] & b[242])^(a[160] & b[243])^(a[159] & b[244])^(a[158] & b[245])^(a[157] & b[246])^(a[156] & b[247])^(a[155] & b[248])^(a[154] & b[249])^(a[153] & b[250])^(a[152] & b[251])^(a[151] & b[252])^(a[150] & b[253])^(a[149] & b[254])^(a[148] & b[255])^(a[147] & b[256])^(a[146] & b[257])^(a[145] & b[258])^(a[144] & b[259])^(a[143] & b[260])^(a[142] & b[261])^(a[141] & b[262])^(a[140] & b[263])^(a[139] & b[264])^(a[138] & b[265])^(a[137] & b[266])^(a[136] & b[267])^(a[135] & b[268])^(a[134] & b[269])^(a[133] & b[270])^(a[132] & b[271])^(a[131] & b[272])^(a[130] & b[273])^(a[129] & b[274])^(a[128] & b[275])^(a[127] & b[276])^(a[126] & b[277])^(a[125] & b[278])^(a[124] & b[279])^(a[123] & b[280])^(a[122] & b[281])^(a[121] & b[282])^(a[120] & b[283])^(a[119] & b[284])^(a[118] & b[285])^(a[117] & b[286])^(a[116] & b[287])^(a[115] & b[288])^(a[114] & b[289])^(a[113] & b[290])^(a[112] & b[291])^(a[111] & b[292])^(a[110] & b[293])^(a[109] & b[294])^(a[108] & b[295])^(a[107] & b[296])^(a[106] & b[297])^(a[105] & b[298])^(a[104] & b[299])^(a[103] & b[300])^(a[102] & b[301])^(a[101] & b[302])^(a[100] & b[303])^(a[99] & b[304])^(a[98] & b[305])^(a[97] & b[306])^(a[96] & b[307])^(a[95] & b[308])^(a[94] & b[309])^(a[93] & b[310])^(a[92] & b[311])^(a[91] & b[312])^(a[90] & b[313])^(a[89] & b[314])^(a[88] & b[315])^(a[87] & b[316])^(a[86] & b[317])^(a[85] & b[318])^(a[84] & b[319])^(a[83] & b[320])^(a[82] & b[321])^(a[81] & b[322])^(a[80] & b[323])^(a[79] & b[324])^(a[78] & b[325])^(a[77] & b[326])^(a[76] & b[327])^(a[75] & b[328])^(a[74] & b[329])^(a[73] & b[330])^(a[72] & b[331])^(a[71] & b[332])^(a[70] & b[333])^(a[69] & b[334])^(a[68] & b[335])^(a[67] & b[336])^(a[66] & b[337])^(a[65] & b[338])^(a[64] & b[339])^(a[63] & b[340])^(a[62] & b[341])^(a[61] & b[342])^(a[60] & b[343])^(a[59] & b[344])^(a[58] & b[345])^(a[57] & b[346])^(a[56] & b[347])^(a[55] & b[348])^(a[54] & b[349])^(a[53] & b[350])^(a[52] & b[351])^(a[51] & b[352])^(a[50] & b[353])^(a[49] & b[354])^(a[48] & b[355])^(a[47] & b[356])^(a[46] & b[357])^(a[45] & b[358])^(a[44] & b[359])^(a[43] & b[360])^(a[42] & b[361])^(a[41] & b[362])^(a[40] & b[363])^(a[39] & b[364])^(a[38] & b[365])^(a[37] & b[366])^(a[36] & b[367])^(a[35] & b[368])^(a[34] & b[369])^(a[33] & b[370])^(a[32] & b[371])^(a[31] & b[372])^(a[30] & b[373])^(a[29] & b[374])^(a[28] & b[375])^(a[27] & b[376])^(a[26] & b[377])^(a[25] & b[378])^(a[24] & b[379])^(a[23] & b[380])^(a[22] & b[381])^(a[21] & b[382])^(a[20] & b[383])^(a[19] & b[384])^(a[18] & b[385])^(a[17] & b[386])^(a[16] & b[387])^(a[15] & b[388])^(a[14] & b[389])^(a[13] & b[390])^(a[12] & b[391])^(a[11] & b[392])^(a[10] & b[393])^(a[9] & b[394])^(a[8] & b[395])^(a[7] & b[396])^(a[6] & b[397])^(a[5] & b[398])^(a[4] & b[399])^(a[3] & b[400])^(a[2] & b[401])^(a[1] & b[402])^(a[0] & b[403]);
assign y[404] = (a[404] & b[0])^(a[403] & b[1])^(a[402] & b[2])^(a[401] & b[3])^(a[400] & b[4])^(a[399] & b[5])^(a[398] & b[6])^(a[397] & b[7])^(a[396] & b[8])^(a[395] & b[9])^(a[394] & b[10])^(a[393] & b[11])^(a[392] & b[12])^(a[391] & b[13])^(a[390] & b[14])^(a[389] & b[15])^(a[388] & b[16])^(a[387] & b[17])^(a[386] & b[18])^(a[385] & b[19])^(a[384] & b[20])^(a[383] & b[21])^(a[382] & b[22])^(a[381] & b[23])^(a[380] & b[24])^(a[379] & b[25])^(a[378] & b[26])^(a[377] & b[27])^(a[376] & b[28])^(a[375] & b[29])^(a[374] & b[30])^(a[373] & b[31])^(a[372] & b[32])^(a[371] & b[33])^(a[370] & b[34])^(a[369] & b[35])^(a[368] & b[36])^(a[367] & b[37])^(a[366] & b[38])^(a[365] & b[39])^(a[364] & b[40])^(a[363] & b[41])^(a[362] & b[42])^(a[361] & b[43])^(a[360] & b[44])^(a[359] & b[45])^(a[358] & b[46])^(a[357] & b[47])^(a[356] & b[48])^(a[355] & b[49])^(a[354] & b[50])^(a[353] & b[51])^(a[352] & b[52])^(a[351] & b[53])^(a[350] & b[54])^(a[349] & b[55])^(a[348] & b[56])^(a[347] & b[57])^(a[346] & b[58])^(a[345] & b[59])^(a[344] & b[60])^(a[343] & b[61])^(a[342] & b[62])^(a[341] & b[63])^(a[340] & b[64])^(a[339] & b[65])^(a[338] & b[66])^(a[337] & b[67])^(a[336] & b[68])^(a[335] & b[69])^(a[334] & b[70])^(a[333] & b[71])^(a[332] & b[72])^(a[331] & b[73])^(a[330] & b[74])^(a[329] & b[75])^(a[328] & b[76])^(a[327] & b[77])^(a[326] & b[78])^(a[325] & b[79])^(a[324] & b[80])^(a[323] & b[81])^(a[322] & b[82])^(a[321] & b[83])^(a[320] & b[84])^(a[319] & b[85])^(a[318] & b[86])^(a[317] & b[87])^(a[316] & b[88])^(a[315] & b[89])^(a[314] & b[90])^(a[313] & b[91])^(a[312] & b[92])^(a[311] & b[93])^(a[310] & b[94])^(a[309] & b[95])^(a[308] & b[96])^(a[307] & b[97])^(a[306] & b[98])^(a[305] & b[99])^(a[304] & b[100])^(a[303] & b[101])^(a[302] & b[102])^(a[301] & b[103])^(a[300] & b[104])^(a[299] & b[105])^(a[298] & b[106])^(a[297] & b[107])^(a[296] & b[108])^(a[295] & b[109])^(a[294] & b[110])^(a[293] & b[111])^(a[292] & b[112])^(a[291] & b[113])^(a[290] & b[114])^(a[289] & b[115])^(a[288] & b[116])^(a[287] & b[117])^(a[286] & b[118])^(a[285] & b[119])^(a[284] & b[120])^(a[283] & b[121])^(a[282] & b[122])^(a[281] & b[123])^(a[280] & b[124])^(a[279] & b[125])^(a[278] & b[126])^(a[277] & b[127])^(a[276] & b[128])^(a[275] & b[129])^(a[274] & b[130])^(a[273] & b[131])^(a[272] & b[132])^(a[271] & b[133])^(a[270] & b[134])^(a[269] & b[135])^(a[268] & b[136])^(a[267] & b[137])^(a[266] & b[138])^(a[265] & b[139])^(a[264] & b[140])^(a[263] & b[141])^(a[262] & b[142])^(a[261] & b[143])^(a[260] & b[144])^(a[259] & b[145])^(a[258] & b[146])^(a[257] & b[147])^(a[256] & b[148])^(a[255] & b[149])^(a[254] & b[150])^(a[253] & b[151])^(a[252] & b[152])^(a[251] & b[153])^(a[250] & b[154])^(a[249] & b[155])^(a[248] & b[156])^(a[247] & b[157])^(a[246] & b[158])^(a[245] & b[159])^(a[244] & b[160])^(a[243] & b[161])^(a[242] & b[162])^(a[241] & b[163])^(a[240] & b[164])^(a[239] & b[165])^(a[238] & b[166])^(a[237] & b[167])^(a[236] & b[168])^(a[235] & b[169])^(a[234] & b[170])^(a[233] & b[171])^(a[232] & b[172])^(a[231] & b[173])^(a[230] & b[174])^(a[229] & b[175])^(a[228] & b[176])^(a[227] & b[177])^(a[226] & b[178])^(a[225] & b[179])^(a[224] & b[180])^(a[223] & b[181])^(a[222] & b[182])^(a[221] & b[183])^(a[220] & b[184])^(a[219] & b[185])^(a[218] & b[186])^(a[217] & b[187])^(a[216] & b[188])^(a[215] & b[189])^(a[214] & b[190])^(a[213] & b[191])^(a[212] & b[192])^(a[211] & b[193])^(a[210] & b[194])^(a[209] & b[195])^(a[208] & b[196])^(a[207] & b[197])^(a[206] & b[198])^(a[205] & b[199])^(a[204] & b[200])^(a[203] & b[201])^(a[202] & b[202])^(a[201] & b[203])^(a[200] & b[204])^(a[199] & b[205])^(a[198] & b[206])^(a[197] & b[207])^(a[196] & b[208])^(a[195] & b[209])^(a[194] & b[210])^(a[193] & b[211])^(a[192] & b[212])^(a[191] & b[213])^(a[190] & b[214])^(a[189] & b[215])^(a[188] & b[216])^(a[187] & b[217])^(a[186] & b[218])^(a[185] & b[219])^(a[184] & b[220])^(a[183] & b[221])^(a[182] & b[222])^(a[181] & b[223])^(a[180] & b[224])^(a[179] & b[225])^(a[178] & b[226])^(a[177] & b[227])^(a[176] & b[228])^(a[175] & b[229])^(a[174] & b[230])^(a[173] & b[231])^(a[172] & b[232])^(a[171] & b[233])^(a[170] & b[234])^(a[169] & b[235])^(a[168] & b[236])^(a[167] & b[237])^(a[166] & b[238])^(a[165] & b[239])^(a[164] & b[240])^(a[163] & b[241])^(a[162] & b[242])^(a[161] & b[243])^(a[160] & b[244])^(a[159] & b[245])^(a[158] & b[246])^(a[157] & b[247])^(a[156] & b[248])^(a[155] & b[249])^(a[154] & b[250])^(a[153] & b[251])^(a[152] & b[252])^(a[151] & b[253])^(a[150] & b[254])^(a[149] & b[255])^(a[148] & b[256])^(a[147] & b[257])^(a[146] & b[258])^(a[145] & b[259])^(a[144] & b[260])^(a[143] & b[261])^(a[142] & b[262])^(a[141] & b[263])^(a[140] & b[264])^(a[139] & b[265])^(a[138] & b[266])^(a[137] & b[267])^(a[136] & b[268])^(a[135] & b[269])^(a[134] & b[270])^(a[133] & b[271])^(a[132] & b[272])^(a[131] & b[273])^(a[130] & b[274])^(a[129] & b[275])^(a[128] & b[276])^(a[127] & b[277])^(a[126] & b[278])^(a[125] & b[279])^(a[124] & b[280])^(a[123] & b[281])^(a[122] & b[282])^(a[121] & b[283])^(a[120] & b[284])^(a[119] & b[285])^(a[118] & b[286])^(a[117] & b[287])^(a[116] & b[288])^(a[115] & b[289])^(a[114] & b[290])^(a[113] & b[291])^(a[112] & b[292])^(a[111] & b[293])^(a[110] & b[294])^(a[109] & b[295])^(a[108] & b[296])^(a[107] & b[297])^(a[106] & b[298])^(a[105] & b[299])^(a[104] & b[300])^(a[103] & b[301])^(a[102] & b[302])^(a[101] & b[303])^(a[100] & b[304])^(a[99] & b[305])^(a[98] & b[306])^(a[97] & b[307])^(a[96] & b[308])^(a[95] & b[309])^(a[94] & b[310])^(a[93] & b[311])^(a[92] & b[312])^(a[91] & b[313])^(a[90] & b[314])^(a[89] & b[315])^(a[88] & b[316])^(a[87] & b[317])^(a[86] & b[318])^(a[85] & b[319])^(a[84] & b[320])^(a[83] & b[321])^(a[82] & b[322])^(a[81] & b[323])^(a[80] & b[324])^(a[79] & b[325])^(a[78] & b[326])^(a[77] & b[327])^(a[76] & b[328])^(a[75] & b[329])^(a[74] & b[330])^(a[73] & b[331])^(a[72] & b[332])^(a[71] & b[333])^(a[70] & b[334])^(a[69] & b[335])^(a[68] & b[336])^(a[67] & b[337])^(a[66] & b[338])^(a[65] & b[339])^(a[64] & b[340])^(a[63] & b[341])^(a[62] & b[342])^(a[61] & b[343])^(a[60] & b[344])^(a[59] & b[345])^(a[58] & b[346])^(a[57] & b[347])^(a[56] & b[348])^(a[55] & b[349])^(a[54] & b[350])^(a[53] & b[351])^(a[52] & b[352])^(a[51] & b[353])^(a[50] & b[354])^(a[49] & b[355])^(a[48] & b[356])^(a[47] & b[357])^(a[46] & b[358])^(a[45] & b[359])^(a[44] & b[360])^(a[43] & b[361])^(a[42] & b[362])^(a[41] & b[363])^(a[40] & b[364])^(a[39] & b[365])^(a[38] & b[366])^(a[37] & b[367])^(a[36] & b[368])^(a[35] & b[369])^(a[34] & b[370])^(a[33] & b[371])^(a[32] & b[372])^(a[31] & b[373])^(a[30] & b[374])^(a[29] & b[375])^(a[28] & b[376])^(a[27] & b[377])^(a[26] & b[378])^(a[25] & b[379])^(a[24] & b[380])^(a[23] & b[381])^(a[22] & b[382])^(a[21] & b[383])^(a[20] & b[384])^(a[19] & b[385])^(a[18] & b[386])^(a[17] & b[387])^(a[16] & b[388])^(a[15] & b[389])^(a[14] & b[390])^(a[13] & b[391])^(a[12] & b[392])^(a[11] & b[393])^(a[10] & b[394])^(a[9] & b[395])^(a[8] & b[396])^(a[7] & b[397])^(a[6] & b[398])^(a[5] & b[399])^(a[4] & b[400])^(a[3] & b[401])^(a[2] & b[402])^(a[1] & b[403])^(a[0] & b[404]);
assign y[405] = (a[405] & b[0])^(a[404] & b[1])^(a[403] & b[2])^(a[402] & b[3])^(a[401] & b[4])^(a[400] & b[5])^(a[399] & b[6])^(a[398] & b[7])^(a[397] & b[8])^(a[396] & b[9])^(a[395] & b[10])^(a[394] & b[11])^(a[393] & b[12])^(a[392] & b[13])^(a[391] & b[14])^(a[390] & b[15])^(a[389] & b[16])^(a[388] & b[17])^(a[387] & b[18])^(a[386] & b[19])^(a[385] & b[20])^(a[384] & b[21])^(a[383] & b[22])^(a[382] & b[23])^(a[381] & b[24])^(a[380] & b[25])^(a[379] & b[26])^(a[378] & b[27])^(a[377] & b[28])^(a[376] & b[29])^(a[375] & b[30])^(a[374] & b[31])^(a[373] & b[32])^(a[372] & b[33])^(a[371] & b[34])^(a[370] & b[35])^(a[369] & b[36])^(a[368] & b[37])^(a[367] & b[38])^(a[366] & b[39])^(a[365] & b[40])^(a[364] & b[41])^(a[363] & b[42])^(a[362] & b[43])^(a[361] & b[44])^(a[360] & b[45])^(a[359] & b[46])^(a[358] & b[47])^(a[357] & b[48])^(a[356] & b[49])^(a[355] & b[50])^(a[354] & b[51])^(a[353] & b[52])^(a[352] & b[53])^(a[351] & b[54])^(a[350] & b[55])^(a[349] & b[56])^(a[348] & b[57])^(a[347] & b[58])^(a[346] & b[59])^(a[345] & b[60])^(a[344] & b[61])^(a[343] & b[62])^(a[342] & b[63])^(a[341] & b[64])^(a[340] & b[65])^(a[339] & b[66])^(a[338] & b[67])^(a[337] & b[68])^(a[336] & b[69])^(a[335] & b[70])^(a[334] & b[71])^(a[333] & b[72])^(a[332] & b[73])^(a[331] & b[74])^(a[330] & b[75])^(a[329] & b[76])^(a[328] & b[77])^(a[327] & b[78])^(a[326] & b[79])^(a[325] & b[80])^(a[324] & b[81])^(a[323] & b[82])^(a[322] & b[83])^(a[321] & b[84])^(a[320] & b[85])^(a[319] & b[86])^(a[318] & b[87])^(a[317] & b[88])^(a[316] & b[89])^(a[315] & b[90])^(a[314] & b[91])^(a[313] & b[92])^(a[312] & b[93])^(a[311] & b[94])^(a[310] & b[95])^(a[309] & b[96])^(a[308] & b[97])^(a[307] & b[98])^(a[306] & b[99])^(a[305] & b[100])^(a[304] & b[101])^(a[303] & b[102])^(a[302] & b[103])^(a[301] & b[104])^(a[300] & b[105])^(a[299] & b[106])^(a[298] & b[107])^(a[297] & b[108])^(a[296] & b[109])^(a[295] & b[110])^(a[294] & b[111])^(a[293] & b[112])^(a[292] & b[113])^(a[291] & b[114])^(a[290] & b[115])^(a[289] & b[116])^(a[288] & b[117])^(a[287] & b[118])^(a[286] & b[119])^(a[285] & b[120])^(a[284] & b[121])^(a[283] & b[122])^(a[282] & b[123])^(a[281] & b[124])^(a[280] & b[125])^(a[279] & b[126])^(a[278] & b[127])^(a[277] & b[128])^(a[276] & b[129])^(a[275] & b[130])^(a[274] & b[131])^(a[273] & b[132])^(a[272] & b[133])^(a[271] & b[134])^(a[270] & b[135])^(a[269] & b[136])^(a[268] & b[137])^(a[267] & b[138])^(a[266] & b[139])^(a[265] & b[140])^(a[264] & b[141])^(a[263] & b[142])^(a[262] & b[143])^(a[261] & b[144])^(a[260] & b[145])^(a[259] & b[146])^(a[258] & b[147])^(a[257] & b[148])^(a[256] & b[149])^(a[255] & b[150])^(a[254] & b[151])^(a[253] & b[152])^(a[252] & b[153])^(a[251] & b[154])^(a[250] & b[155])^(a[249] & b[156])^(a[248] & b[157])^(a[247] & b[158])^(a[246] & b[159])^(a[245] & b[160])^(a[244] & b[161])^(a[243] & b[162])^(a[242] & b[163])^(a[241] & b[164])^(a[240] & b[165])^(a[239] & b[166])^(a[238] & b[167])^(a[237] & b[168])^(a[236] & b[169])^(a[235] & b[170])^(a[234] & b[171])^(a[233] & b[172])^(a[232] & b[173])^(a[231] & b[174])^(a[230] & b[175])^(a[229] & b[176])^(a[228] & b[177])^(a[227] & b[178])^(a[226] & b[179])^(a[225] & b[180])^(a[224] & b[181])^(a[223] & b[182])^(a[222] & b[183])^(a[221] & b[184])^(a[220] & b[185])^(a[219] & b[186])^(a[218] & b[187])^(a[217] & b[188])^(a[216] & b[189])^(a[215] & b[190])^(a[214] & b[191])^(a[213] & b[192])^(a[212] & b[193])^(a[211] & b[194])^(a[210] & b[195])^(a[209] & b[196])^(a[208] & b[197])^(a[207] & b[198])^(a[206] & b[199])^(a[205] & b[200])^(a[204] & b[201])^(a[203] & b[202])^(a[202] & b[203])^(a[201] & b[204])^(a[200] & b[205])^(a[199] & b[206])^(a[198] & b[207])^(a[197] & b[208])^(a[196] & b[209])^(a[195] & b[210])^(a[194] & b[211])^(a[193] & b[212])^(a[192] & b[213])^(a[191] & b[214])^(a[190] & b[215])^(a[189] & b[216])^(a[188] & b[217])^(a[187] & b[218])^(a[186] & b[219])^(a[185] & b[220])^(a[184] & b[221])^(a[183] & b[222])^(a[182] & b[223])^(a[181] & b[224])^(a[180] & b[225])^(a[179] & b[226])^(a[178] & b[227])^(a[177] & b[228])^(a[176] & b[229])^(a[175] & b[230])^(a[174] & b[231])^(a[173] & b[232])^(a[172] & b[233])^(a[171] & b[234])^(a[170] & b[235])^(a[169] & b[236])^(a[168] & b[237])^(a[167] & b[238])^(a[166] & b[239])^(a[165] & b[240])^(a[164] & b[241])^(a[163] & b[242])^(a[162] & b[243])^(a[161] & b[244])^(a[160] & b[245])^(a[159] & b[246])^(a[158] & b[247])^(a[157] & b[248])^(a[156] & b[249])^(a[155] & b[250])^(a[154] & b[251])^(a[153] & b[252])^(a[152] & b[253])^(a[151] & b[254])^(a[150] & b[255])^(a[149] & b[256])^(a[148] & b[257])^(a[147] & b[258])^(a[146] & b[259])^(a[145] & b[260])^(a[144] & b[261])^(a[143] & b[262])^(a[142] & b[263])^(a[141] & b[264])^(a[140] & b[265])^(a[139] & b[266])^(a[138] & b[267])^(a[137] & b[268])^(a[136] & b[269])^(a[135] & b[270])^(a[134] & b[271])^(a[133] & b[272])^(a[132] & b[273])^(a[131] & b[274])^(a[130] & b[275])^(a[129] & b[276])^(a[128] & b[277])^(a[127] & b[278])^(a[126] & b[279])^(a[125] & b[280])^(a[124] & b[281])^(a[123] & b[282])^(a[122] & b[283])^(a[121] & b[284])^(a[120] & b[285])^(a[119] & b[286])^(a[118] & b[287])^(a[117] & b[288])^(a[116] & b[289])^(a[115] & b[290])^(a[114] & b[291])^(a[113] & b[292])^(a[112] & b[293])^(a[111] & b[294])^(a[110] & b[295])^(a[109] & b[296])^(a[108] & b[297])^(a[107] & b[298])^(a[106] & b[299])^(a[105] & b[300])^(a[104] & b[301])^(a[103] & b[302])^(a[102] & b[303])^(a[101] & b[304])^(a[100] & b[305])^(a[99] & b[306])^(a[98] & b[307])^(a[97] & b[308])^(a[96] & b[309])^(a[95] & b[310])^(a[94] & b[311])^(a[93] & b[312])^(a[92] & b[313])^(a[91] & b[314])^(a[90] & b[315])^(a[89] & b[316])^(a[88] & b[317])^(a[87] & b[318])^(a[86] & b[319])^(a[85] & b[320])^(a[84] & b[321])^(a[83] & b[322])^(a[82] & b[323])^(a[81] & b[324])^(a[80] & b[325])^(a[79] & b[326])^(a[78] & b[327])^(a[77] & b[328])^(a[76] & b[329])^(a[75] & b[330])^(a[74] & b[331])^(a[73] & b[332])^(a[72] & b[333])^(a[71] & b[334])^(a[70] & b[335])^(a[69] & b[336])^(a[68] & b[337])^(a[67] & b[338])^(a[66] & b[339])^(a[65] & b[340])^(a[64] & b[341])^(a[63] & b[342])^(a[62] & b[343])^(a[61] & b[344])^(a[60] & b[345])^(a[59] & b[346])^(a[58] & b[347])^(a[57] & b[348])^(a[56] & b[349])^(a[55] & b[350])^(a[54] & b[351])^(a[53] & b[352])^(a[52] & b[353])^(a[51] & b[354])^(a[50] & b[355])^(a[49] & b[356])^(a[48] & b[357])^(a[47] & b[358])^(a[46] & b[359])^(a[45] & b[360])^(a[44] & b[361])^(a[43] & b[362])^(a[42] & b[363])^(a[41] & b[364])^(a[40] & b[365])^(a[39] & b[366])^(a[38] & b[367])^(a[37] & b[368])^(a[36] & b[369])^(a[35] & b[370])^(a[34] & b[371])^(a[33] & b[372])^(a[32] & b[373])^(a[31] & b[374])^(a[30] & b[375])^(a[29] & b[376])^(a[28] & b[377])^(a[27] & b[378])^(a[26] & b[379])^(a[25] & b[380])^(a[24] & b[381])^(a[23] & b[382])^(a[22] & b[383])^(a[21] & b[384])^(a[20] & b[385])^(a[19] & b[386])^(a[18] & b[387])^(a[17] & b[388])^(a[16] & b[389])^(a[15] & b[390])^(a[14] & b[391])^(a[13] & b[392])^(a[12] & b[393])^(a[11] & b[394])^(a[10] & b[395])^(a[9] & b[396])^(a[8] & b[397])^(a[7] & b[398])^(a[6] & b[399])^(a[5] & b[400])^(a[4] & b[401])^(a[3] & b[402])^(a[2] & b[403])^(a[1] & b[404])^(a[0] & b[405]);
assign y[406] = (a[406] & b[0])^(a[405] & b[1])^(a[404] & b[2])^(a[403] & b[3])^(a[402] & b[4])^(a[401] & b[5])^(a[400] & b[6])^(a[399] & b[7])^(a[398] & b[8])^(a[397] & b[9])^(a[396] & b[10])^(a[395] & b[11])^(a[394] & b[12])^(a[393] & b[13])^(a[392] & b[14])^(a[391] & b[15])^(a[390] & b[16])^(a[389] & b[17])^(a[388] & b[18])^(a[387] & b[19])^(a[386] & b[20])^(a[385] & b[21])^(a[384] & b[22])^(a[383] & b[23])^(a[382] & b[24])^(a[381] & b[25])^(a[380] & b[26])^(a[379] & b[27])^(a[378] & b[28])^(a[377] & b[29])^(a[376] & b[30])^(a[375] & b[31])^(a[374] & b[32])^(a[373] & b[33])^(a[372] & b[34])^(a[371] & b[35])^(a[370] & b[36])^(a[369] & b[37])^(a[368] & b[38])^(a[367] & b[39])^(a[366] & b[40])^(a[365] & b[41])^(a[364] & b[42])^(a[363] & b[43])^(a[362] & b[44])^(a[361] & b[45])^(a[360] & b[46])^(a[359] & b[47])^(a[358] & b[48])^(a[357] & b[49])^(a[356] & b[50])^(a[355] & b[51])^(a[354] & b[52])^(a[353] & b[53])^(a[352] & b[54])^(a[351] & b[55])^(a[350] & b[56])^(a[349] & b[57])^(a[348] & b[58])^(a[347] & b[59])^(a[346] & b[60])^(a[345] & b[61])^(a[344] & b[62])^(a[343] & b[63])^(a[342] & b[64])^(a[341] & b[65])^(a[340] & b[66])^(a[339] & b[67])^(a[338] & b[68])^(a[337] & b[69])^(a[336] & b[70])^(a[335] & b[71])^(a[334] & b[72])^(a[333] & b[73])^(a[332] & b[74])^(a[331] & b[75])^(a[330] & b[76])^(a[329] & b[77])^(a[328] & b[78])^(a[327] & b[79])^(a[326] & b[80])^(a[325] & b[81])^(a[324] & b[82])^(a[323] & b[83])^(a[322] & b[84])^(a[321] & b[85])^(a[320] & b[86])^(a[319] & b[87])^(a[318] & b[88])^(a[317] & b[89])^(a[316] & b[90])^(a[315] & b[91])^(a[314] & b[92])^(a[313] & b[93])^(a[312] & b[94])^(a[311] & b[95])^(a[310] & b[96])^(a[309] & b[97])^(a[308] & b[98])^(a[307] & b[99])^(a[306] & b[100])^(a[305] & b[101])^(a[304] & b[102])^(a[303] & b[103])^(a[302] & b[104])^(a[301] & b[105])^(a[300] & b[106])^(a[299] & b[107])^(a[298] & b[108])^(a[297] & b[109])^(a[296] & b[110])^(a[295] & b[111])^(a[294] & b[112])^(a[293] & b[113])^(a[292] & b[114])^(a[291] & b[115])^(a[290] & b[116])^(a[289] & b[117])^(a[288] & b[118])^(a[287] & b[119])^(a[286] & b[120])^(a[285] & b[121])^(a[284] & b[122])^(a[283] & b[123])^(a[282] & b[124])^(a[281] & b[125])^(a[280] & b[126])^(a[279] & b[127])^(a[278] & b[128])^(a[277] & b[129])^(a[276] & b[130])^(a[275] & b[131])^(a[274] & b[132])^(a[273] & b[133])^(a[272] & b[134])^(a[271] & b[135])^(a[270] & b[136])^(a[269] & b[137])^(a[268] & b[138])^(a[267] & b[139])^(a[266] & b[140])^(a[265] & b[141])^(a[264] & b[142])^(a[263] & b[143])^(a[262] & b[144])^(a[261] & b[145])^(a[260] & b[146])^(a[259] & b[147])^(a[258] & b[148])^(a[257] & b[149])^(a[256] & b[150])^(a[255] & b[151])^(a[254] & b[152])^(a[253] & b[153])^(a[252] & b[154])^(a[251] & b[155])^(a[250] & b[156])^(a[249] & b[157])^(a[248] & b[158])^(a[247] & b[159])^(a[246] & b[160])^(a[245] & b[161])^(a[244] & b[162])^(a[243] & b[163])^(a[242] & b[164])^(a[241] & b[165])^(a[240] & b[166])^(a[239] & b[167])^(a[238] & b[168])^(a[237] & b[169])^(a[236] & b[170])^(a[235] & b[171])^(a[234] & b[172])^(a[233] & b[173])^(a[232] & b[174])^(a[231] & b[175])^(a[230] & b[176])^(a[229] & b[177])^(a[228] & b[178])^(a[227] & b[179])^(a[226] & b[180])^(a[225] & b[181])^(a[224] & b[182])^(a[223] & b[183])^(a[222] & b[184])^(a[221] & b[185])^(a[220] & b[186])^(a[219] & b[187])^(a[218] & b[188])^(a[217] & b[189])^(a[216] & b[190])^(a[215] & b[191])^(a[214] & b[192])^(a[213] & b[193])^(a[212] & b[194])^(a[211] & b[195])^(a[210] & b[196])^(a[209] & b[197])^(a[208] & b[198])^(a[207] & b[199])^(a[206] & b[200])^(a[205] & b[201])^(a[204] & b[202])^(a[203] & b[203])^(a[202] & b[204])^(a[201] & b[205])^(a[200] & b[206])^(a[199] & b[207])^(a[198] & b[208])^(a[197] & b[209])^(a[196] & b[210])^(a[195] & b[211])^(a[194] & b[212])^(a[193] & b[213])^(a[192] & b[214])^(a[191] & b[215])^(a[190] & b[216])^(a[189] & b[217])^(a[188] & b[218])^(a[187] & b[219])^(a[186] & b[220])^(a[185] & b[221])^(a[184] & b[222])^(a[183] & b[223])^(a[182] & b[224])^(a[181] & b[225])^(a[180] & b[226])^(a[179] & b[227])^(a[178] & b[228])^(a[177] & b[229])^(a[176] & b[230])^(a[175] & b[231])^(a[174] & b[232])^(a[173] & b[233])^(a[172] & b[234])^(a[171] & b[235])^(a[170] & b[236])^(a[169] & b[237])^(a[168] & b[238])^(a[167] & b[239])^(a[166] & b[240])^(a[165] & b[241])^(a[164] & b[242])^(a[163] & b[243])^(a[162] & b[244])^(a[161] & b[245])^(a[160] & b[246])^(a[159] & b[247])^(a[158] & b[248])^(a[157] & b[249])^(a[156] & b[250])^(a[155] & b[251])^(a[154] & b[252])^(a[153] & b[253])^(a[152] & b[254])^(a[151] & b[255])^(a[150] & b[256])^(a[149] & b[257])^(a[148] & b[258])^(a[147] & b[259])^(a[146] & b[260])^(a[145] & b[261])^(a[144] & b[262])^(a[143] & b[263])^(a[142] & b[264])^(a[141] & b[265])^(a[140] & b[266])^(a[139] & b[267])^(a[138] & b[268])^(a[137] & b[269])^(a[136] & b[270])^(a[135] & b[271])^(a[134] & b[272])^(a[133] & b[273])^(a[132] & b[274])^(a[131] & b[275])^(a[130] & b[276])^(a[129] & b[277])^(a[128] & b[278])^(a[127] & b[279])^(a[126] & b[280])^(a[125] & b[281])^(a[124] & b[282])^(a[123] & b[283])^(a[122] & b[284])^(a[121] & b[285])^(a[120] & b[286])^(a[119] & b[287])^(a[118] & b[288])^(a[117] & b[289])^(a[116] & b[290])^(a[115] & b[291])^(a[114] & b[292])^(a[113] & b[293])^(a[112] & b[294])^(a[111] & b[295])^(a[110] & b[296])^(a[109] & b[297])^(a[108] & b[298])^(a[107] & b[299])^(a[106] & b[300])^(a[105] & b[301])^(a[104] & b[302])^(a[103] & b[303])^(a[102] & b[304])^(a[101] & b[305])^(a[100] & b[306])^(a[99] & b[307])^(a[98] & b[308])^(a[97] & b[309])^(a[96] & b[310])^(a[95] & b[311])^(a[94] & b[312])^(a[93] & b[313])^(a[92] & b[314])^(a[91] & b[315])^(a[90] & b[316])^(a[89] & b[317])^(a[88] & b[318])^(a[87] & b[319])^(a[86] & b[320])^(a[85] & b[321])^(a[84] & b[322])^(a[83] & b[323])^(a[82] & b[324])^(a[81] & b[325])^(a[80] & b[326])^(a[79] & b[327])^(a[78] & b[328])^(a[77] & b[329])^(a[76] & b[330])^(a[75] & b[331])^(a[74] & b[332])^(a[73] & b[333])^(a[72] & b[334])^(a[71] & b[335])^(a[70] & b[336])^(a[69] & b[337])^(a[68] & b[338])^(a[67] & b[339])^(a[66] & b[340])^(a[65] & b[341])^(a[64] & b[342])^(a[63] & b[343])^(a[62] & b[344])^(a[61] & b[345])^(a[60] & b[346])^(a[59] & b[347])^(a[58] & b[348])^(a[57] & b[349])^(a[56] & b[350])^(a[55] & b[351])^(a[54] & b[352])^(a[53] & b[353])^(a[52] & b[354])^(a[51] & b[355])^(a[50] & b[356])^(a[49] & b[357])^(a[48] & b[358])^(a[47] & b[359])^(a[46] & b[360])^(a[45] & b[361])^(a[44] & b[362])^(a[43] & b[363])^(a[42] & b[364])^(a[41] & b[365])^(a[40] & b[366])^(a[39] & b[367])^(a[38] & b[368])^(a[37] & b[369])^(a[36] & b[370])^(a[35] & b[371])^(a[34] & b[372])^(a[33] & b[373])^(a[32] & b[374])^(a[31] & b[375])^(a[30] & b[376])^(a[29] & b[377])^(a[28] & b[378])^(a[27] & b[379])^(a[26] & b[380])^(a[25] & b[381])^(a[24] & b[382])^(a[23] & b[383])^(a[22] & b[384])^(a[21] & b[385])^(a[20] & b[386])^(a[19] & b[387])^(a[18] & b[388])^(a[17] & b[389])^(a[16] & b[390])^(a[15] & b[391])^(a[14] & b[392])^(a[13] & b[393])^(a[12] & b[394])^(a[11] & b[395])^(a[10] & b[396])^(a[9] & b[397])^(a[8] & b[398])^(a[7] & b[399])^(a[6] & b[400])^(a[5] & b[401])^(a[4] & b[402])^(a[3] & b[403])^(a[2] & b[404])^(a[1] & b[405])^(a[0] & b[406]);
assign y[407] = (a[407] & b[0])^(a[406] & b[1])^(a[405] & b[2])^(a[404] & b[3])^(a[403] & b[4])^(a[402] & b[5])^(a[401] & b[6])^(a[400] & b[7])^(a[399] & b[8])^(a[398] & b[9])^(a[397] & b[10])^(a[396] & b[11])^(a[395] & b[12])^(a[394] & b[13])^(a[393] & b[14])^(a[392] & b[15])^(a[391] & b[16])^(a[390] & b[17])^(a[389] & b[18])^(a[388] & b[19])^(a[387] & b[20])^(a[386] & b[21])^(a[385] & b[22])^(a[384] & b[23])^(a[383] & b[24])^(a[382] & b[25])^(a[381] & b[26])^(a[380] & b[27])^(a[379] & b[28])^(a[378] & b[29])^(a[377] & b[30])^(a[376] & b[31])^(a[375] & b[32])^(a[374] & b[33])^(a[373] & b[34])^(a[372] & b[35])^(a[371] & b[36])^(a[370] & b[37])^(a[369] & b[38])^(a[368] & b[39])^(a[367] & b[40])^(a[366] & b[41])^(a[365] & b[42])^(a[364] & b[43])^(a[363] & b[44])^(a[362] & b[45])^(a[361] & b[46])^(a[360] & b[47])^(a[359] & b[48])^(a[358] & b[49])^(a[357] & b[50])^(a[356] & b[51])^(a[355] & b[52])^(a[354] & b[53])^(a[353] & b[54])^(a[352] & b[55])^(a[351] & b[56])^(a[350] & b[57])^(a[349] & b[58])^(a[348] & b[59])^(a[347] & b[60])^(a[346] & b[61])^(a[345] & b[62])^(a[344] & b[63])^(a[343] & b[64])^(a[342] & b[65])^(a[341] & b[66])^(a[340] & b[67])^(a[339] & b[68])^(a[338] & b[69])^(a[337] & b[70])^(a[336] & b[71])^(a[335] & b[72])^(a[334] & b[73])^(a[333] & b[74])^(a[332] & b[75])^(a[331] & b[76])^(a[330] & b[77])^(a[329] & b[78])^(a[328] & b[79])^(a[327] & b[80])^(a[326] & b[81])^(a[325] & b[82])^(a[324] & b[83])^(a[323] & b[84])^(a[322] & b[85])^(a[321] & b[86])^(a[320] & b[87])^(a[319] & b[88])^(a[318] & b[89])^(a[317] & b[90])^(a[316] & b[91])^(a[315] & b[92])^(a[314] & b[93])^(a[313] & b[94])^(a[312] & b[95])^(a[311] & b[96])^(a[310] & b[97])^(a[309] & b[98])^(a[308] & b[99])^(a[307] & b[100])^(a[306] & b[101])^(a[305] & b[102])^(a[304] & b[103])^(a[303] & b[104])^(a[302] & b[105])^(a[301] & b[106])^(a[300] & b[107])^(a[299] & b[108])^(a[298] & b[109])^(a[297] & b[110])^(a[296] & b[111])^(a[295] & b[112])^(a[294] & b[113])^(a[293] & b[114])^(a[292] & b[115])^(a[291] & b[116])^(a[290] & b[117])^(a[289] & b[118])^(a[288] & b[119])^(a[287] & b[120])^(a[286] & b[121])^(a[285] & b[122])^(a[284] & b[123])^(a[283] & b[124])^(a[282] & b[125])^(a[281] & b[126])^(a[280] & b[127])^(a[279] & b[128])^(a[278] & b[129])^(a[277] & b[130])^(a[276] & b[131])^(a[275] & b[132])^(a[274] & b[133])^(a[273] & b[134])^(a[272] & b[135])^(a[271] & b[136])^(a[270] & b[137])^(a[269] & b[138])^(a[268] & b[139])^(a[267] & b[140])^(a[266] & b[141])^(a[265] & b[142])^(a[264] & b[143])^(a[263] & b[144])^(a[262] & b[145])^(a[261] & b[146])^(a[260] & b[147])^(a[259] & b[148])^(a[258] & b[149])^(a[257] & b[150])^(a[256] & b[151])^(a[255] & b[152])^(a[254] & b[153])^(a[253] & b[154])^(a[252] & b[155])^(a[251] & b[156])^(a[250] & b[157])^(a[249] & b[158])^(a[248] & b[159])^(a[247] & b[160])^(a[246] & b[161])^(a[245] & b[162])^(a[244] & b[163])^(a[243] & b[164])^(a[242] & b[165])^(a[241] & b[166])^(a[240] & b[167])^(a[239] & b[168])^(a[238] & b[169])^(a[237] & b[170])^(a[236] & b[171])^(a[235] & b[172])^(a[234] & b[173])^(a[233] & b[174])^(a[232] & b[175])^(a[231] & b[176])^(a[230] & b[177])^(a[229] & b[178])^(a[228] & b[179])^(a[227] & b[180])^(a[226] & b[181])^(a[225] & b[182])^(a[224] & b[183])^(a[223] & b[184])^(a[222] & b[185])^(a[221] & b[186])^(a[220] & b[187])^(a[219] & b[188])^(a[218] & b[189])^(a[217] & b[190])^(a[216] & b[191])^(a[215] & b[192])^(a[214] & b[193])^(a[213] & b[194])^(a[212] & b[195])^(a[211] & b[196])^(a[210] & b[197])^(a[209] & b[198])^(a[208] & b[199])^(a[207] & b[200])^(a[206] & b[201])^(a[205] & b[202])^(a[204] & b[203])^(a[203] & b[204])^(a[202] & b[205])^(a[201] & b[206])^(a[200] & b[207])^(a[199] & b[208])^(a[198] & b[209])^(a[197] & b[210])^(a[196] & b[211])^(a[195] & b[212])^(a[194] & b[213])^(a[193] & b[214])^(a[192] & b[215])^(a[191] & b[216])^(a[190] & b[217])^(a[189] & b[218])^(a[188] & b[219])^(a[187] & b[220])^(a[186] & b[221])^(a[185] & b[222])^(a[184] & b[223])^(a[183] & b[224])^(a[182] & b[225])^(a[181] & b[226])^(a[180] & b[227])^(a[179] & b[228])^(a[178] & b[229])^(a[177] & b[230])^(a[176] & b[231])^(a[175] & b[232])^(a[174] & b[233])^(a[173] & b[234])^(a[172] & b[235])^(a[171] & b[236])^(a[170] & b[237])^(a[169] & b[238])^(a[168] & b[239])^(a[167] & b[240])^(a[166] & b[241])^(a[165] & b[242])^(a[164] & b[243])^(a[163] & b[244])^(a[162] & b[245])^(a[161] & b[246])^(a[160] & b[247])^(a[159] & b[248])^(a[158] & b[249])^(a[157] & b[250])^(a[156] & b[251])^(a[155] & b[252])^(a[154] & b[253])^(a[153] & b[254])^(a[152] & b[255])^(a[151] & b[256])^(a[150] & b[257])^(a[149] & b[258])^(a[148] & b[259])^(a[147] & b[260])^(a[146] & b[261])^(a[145] & b[262])^(a[144] & b[263])^(a[143] & b[264])^(a[142] & b[265])^(a[141] & b[266])^(a[140] & b[267])^(a[139] & b[268])^(a[138] & b[269])^(a[137] & b[270])^(a[136] & b[271])^(a[135] & b[272])^(a[134] & b[273])^(a[133] & b[274])^(a[132] & b[275])^(a[131] & b[276])^(a[130] & b[277])^(a[129] & b[278])^(a[128] & b[279])^(a[127] & b[280])^(a[126] & b[281])^(a[125] & b[282])^(a[124] & b[283])^(a[123] & b[284])^(a[122] & b[285])^(a[121] & b[286])^(a[120] & b[287])^(a[119] & b[288])^(a[118] & b[289])^(a[117] & b[290])^(a[116] & b[291])^(a[115] & b[292])^(a[114] & b[293])^(a[113] & b[294])^(a[112] & b[295])^(a[111] & b[296])^(a[110] & b[297])^(a[109] & b[298])^(a[108] & b[299])^(a[107] & b[300])^(a[106] & b[301])^(a[105] & b[302])^(a[104] & b[303])^(a[103] & b[304])^(a[102] & b[305])^(a[101] & b[306])^(a[100] & b[307])^(a[99] & b[308])^(a[98] & b[309])^(a[97] & b[310])^(a[96] & b[311])^(a[95] & b[312])^(a[94] & b[313])^(a[93] & b[314])^(a[92] & b[315])^(a[91] & b[316])^(a[90] & b[317])^(a[89] & b[318])^(a[88] & b[319])^(a[87] & b[320])^(a[86] & b[321])^(a[85] & b[322])^(a[84] & b[323])^(a[83] & b[324])^(a[82] & b[325])^(a[81] & b[326])^(a[80] & b[327])^(a[79] & b[328])^(a[78] & b[329])^(a[77] & b[330])^(a[76] & b[331])^(a[75] & b[332])^(a[74] & b[333])^(a[73] & b[334])^(a[72] & b[335])^(a[71] & b[336])^(a[70] & b[337])^(a[69] & b[338])^(a[68] & b[339])^(a[67] & b[340])^(a[66] & b[341])^(a[65] & b[342])^(a[64] & b[343])^(a[63] & b[344])^(a[62] & b[345])^(a[61] & b[346])^(a[60] & b[347])^(a[59] & b[348])^(a[58] & b[349])^(a[57] & b[350])^(a[56] & b[351])^(a[55] & b[352])^(a[54] & b[353])^(a[53] & b[354])^(a[52] & b[355])^(a[51] & b[356])^(a[50] & b[357])^(a[49] & b[358])^(a[48] & b[359])^(a[47] & b[360])^(a[46] & b[361])^(a[45] & b[362])^(a[44] & b[363])^(a[43] & b[364])^(a[42] & b[365])^(a[41] & b[366])^(a[40] & b[367])^(a[39] & b[368])^(a[38] & b[369])^(a[37] & b[370])^(a[36] & b[371])^(a[35] & b[372])^(a[34] & b[373])^(a[33] & b[374])^(a[32] & b[375])^(a[31] & b[376])^(a[30] & b[377])^(a[29] & b[378])^(a[28] & b[379])^(a[27] & b[380])^(a[26] & b[381])^(a[25] & b[382])^(a[24] & b[383])^(a[23] & b[384])^(a[22] & b[385])^(a[21] & b[386])^(a[20] & b[387])^(a[19] & b[388])^(a[18] & b[389])^(a[17] & b[390])^(a[16] & b[391])^(a[15] & b[392])^(a[14] & b[393])^(a[13] & b[394])^(a[12] & b[395])^(a[11] & b[396])^(a[10] & b[397])^(a[9] & b[398])^(a[8] & b[399])^(a[7] & b[400])^(a[6] & b[401])^(a[5] & b[402])^(a[4] & b[403])^(a[3] & b[404])^(a[2] & b[405])^(a[1] & b[406])^(a[0] & b[407]);
assign y[408] = (a[408] & b[0])^(a[407] & b[1])^(a[406] & b[2])^(a[405] & b[3])^(a[404] & b[4])^(a[403] & b[5])^(a[402] & b[6])^(a[401] & b[7])^(a[400] & b[8])^(a[399] & b[9])^(a[398] & b[10])^(a[397] & b[11])^(a[396] & b[12])^(a[395] & b[13])^(a[394] & b[14])^(a[393] & b[15])^(a[392] & b[16])^(a[391] & b[17])^(a[390] & b[18])^(a[389] & b[19])^(a[388] & b[20])^(a[387] & b[21])^(a[386] & b[22])^(a[385] & b[23])^(a[384] & b[24])^(a[383] & b[25])^(a[382] & b[26])^(a[381] & b[27])^(a[380] & b[28])^(a[379] & b[29])^(a[378] & b[30])^(a[377] & b[31])^(a[376] & b[32])^(a[375] & b[33])^(a[374] & b[34])^(a[373] & b[35])^(a[372] & b[36])^(a[371] & b[37])^(a[370] & b[38])^(a[369] & b[39])^(a[368] & b[40])^(a[367] & b[41])^(a[366] & b[42])^(a[365] & b[43])^(a[364] & b[44])^(a[363] & b[45])^(a[362] & b[46])^(a[361] & b[47])^(a[360] & b[48])^(a[359] & b[49])^(a[358] & b[50])^(a[357] & b[51])^(a[356] & b[52])^(a[355] & b[53])^(a[354] & b[54])^(a[353] & b[55])^(a[352] & b[56])^(a[351] & b[57])^(a[350] & b[58])^(a[349] & b[59])^(a[348] & b[60])^(a[347] & b[61])^(a[346] & b[62])^(a[345] & b[63])^(a[344] & b[64])^(a[343] & b[65])^(a[342] & b[66])^(a[341] & b[67])^(a[340] & b[68])^(a[339] & b[69])^(a[338] & b[70])^(a[337] & b[71])^(a[336] & b[72])^(a[335] & b[73])^(a[334] & b[74])^(a[333] & b[75])^(a[332] & b[76])^(a[331] & b[77])^(a[330] & b[78])^(a[329] & b[79])^(a[328] & b[80])^(a[327] & b[81])^(a[326] & b[82])^(a[325] & b[83])^(a[324] & b[84])^(a[323] & b[85])^(a[322] & b[86])^(a[321] & b[87])^(a[320] & b[88])^(a[319] & b[89])^(a[318] & b[90])^(a[317] & b[91])^(a[316] & b[92])^(a[315] & b[93])^(a[314] & b[94])^(a[313] & b[95])^(a[312] & b[96])^(a[311] & b[97])^(a[310] & b[98])^(a[309] & b[99])^(a[308] & b[100])^(a[307] & b[101])^(a[306] & b[102])^(a[305] & b[103])^(a[304] & b[104])^(a[303] & b[105])^(a[302] & b[106])^(a[301] & b[107])^(a[300] & b[108])^(a[299] & b[109])^(a[298] & b[110])^(a[297] & b[111])^(a[296] & b[112])^(a[295] & b[113])^(a[294] & b[114])^(a[293] & b[115])^(a[292] & b[116])^(a[291] & b[117])^(a[290] & b[118])^(a[289] & b[119])^(a[288] & b[120])^(a[287] & b[121])^(a[286] & b[122])^(a[285] & b[123])^(a[284] & b[124])^(a[283] & b[125])^(a[282] & b[126])^(a[281] & b[127])^(a[280] & b[128])^(a[279] & b[129])^(a[278] & b[130])^(a[277] & b[131])^(a[276] & b[132])^(a[275] & b[133])^(a[274] & b[134])^(a[273] & b[135])^(a[272] & b[136])^(a[271] & b[137])^(a[270] & b[138])^(a[269] & b[139])^(a[268] & b[140])^(a[267] & b[141])^(a[266] & b[142])^(a[265] & b[143])^(a[264] & b[144])^(a[263] & b[145])^(a[262] & b[146])^(a[261] & b[147])^(a[260] & b[148])^(a[259] & b[149])^(a[258] & b[150])^(a[257] & b[151])^(a[256] & b[152])^(a[255] & b[153])^(a[254] & b[154])^(a[253] & b[155])^(a[252] & b[156])^(a[251] & b[157])^(a[250] & b[158])^(a[249] & b[159])^(a[248] & b[160])^(a[247] & b[161])^(a[246] & b[162])^(a[245] & b[163])^(a[244] & b[164])^(a[243] & b[165])^(a[242] & b[166])^(a[241] & b[167])^(a[240] & b[168])^(a[239] & b[169])^(a[238] & b[170])^(a[237] & b[171])^(a[236] & b[172])^(a[235] & b[173])^(a[234] & b[174])^(a[233] & b[175])^(a[232] & b[176])^(a[231] & b[177])^(a[230] & b[178])^(a[229] & b[179])^(a[228] & b[180])^(a[227] & b[181])^(a[226] & b[182])^(a[225] & b[183])^(a[224] & b[184])^(a[223] & b[185])^(a[222] & b[186])^(a[221] & b[187])^(a[220] & b[188])^(a[219] & b[189])^(a[218] & b[190])^(a[217] & b[191])^(a[216] & b[192])^(a[215] & b[193])^(a[214] & b[194])^(a[213] & b[195])^(a[212] & b[196])^(a[211] & b[197])^(a[210] & b[198])^(a[209] & b[199])^(a[208] & b[200])^(a[207] & b[201])^(a[206] & b[202])^(a[205] & b[203])^(a[204] & b[204])^(a[203] & b[205])^(a[202] & b[206])^(a[201] & b[207])^(a[200] & b[208])^(a[199] & b[209])^(a[198] & b[210])^(a[197] & b[211])^(a[196] & b[212])^(a[195] & b[213])^(a[194] & b[214])^(a[193] & b[215])^(a[192] & b[216])^(a[191] & b[217])^(a[190] & b[218])^(a[189] & b[219])^(a[188] & b[220])^(a[187] & b[221])^(a[186] & b[222])^(a[185] & b[223])^(a[184] & b[224])^(a[183] & b[225])^(a[182] & b[226])^(a[181] & b[227])^(a[180] & b[228])^(a[179] & b[229])^(a[178] & b[230])^(a[177] & b[231])^(a[176] & b[232])^(a[175] & b[233])^(a[174] & b[234])^(a[173] & b[235])^(a[172] & b[236])^(a[171] & b[237])^(a[170] & b[238])^(a[169] & b[239])^(a[168] & b[240])^(a[167] & b[241])^(a[166] & b[242])^(a[165] & b[243])^(a[164] & b[244])^(a[163] & b[245])^(a[162] & b[246])^(a[161] & b[247])^(a[160] & b[248])^(a[159] & b[249])^(a[158] & b[250])^(a[157] & b[251])^(a[156] & b[252])^(a[155] & b[253])^(a[154] & b[254])^(a[153] & b[255])^(a[152] & b[256])^(a[151] & b[257])^(a[150] & b[258])^(a[149] & b[259])^(a[148] & b[260])^(a[147] & b[261])^(a[146] & b[262])^(a[145] & b[263])^(a[144] & b[264])^(a[143] & b[265])^(a[142] & b[266])^(a[141] & b[267])^(a[140] & b[268])^(a[139] & b[269])^(a[138] & b[270])^(a[137] & b[271])^(a[136] & b[272])^(a[135] & b[273])^(a[134] & b[274])^(a[133] & b[275])^(a[132] & b[276])^(a[131] & b[277])^(a[130] & b[278])^(a[129] & b[279])^(a[128] & b[280])^(a[127] & b[281])^(a[126] & b[282])^(a[125] & b[283])^(a[124] & b[284])^(a[123] & b[285])^(a[122] & b[286])^(a[121] & b[287])^(a[120] & b[288])^(a[119] & b[289])^(a[118] & b[290])^(a[117] & b[291])^(a[116] & b[292])^(a[115] & b[293])^(a[114] & b[294])^(a[113] & b[295])^(a[112] & b[296])^(a[111] & b[297])^(a[110] & b[298])^(a[109] & b[299])^(a[108] & b[300])^(a[107] & b[301])^(a[106] & b[302])^(a[105] & b[303])^(a[104] & b[304])^(a[103] & b[305])^(a[102] & b[306])^(a[101] & b[307])^(a[100] & b[308])^(a[99] & b[309])^(a[98] & b[310])^(a[97] & b[311])^(a[96] & b[312])^(a[95] & b[313])^(a[94] & b[314])^(a[93] & b[315])^(a[92] & b[316])^(a[91] & b[317])^(a[90] & b[318])^(a[89] & b[319])^(a[88] & b[320])^(a[87] & b[321])^(a[86] & b[322])^(a[85] & b[323])^(a[84] & b[324])^(a[83] & b[325])^(a[82] & b[326])^(a[81] & b[327])^(a[80] & b[328])^(a[79] & b[329])^(a[78] & b[330])^(a[77] & b[331])^(a[76] & b[332])^(a[75] & b[333])^(a[74] & b[334])^(a[73] & b[335])^(a[72] & b[336])^(a[71] & b[337])^(a[70] & b[338])^(a[69] & b[339])^(a[68] & b[340])^(a[67] & b[341])^(a[66] & b[342])^(a[65] & b[343])^(a[64] & b[344])^(a[63] & b[345])^(a[62] & b[346])^(a[61] & b[347])^(a[60] & b[348])^(a[59] & b[349])^(a[58] & b[350])^(a[57] & b[351])^(a[56] & b[352])^(a[55] & b[353])^(a[54] & b[354])^(a[53] & b[355])^(a[52] & b[356])^(a[51] & b[357])^(a[50] & b[358])^(a[49] & b[359])^(a[48] & b[360])^(a[47] & b[361])^(a[46] & b[362])^(a[45] & b[363])^(a[44] & b[364])^(a[43] & b[365])^(a[42] & b[366])^(a[41] & b[367])^(a[40] & b[368])^(a[39] & b[369])^(a[38] & b[370])^(a[37] & b[371])^(a[36] & b[372])^(a[35] & b[373])^(a[34] & b[374])^(a[33] & b[375])^(a[32] & b[376])^(a[31] & b[377])^(a[30] & b[378])^(a[29] & b[379])^(a[28] & b[380])^(a[27] & b[381])^(a[26] & b[382])^(a[25] & b[383])^(a[24] & b[384])^(a[23] & b[385])^(a[22] & b[386])^(a[21] & b[387])^(a[20] & b[388])^(a[19] & b[389])^(a[18] & b[390])^(a[17] & b[391])^(a[16] & b[392])^(a[15] & b[393])^(a[14] & b[394])^(a[13] & b[395])^(a[12] & b[396])^(a[11] & b[397])^(a[10] & b[398])^(a[9] & b[399])^(a[8] & b[400])^(a[7] & b[401])^(a[6] & b[402])^(a[5] & b[403])^(a[4] & b[404])^(a[3] & b[405])^(a[2] & b[406])^(a[1] & b[407])^(a[0] & b[408]);
assign y[409] = (a[408] & b[1])^(a[407] & b[2])^(a[406] & b[3])^(a[405] & b[4])^(a[404] & b[5])^(a[403] & b[6])^(a[402] & b[7])^(a[401] & b[8])^(a[400] & b[9])^(a[399] & b[10])^(a[398] & b[11])^(a[397] & b[12])^(a[396] & b[13])^(a[395] & b[14])^(a[394] & b[15])^(a[393] & b[16])^(a[392] & b[17])^(a[391] & b[18])^(a[390] & b[19])^(a[389] & b[20])^(a[388] & b[21])^(a[387] & b[22])^(a[386] & b[23])^(a[385] & b[24])^(a[384] & b[25])^(a[383] & b[26])^(a[382] & b[27])^(a[381] & b[28])^(a[380] & b[29])^(a[379] & b[30])^(a[378] & b[31])^(a[377] & b[32])^(a[376] & b[33])^(a[375] & b[34])^(a[374] & b[35])^(a[373] & b[36])^(a[372] & b[37])^(a[371] & b[38])^(a[370] & b[39])^(a[369] & b[40])^(a[368] & b[41])^(a[367] & b[42])^(a[366] & b[43])^(a[365] & b[44])^(a[364] & b[45])^(a[363] & b[46])^(a[362] & b[47])^(a[361] & b[48])^(a[360] & b[49])^(a[359] & b[50])^(a[358] & b[51])^(a[357] & b[52])^(a[356] & b[53])^(a[355] & b[54])^(a[354] & b[55])^(a[353] & b[56])^(a[352] & b[57])^(a[351] & b[58])^(a[350] & b[59])^(a[349] & b[60])^(a[348] & b[61])^(a[347] & b[62])^(a[346] & b[63])^(a[345] & b[64])^(a[344] & b[65])^(a[343] & b[66])^(a[342] & b[67])^(a[341] & b[68])^(a[340] & b[69])^(a[339] & b[70])^(a[338] & b[71])^(a[337] & b[72])^(a[336] & b[73])^(a[335] & b[74])^(a[334] & b[75])^(a[333] & b[76])^(a[332] & b[77])^(a[331] & b[78])^(a[330] & b[79])^(a[329] & b[80])^(a[328] & b[81])^(a[327] & b[82])^(a[326] & b[83])^(a[325] & b[84])^(a[324] & b[85])^(a[323] & b[86])^(a[322] & b[87])^(a[321] & b[88])^(a[320] & b[89])^(a[319] & b[90])^(a[318] & b[91])^(a[317] & b[92])^(a[316] & b[93])^(a[315] & b[94])^(a[314] & b[95])^(a[313] & b[96])^(a[312] & b[97])^(a[311] & b[98])^(a[310] & b[99])^(a[309] & b[100])^(a[308] & b[101])^(a[307] & b[102])^(a[306] & b[103])^(a[305] & b[104])^(a[304] & b[105])^(a[303] & b[106])^(a[302] & b[107])^(a[301] & b[108])^(a[300] & b[109])^(a[299] & b[110])^(a[298] & b[111])^(a[297] & b[112])^(a[296] & b[113])^(a[295] & b[114])^(a[294] & b[115])^(a[293] & b[116])^(a[292] & b[117])^(a[291] & b[118])^(a[290] & b[119])^(a[289] & b[120])^(a[288] & b[121])^(a[287] & b[122])^(a[286] & b[123])^(a[285] & b[124])^(a[284] & b[125])^(a[283] & b[126])^(a[282] & b[127])^(a[281] & b[128])^(a[280] & b[129])^(a[279] & b[130])^(a[278] & b[131])^(a[277] & b[132])^(a[276] & b[133])^(a[275] & b[134])^(a[274] & b[135])^(a[273] & b[136])^(a[272] & b[137])^(a[271] & b[138])^(a[270] & b[139])^(a[269] & b[140])^(a[268] & b[141])^(a[267] & b[142])^(a[266] & b[143])^(a[265] & b[144])^(a[264] & b[145])^(a[263] & b[146])^(a[262] & b[147])^(a[261] & b[148])^(a[260] & b[149])^(a[259] & b[150])^(a[258] & b[151])^(a[257] & b[152])^(a[256] & b[153])^(a[255] & b[154])^(a[254] & b[155])^(a[253] & b[156])^(a[252] & b[157])^(a[251] & b[158])^(a[250] & b[159])^(a[249] & b[160])^(a[248] & b[161])^(a[247] & b[162])^(a[246] & b[163])^(a[245] & b[164])^(a[244] & b[165])^(a[243] & b[166])^(a[242] & b[167])^(a[241] & b[168])^(a[240] & b[169])^(a[239] & b[170])^(a[238] & b[171])^(a[237] & b[172])^(a[236] & b[173])^(a[235] & b[174])^(a[234] & b[175])^(a[233] & b[176])^(a[232] & b[177])^(a[231] & b[178])^(a[230] & b[179])^(a[229] & b[180])^(a[228] & b[181])^(a[227] & b[182])^(a[226] & b[183])^(a[225] & b[184])^(a[224] & b[185])^(a[223] & b[186])^(a[222] & b[187])^(a[221] & b[188])^(a[220] & b[189])^(a[219] & b[190])^(a[218] & b[191])^(a[217] & b[192])^(a[216] & b[193])^(a[215] & b[194])^(a[214] & b[195])^(a[213] & b[196])^(a[212] & b[197])^(a[211] & b[198])^(a[210] & b[199])^(a[209] & b[200])^(a[208] & b[201])^(a[207] & b[202])^(a[206] & b[203])^(a[205] & b[204])^(a[204] & b[205])^(a[203] & b[206])^(a[202] & b[207])^(a[201] & b[208])^(a[200] & b[209])^(a[199] & b[210])^(a[198] & b[211])^(a[197] & b[212])^(a[196] & b[213])^(a[195] & b[214])^(a[194] & b[215])^(a[193] & b[216])^(a[192] & b[217])^(a[191] & b[218])^(a[190] & b[219])^(a[189] & b[220])^(a[188] & b[221])^(a[187] & b[222])^(a[186] & b[223])^(a[185] & b[224])^(a[184] & b[225])^(a[183] & b[226])^(a[182] & b[227])^(a[181] & b[228])^(a[180] & b[229])^(a[179] & b[230])^(a[178] & b[231])^(a[177] & b[232])^(a[176] & b[233])^(a[175] & b[234])^(a[174] & b[235])^(a[173] & b[236])^(a[172] & b[237])^(a[171] & b[238])^(a[170] & b[239])^(a[169] & b[240])^(a[168] & b[241])^(a[167] & b[242])^(a[166] & b[243])^(a[165] & b[244])^(a[164] & b[245])^(a[163] & b[246])^(a[162] & b[247])^(a[161] & b[248])^(a[160] & b[249])^(a[159] & b[250])^(a[158] & b[251])^(a[157] & b[252])^(a[156] & b[253])^(a[155] & b[254])^(a[154] & b[255])^(a[153] & b[256])^(a[152] & b[257])^(a[151] & b[258])^(a[150] & b[259])^(a[149] & b[260])^(a[148] & b[261])^(a[147] & b[262])^(a[146] & b[263])^(a[145] & b[264])^(a[144] & b[265])^(a[143] & b[266])^(a[142] & b[267])^(a[141] & b[268])^(a[140] & b[269])^(a[139] & b[270])^(a[138] & b[271])^(a[137] & b[272])^(a[136] & b[273])^(a[135] & b[274])^(a[134] & b[275])^(a[133] & b[276])^(a[132] & b[277])^(a[131] & b[278])^(a[130] & b[279])^(a[129] & b[280])^(a[128] & b[281])^(a[127] & b[282])^(a[126] & b[283])^(a[125] & b[284])^(a[124] & b[285])^(a[123] & b[286])^(a[122] & b[287])^(a[121] & b[288])^(a[120] & b[289])^(a[119] & b[290])^(a[118] & b[291])^(a[117] & b[292])^(a[116] & b[293])^(a[115] & b[294])^(a[114] & b[295])^(a[113] & b[296])^(a[112] & b[297])^(a[111] & b[298])^(a[110] & b[299])^(a[109] & b[300])^(a[108] & b[301])^(a[107] & b[302])^(a[106] & b[303])^(a[105] & b[304])^(a[104] & b[305])^(a[103] & b[306])^(a[102] & b[307])^(a[101] & b[308])^(a[100] & b[309])^(a[99] & b[310])^(a[98] & b[311])^(a[97] & b[312])^(a[96] & b[313])^(a[95] & b[314])^(a[94] & b[315])^(a[93] & b[316])^(a[92] & b[317])^(a[91] & b[318])^(a[90] & b[319])^(a[89] & b[320])^(a[88] & b[321])^(a[87] & b[322])^(a[86] & b[323])^(a[85] & b[324])^(a[84] & b[325])^(a[83] & b[326])^(a[82] & b[327])^(a[81] & b[328])^(a[80] & b[329])^(a[79] & b[330])^(a[78] & b[331])^(a[77] & b[332])^(a[76] & b[333])^(a[75] & b[334])^(a[74] & b[335])^(a[73] & b[336])^(a[72] & b[337])^(a[71] & b[338])^(a[70] & b[339])^(a[69] & b[340])^(a[68] & b[341])^(a[67] & b[342])^(a[66] & b[343])^(a[65] & b[344])^(a[64] & b[345])^(a[63] & b[346])^(a[62] & b[347])^(a[61] & b[348])^(a[60] & b[349])^(a[59] & b[350])^(a[58] & b[351])^(a[57] & b[352])^(a[56] & b[353])^(a[55] & b[354])^(a[54] & b[355])^(a[53] & b[356])^(a[52] & b[357])^(a[51] & b[358])^(a[50] & b[359])^(a[49] & b[360])^(a[48] & b[361])^(a[47] & b[362])^(a[46] & b[363])^(a[45] & b[364])^(a[44] & b[365])^(a[43] & b[366])^(a[42] & b[367])^(a[41] & b[368])^(a[40] & b[369])^(a[39] & b[370])^(a[38] & b[371])^(a[37] & b[372])^(a[36] & b[373])^(a[35] & b[374])^(a[34] & b[375])^(a[33] & b[376])^(a[32] & b[377])^(a[31] & b[378])^(a[30] & b[379])^(a[29] & b[380])^(a[28] & b[381])^(a[27] & b[382])^(a[26] & b[383])^(a[25] & b[384])^(a[24] & b[385])^(a[23] & b[386])^(a[22] & b[387])^(a[21] & b[388])^(a[20] & b[389])^(a[19] & b[390])^(a[18] & b[391])^(a[17] & b[392])^(a[16] & b[393])^(a[15] & b[394])^(a[14] & b[395])^(a[13] & b[396])^(a[12] & b[397])^(a[11] & b[398])^(a[10] & b[399])^(a[9] & b[400])^(a[8] & b[401])^(a[7] & b[402])^(a[6] & b[403])^(a[5] & b[404])^(a[4] & b[405])^(a[3] & b[406])^(a[2] & b[407])^(a[1] & b[408]);
assign y[410] = (a[408] & b[2])^(a[407] & b[3])^(a[406] & b[4])^(a[405] & b[5])^(a[404] & b[6])^(a[403] & b[7])^(a[402] & b[8])^(a[401] & b[9])^(a[400] & b[10])^(a[399] & b[11])^(a[398] & b[12])^(a[397] & b[13])^(a[396] & b[14])^(a[395] & b[15])^(a[394] & b[16])^(a[393] & b[17])^(a[392] & b[18])^(a[391] & b[19])^(a[390] & b[20])^(a[389] & b[21])^(a[388] & b[22])^(a[387] & b[23])^(a[386] & b[24])^(a[385] & b[25])^(a[384] & b[26])^(a[383] & b[27])^(a[382] & b[28])^(a[381] & b[29])^(a[380] & b[30])^(a[379] & b[31])^(a[378] & b[32])^(a[377] & b[33])^(a[376] & b[34])^(a[375] & b[35])^(a[374] & b[36])^(a[373] & b[37])^(a[372] & b[38])^(a[371] & b[39])^(a[370] & b[40])^(a[369] & b[41])^(a[368] & b[42])^(a[367] & b[43])^(a[366] & b[44])^(a[365] & b[45])^(a[364] & b[46])^(a[363] & b[47])^(a[362] & b[48])^(a[361] & b[49])^(a[360] & b[50])^(a[359] & b[51])^(a[358] & b[52])^(a[357] & b[53])^(a[356] & b[54])^(a[355] & b[55])^(a[354] & b[56])^(a[353] & b[57])^(a[352] & b[58])^(a[351] & b[59])^(a[350] & b[60])^(a[349] & b[61])^(a[348] & b[62])^(a[347] & b[63])^(a[346] & b[64])^(a[345] & b[65])^(a[344] & b[66])^(a[343] & b[67])^(a[342] & b[68])^(a[341] & b[69])^(a[340] & b[70])^(a[339] & b[71])^(a[338] & b[72])^(a[337] & b[73])^(a[336] & b[74])^(a[335] & b[75])^(a[334] & b[76])^(a[333] & b[77])^(a[332] & b[78])^(a[331] & b[79])^(a[330] & b[80])^(a[329] & b[81])^(a[328] & b[82])^(a[327] & b[83])^(a[326] & b[84])^(a[325] & b[85])^(a[324] & b[86])^(a[323] & b[87])^(a[322] & b[88])^(a[321] & b[89])^(a[320] & b[90])^(a[319] & b[91])^(a[318] & b[92])^(a[317] & b[93])^(a[316] & b[94])^(a[315] & b[95])^(a[314] & b[96])^(a[313] & b[97])^(a[312] & b[98])^(a[311] & b[99])^(a[310] & b[100])^(a[309] & b[101])^(a[308] & b[102])^(a[307] & b[103])^(a[306] & b[104])^(a[305] & b[105])^(a[304] & b[106])^(a[303] & b[107])^(a[302] & b[108])^(a[301] & b[109])^(a[300] & b[110])^(a[299] & b[111])^(a[298] & b[112])^(a[297] & b[113])^(a[296] & b[114])^(a[295] & b[115])^(a[294] & b[116])^(a[293] & b[117])^(a[292] & b[118])^(a[291] & b[119])^(a[290] & b[120])^(a[289] & b[121])^(a[288] & b[122])^(a[287] & b[123])^(a[286] & b[124])^(a[285] & b[125])^(a[284] & b[126])^(a[283] & b[127])^(a[282] & b[128])^(a[281] & b[129])^(a[280] & b[130])^(a[279] & b[131])^(a[278] & b[132])^(a[277] & b[133])^(a[276] & b[134])^(a[275] & b[135])^(a[274] & b[136])^(a[273] & b[137])^(a[272] & b[138])^(a[271] & b[139])^(a[270] & b[140])^(a[269] & b[141])^(a[268] & b[142])^(a[267] & b[143])^(a[266] & b[144])^(a[265] & b[145])^(a[264] & b[146])^(a[263] & b[147])^(a[262] & b[148])^(a[261] & b[149])^(a[260] & b[150])^(a[259] & b[151])^(a[258] & b[152])^(a[257] & b[153])^(a[256] & b[154])^(a[255] & b[155])^(a[254] & b[156])^(a[253] & b[157])^(a[252] & b[158])^(a[251] & b[159])^(a[250] & b[160])^(a[249] & b[161])^(a[248] & b[162])^(a[247] & b[163])^(a[246] & b[164])^(a[245] & b[165])^(a[244] & b[166])^(a[243] & b[167])^(a[242] & b[168])^(a[241] & b[169])^(a[240] & b[170])^(a[239] & b[171])^(a[238] & b[172])^(a[237] & b[173])^(a[236] & b[174])^(a[235] & b[175])^(a[234] & b[176])^(a[233] & b[177])^(a[232] & b[178])^(a[231] & b[179])^(a[230] & b[180])^(a[229] & b[181])^(a[228] & b[182])^(a[227] & b[183])^(a[226] & b[184])^(a[225] & b[185])^(a[224] & b[186])^(a[223] & b[187])^(a[222] & b[188])^(a[221] & b[189])^(a[220] & b[190])^(a[219] & b[191])^(a[218] & b[192])^(a[217] & b[193])^(a[216] & b[194])^(a[215] & b[195])^(a[214] & b[196])^(a[213] & b[197])^(a[212] & b[198])^(a[211] & b[199])^(a[210] & b[200])^(a[209] & b[201])^(a[208] & b[202])^(a[207] & b[203])^(a[206] & b[204])^(a[205] & b[205])^(a[204] & b[206])^(a[203] & b[207])^(a[202] & b[208])^(a[201] & b[209])^(a[200] & b[210])^(a[199] & b[211])^(a[198] & b[212])^(a[197] & b[213])^(a[196] & b[214])^(a[195] & b[215])^(a[194] & b[216])^(a[193] & b[217])^(a[192] & b[218])^(a[191] & b[219])^(a[190] & b[220])^(a[189] & b[221])^(a[188] & b[222])^(a[187] & b[223])^(a[186] & b[224])^(a[185] & b[225])^(a[184] & b[226])^(a[183] & b[227])^(a[182] & b[228])^(a[181] & b[229])^(a[180] & b[230])^(a[179] & b[231])^(a[178] & b[232])^(a[177] & b[233])^(a[176] & b[234])^(a[175] & b[235])^(a[174] & b[236])^(a[173] & b[237])^(a[172] & b[238])^(a[171] & b[239])^(a[170] & b[240])^(a[169] & b[241])^(a[168] & b[242])^(a[167] & b[243])^(a[166] & b[244])^(a[165] & b[245])^(a[164] & b[246])^(a[163] & b[247])^(a[162] & b[248])^(a[161] & b[249])^(a[160] & b[250])^(a[159] & b[251])^(a[158] & b[252])^(a[157] & b[253])^(a[156] & b[254])^(a[155] & b[255])^(a[154] & b[256])^(a[153] & b[257])^(a[152] & b[258])^(a[151] & b[259])^(a[150] & b[260])^(a[149] & b[261])^(a[148] & b[262])^(a[147] & b[263])^(a[146] & b[264])^(a[145] & b[265])^(a[144] & b[266])^(a[143] & b[267])^(a[142] & b[268])^(a[141] & b[269])^(a[140] & b[270])^(a[139] & b[271])^(a[138] & b[272])^(a[137] & b[273])^(a[136] & b[274])^(a[135] & b[275])^(a[134] & b[276])^(a[133] & b[277])^(a[132] & b[278])^(a[131] & b[279])^(a[130] & b[280])^(a[129] & b[281])^(a[128] & b[282])^(a[127] & b[283])^(a[126] & b[284])^(a[125] & b[285])^(a[124] & b[286])^(a[123] & b[287])^(a[122] & b[288])^(a[121] & b[289])^(a[120] & b[290])^(a[119] & b[291])^(a[118] & b[292])^(a[117] & b[293])^(a[116] & b[294])^(a[115] & b[295])^(a[114] & b[296])^(a[113] & b[297])^(a[112] & b[298])^(a[111] & b[299])^(a[110] & b[300])^(a[109] & b[301])^(a[108] & b[302])^(a[107] & b[303])^(a[106] & b[304])^(a[105] & b[305])^(a[104] & b[306])^(a[103] & b[307])^(a[102] & b[308])^(a[101] & b[309])^(a[100] & b[310])^(a[99] & b[311])^(a[98] & b[312])^(a[97] & b[313])^(a[96] & b[314])^(a[95] & b[315])^(a[94] & b[316])^(a[93] & b[317])^(a[92] & b[318])^(a[91] & b[319])^(a[90] & b[320])^(a[89] & b[321])^(a[88] & b[322])^(a[87] & b[323])^(a[86] & b[324])^(a[85] & b[325])^(a[84] & b[326])^(a[83] & b[327])^(a[82] & b[328])^(a[81] & b[329])^(a[80] & b[330])^(a[79] & b[331])^(a[78] & b[332])^(a[77] & b[333])^(a[76] & b[334])^(a[75] & b[335])^(a[74] & b[336])^(a[73] & b[337])^(a[72] & b[338])^(a[71] & b[339])^(a[70] & b[340])^(a[69] & b[341])^(a[68] & b[342])^(a[67] & b[343])^(a[66] & b[344])^(a[65] & b[345])^(a[64] & b[346])^(a[63] & b[347])^(a[62] & b[348])^(a[61] & b[349])^(a[60] & b[350])^(a[59] & b[351])^(a[58] & b[352])^(a[57] & b[353])^(a[56] & b[354])^(a[55] & b[355])^(a[54] & b[356])^(a[53] & b[357])^(a[52] & b[358])^(a[51] & b[359])^(a[50] & b[360])^(a[49] & b[361])^(a[48] & b[362])^(a[47] & b[363])^(a[46] & b[364])^(a[45] & b[365])^(a[44] & b[366])^(a[43] & b[367])^(a[42] & b[368])^(a[41] & b[369])^(a[40] & b[370])^(a[39] & b[371])^(a[38] & b[372])^(a[37] & b[373])^(a[36] & b[374])^(a[35] & b[375])^(a[34] & b[376])^(a[33] & b[377])^(a[32] & b[378])^(a[31] & b[379])^(a[30] & b[380])^(a[29] & b[381])^(a[28] & b[382])^(a[27] & b[383])^(a[26] & b[384])^(a[25] & b[385])^(a[24] & b[386])^(a[23] & b[387])^(a[22] & b[388])^(a[21] & b[389])^(a[20] & b[390])^(a[19] & b[391])^(a[18] & b[392])^(a[17] & b[393])^(a[16] & b[394])^(a[15] & b[395])^(a[14] & b[396])^(a[13] & b[397])^(a[12] & b[398])^(a[11] & b[399])^(a[10] & b[400])^(a[9] & b[401])^(a[8] & b[402])^(a[7] & b[403])^(a[6] & b[404])^(a[5] & b[405])^(a[4] & b[406])^(a[3] & b[407])^(a[2] & b[408]);
assign y[411] = (a[408] & b[3])^(a[407] & b[4])^(a[406] & b[5])^(a[405] & b[6])^(a[404] & b[7])^(a[403] & b[8])^(a[402] & b[9])^(a[401] & b[10])^(a[400] & b[11])^(a[399] & b[12])^(a[398] & b[13])^(a[397] & b[14])^(a[396] & b[15])^(a[395] & b[16])^(a[394] & b[17])^(a[393] & b[18])^(a[392] & b[19])^(a[391] & b[20])^(a[390] & b[21])^(a[389] & b[22])^(a[388] & b[23])^(a[387] & b[24])^(a[386] & b[25])^(a[385] & b[26])^(a[384] & b[27])^(a[383] & b[28])^(a[382] & b[29])^(a[381] & b[30])^(a[380] & b[31])^(a[379] & b[32])^(a[378] & b[33])^(a[377] & b[34])^(a[376] & b[35])^(a[375] & b[36])^(a[374] & b[37])^(a[373] & b[38])^(a[372] & b[39])^(a[371] & b[40])^(a[370] & b[41])^(a[369] & b[42])^(a[368] & b[43])^(a[367] & b[44])^(a[366] & b[45])^(a[365] & b[46])^(a[364] & b[47])^(a[363] & b[48])^(a[362] & b[49])^(a[361] & b[50])^(a[360] & b[51])^(a[359] & b[52])^(a[358] & b[53])^(a[357] & b[54])^(a[356] & b[55])^(a[355] & b[56])^(a[354] & b[57])^(a[353] & b[58])^(a[352] & b[59])^(a[351] & b[60])^(a[350] & b[61])^(a[349] & b[62])^(a[348] & b[63])^(a[347] & b[64])^(a[346] & b[65])^(a[345] & b[66])^(a[344] & b[67])^(a[343] & b[68])^(a[342] & b[69])^(a[341] & b[70])^(a[340] & b[71])^(a[339] & b[72])^(a[338] & b[73])^(a[337] & b[74])^(a[336] & b[75])^(a[335] & b[76])^(a[334] & b[77])^(a[333] & b[78])^(a[332] & b[79])^(a[331] & b[80])^(a[330] & b[81])^(a[329] & b[82])^(a[328] & b[83])^(a[327] & b[84])^(a[326] & b[85])^(a[325] & b[86])^(a[324] & b[87])^(a[323] & b[88])^(a[322] & b[89])^(a[321] & b[90])^(a[320] & b[91])^(a[319] & b[92])^(a[318] & b[93])^(a[317] & b[94])^(a[316] & b[95])^(a[315] & b[96])^(a[314] & b[97])^(a[313] & b[98])^(a[312] & b[99])^(a[311] & b[100])^(a[310] & b[101])^(a[309] & b[102])^(a[308] & b[103])^(a[307] & b[104])^(a[306] & b[105])^(a[305] & b[106])^(a[304] & b[107])^(a[303] & b[108])^(a[302] & b[109])^(a[301] & b[110])^(a[300] & b[111])^(a[299] & b[112])^(a[298] & b[113])^(a[297] & b[114])^(a[296] & b[115])^(a[295] & b[116])^(a[294] & b[117])^(a[293] & b[118])^(a[292] & b[119])^(a[291] & b[120])^(a[290] & b[121])^(a[289] & b[122])^(a[288] & b[123])^(a[287] & b[124])^(a[286] & b[125])^(a[285] & b[126])^(a[284] & b[127])^(a[283] & b[128])^(a[282] & b[129])^(a[281] & b[130])^(a[280] & b[131])^(a[279] & b[132])^(a[278] & b[133])^(a[277] & b[134])^(a[276] & b[135])^(a[275] & b[136])^(a[274] & b[137])^(a[273] & b[138])^(a[272] & b[139])^(a[271] & b[140])^(a[270] & b[141])^(a[269] & b[142])^(a[268] & b[143])^(a[267] & b[144])^(a[266] & b[145])^(a[265] & b[146])^(a[264] & b[147])^(a[263] & b[148])^(a[262] & b[149])^(a[261] & b[150])^(a[260] & b[151])^(a[259] & b[152])^(a[258] & b[153])^(a[257] & b[154])^(a[256] & b[155])^(a[255] & b[156])^(a[254] & b[157])^(a[253] & b[158])^(a[252] & b[159])^(a[251] & b[160])^(a[250] & b[161])^(a[249] & b[162])^(a[248] & b[163])^(a[247] & b[164])^(a[246] & b[165])^(a[245] & b[166])^(a[244] & b[167])^(a[243] & b[168])^(a[242] & b[169])^(a[241] & b[170])^(a[240] & b[171])^(a[239] & b[172])^(a[238] & b[173])^(a[237] & b[174])^(a[236] & b[175])^(a[235] & b[176])^(a[234] & b[177])^(a[233] & b[178])^(a[232] & b[179])^(a[231] & b[180])^(a[230] & b[181])^(a[229] & b[182])^(a[228] & b[183])^(a[227] & b[184])^(a[226] & b[185])^(a[225] & b[186])^(a[224] & b[187])^(a[223] & b[188])^(a[222] & b[189])^(a[221] & b[190])^(a[220] & b[191])^(a[219] & b[192])^(a[218] & b[193])^(a[217] & b[194])^(a[216] & b[195])^(a[215] & b[196])^(a[214] & b[197])^(a[213] & b[198])^(a[212] & b[199])^(a[211] & b[200])^(a[210] & b[201])^(a[209] & b[202])^(a[208] & b[203])^(a[207] & b[204])^(a[206] & b[205])^(a[205] & b[206])^(a[204] & b[207])^(a[203] & b[208])^(a[202] & b[209])^(a[201] & b[210])^(a[200] & b[211])^(a[199] & b[212])^(a[198] & b[213])^(a[197] & b[214])^(a[196] & b[215])^(a[195] & b[216])^(a[194] & b[217])^(a[193] & b[218])^(a[192] & b[219])^(a[191] & b[220])^(a[190] & b[221])^(a[189] & b[222])^(a[188] & b[223])^(a[187] & b[224])^(a[186] & b[225])^(a[185] & b[226])^(a[184] & b[227])^(a[183] & b[228])^(a[182] & b[229])^(a[181] & b[230])^(a[180] & b[231])^(a[179] & b[232])^(a[178] & b[233])^(a[177] & b[234])^(a[176] & b[235])^(a[175] & b[236])^(a[174] & b[237])^(a[173] & b[238])^(a[172] & b[239])^(a[171] & b[240])^(a[170] & b[241])^(a[169] & b[242])^(a[168] & b[243])^(a[167] & b[244])^(a[166] & b[245])^(a[165] & b[246])^(a[164] & b[247])^(a[163] & b[248])^(a[162] & b[249])^(a[161] & b[250])^(a[160] & b[251])^(a[159] & b[252])^(a[158] & b[253])^(a[157] & b[254])^(a[156] & b[255])^(a[155] & b[256])^(a[154] & b[257])^(a[153] & b[258])^(a[152] & b[259])^(a[151] & b[260])^(a[150] & b[261])^(a[149] & b[262])^(a[148] & b[263])^(a[147] & b[264])^(a[146] & b[265])^(a[145] & b[266])^(a[144] & b[267])^(a[143] & b[268])^(a[142] & b[269])^(a[141] & b[270])^(a[140] & b[271])^(a[139] & b[272])^(a[138] & b[273])^(a[137] & b[274])^(a[136] & b[275])^(a[135] & b[276])^(a[134] & b[277])^(a[133] & b[278])^(a[132] & b[279])^(a[131] & b[280])^(a[130] & b[281])^(a[129] & b[282])^(a[128] & b[283])^(a[127] & b[284])^(a[126] & b[285])^(a[125] & b[286])^(a[124] & b[287])^(a[123] & b[288])^(a[122] & b[289])^(a[121] & b[290])^(a[120] & b[291])^(a[119] & b[292])^(a[118] & b[293])^(a[117] & b[294])^(a[116] & b[295])^(a[115] & b[296])^(a[114] & b[297])^(a[113] & b[298])^(a[112] & b[299])^(a[111] & b[300])^(a[110] & b[301])^(a[109] & b[302])^(a[108] & b[303])^(a[107] & b[304])^(a[106] & b[305])^(a[105] & b[306])^(a[104] & b[307])^(a[103] & b[308])^(a[102] & b[309])^(a[101] & b[310])^(a[100] & b[311])^(a[99] & b[312])^(a[98] & b[313])^(a[97] & b[314])^(a[96] & b[315])^(a[95] & b[316])^(a[94] & b[317])^(a[93] & b[318])^(a[92] & b[319])^(a[91] & b[320])^(a[90] & b[321])^(a[89] & b[322])^(a[88] & b[323])^(a[87] & b[324])^(a[86] & b[325])^(a[85] & b[326])^(a[84] & b[327])^(a[83] & b[328])^(a[82] & b[329])^(a[81] & b[330])^(a[80] & b[331])^(a[79] & b[332])^(a[78] & b[333])^(a[77] & b[334])^(a[76] & b[335])^(a[75] & b[336])^(a[74] & b[337])^(a[73] & b[338])^(a[72] & b[339])^(a[71] & b[340])^(a[70] & b[341])^(a[69] & b[342])^(a[68] & b[343])^(a[67] & b[344])^(a[66] & b[345])^(a[65] & b[346])^(a[64] & b[347])^(a[63] & b[348])^(a[62] & b[349])^(a[61] & b[350])^(a[60] & b[351])^(a[59] & b[352])^(a[58] & b[353])^(a[57] & b[354])^(a[56] & b[355])^(a[55] & b[356])^(a[54] & b[357])^(a[53] & b[358])^(a[52] & b[359])^(a[51] & b[360])^(a[50] & b[361])^(a[49] & b[362])^(a[48] & b[363])^(a[47] & b[364])^(a[46] & b[365])^(a[45] & b[366])^(a[44] & b[367])^(a[43] & b[368])^(a[42] & b[369])^(a[41] & b[370])^(a[40] & b[371])^(a[39] & b[372])^(a[38] & b[373])^(a[37] & b[374])^(a[36] & b[375])^(a[35] & b[376])^(a[34] & b[377])^(a[33] & b[378])^(a[32] & b[379])^(a[31] & b[380])^(a[30] & b[381])^(a[29] & b[382])^(a[28] & b[383])^(a[27] & b[384])^(a[26] & b[385])^(a[25] & b[386])^(a[24] & b[387])^(a[23] & b[388])^(a[22] & b[389])^(a[21] & b[390])^(a[20] & b[391])^(a[19] & b[392])^(a[18] & b[393])^(a[17] & b[394])^(a[16] & b[395])^(a[15] & b[396])^(a[14] & b[397])^(a[13] & b[398])^(a[12] & b[399])^(a[11] & b[400])^(a[10] & b[401])^(a[9] & b[402])^(a[8] & b[403])^(a[7] & b[404])^(a[6] & b[405])^(a[5] & b[406])^(a[4] & b[407])^(a[3] & b[408]);
assign y[412] = (a[408] & b[4])^(a[407] & b[5])^(a[406] & b[6])^(a[405] & b[7])^(a[404] & b[8])^(a[403] & b[9])^(a[402] & b[10])^(a[401] & b[11])^(a[400] & b[12])^(a[399] & b[13])^(a[398] & b[14])^(a[397] & b[15])^(a[396] & b[16])^(a[395] & b[17])^(a[394] & b[18])^(a[393] & b[19])^(a[392] & b[20])^(a[391] & b[21])^(a[390] & b[22])^(a[389] & b[23])^(a[388] & b[24])^(a[387] & b[25])^(a[386] & b[26])^(a[385] & b[27])^(a[384] & b[28])^(a[383] & b[29])^(a[382] & b[30])^(a[381] & b[31])^(a[380] & b[32])^(a[379] & b[33])^(a[378] & b[34])^(a[377] & b[35])^(a[376] & b[36])^(a[375] & b[37])^(a[374] & b[38])^(a[373] & b[39])^(a[372] & b[40])^(a[371] & b[41])^(a[370] & b[42])^(a[369] & b[43])^(a[368] & b[44])^(a[367] & b[45])^(a[366] & b[46])^(a[365] & b[47])^(a[364] & b[48])^(a[363] & b[49])^(a[362] & b[50])^(a[361] & b[51])^(a[360] & b[52])^(a[359] & b[53])^(a[358] & b[54])^(a[357] & b[55])^(a[356] & b[56])^(a[355] & b[57])^(a[354] & b[58])^(a[353] & b[59])^(a[352] & b[60])^(a[351] & b[61])^(a[350] & b[62])^(a[349] & b[63])^(a[348] & b[64])^(a[347] & b[65])^(a[346] & b[66])^(a[345] & b[67])^(a[344] & b[68])^(a[343] & b[69])^(a[342] & b[70])^(a[341] & b[71])^(a[340] & b[72])^(a[339] & b[73])^(a[338] & b[74])^(a[337] & b[75])^(a[336] & b[76])^(a[335] & b[77])^(a[334] & b[78])^(a[333] & b[79])^(a[332] & b[80])^(a[331] & b[81])^(a[330] & b[82])^(a[329] & b[83])^(a[328] & b[84])^(a[327] & b[85])^(a[326] & b[86])^(a[325] & b[87])^(a[324] & b[88])^(a[323] & b[89])^(a[322] & b[90])^(a[321] & b[91])^(a[320] & b[92])^(a[319] & b[93])^(a[318] & b[94])^(a[317] & b[95])^(a[316] & b[96])^(a[315] & b[97])^(a[314] & b[98])^(a[313] & b[99])^(a[312] & b[100])^(a[311] & b[101])^(a[310] & b[102])^(a[309] & b[103])^(a[308] & b[104])^(a[307] & b[105])^(a[306] & b[106])^(a[305] & b[107])^(a[304] & b[108])^(a[303] & b[109])^(a[302] & b[110])^(a[301] & b[111])^(a[300] & b[112])^(a[299] & b[113])^(a[298] & b[114])^(a[297] & b[115])^(a[296] & b[116])^(a[295] & b[117])^(a[294] & b[118])^(a[293] & b[119])^(a[292] & b[120])^(a[291] & b[121])^(a[290] & b[122])^(a[289] & b[123])^(a[288] & b[124])^(a[287] & b[125])^(a[286] & b[126])^(a[285] & b[127])^(a[284] & b[128])^(a[283] & b[129])^(a[282] & b[130])^(a[281] & b[131])^(a[280] & b[132])^(a[279] & b[133])^(a[278] & b[134])^(a[277] & b[135])^(a[276] & b[136])^(a[275] & b[137])^(a[274] & b[138])^(a[273] & b[139])^(a[272] & b[140])^(a[271] & b[141])^(a[270] & b[142])^(a[269] & b[143])^(a[268] & b[144])^(a[267] & b[145])^(a[266] & b[146])^(a[265] & b[147])^(a[264] & b[148])^(a[263] & b[149])^(a[262] & b[150])^(a[261] & b[151])^(a[260] & b[152])^(a[259] & b[153])^(a[258] & b[154])^(a[257] & b[155])^(a[256] & b[156])^(a[255] & b[157])^(a[254] & b[158])^(a[253] & b[159])^(a[252] & b[160])^(a[251] & b[161])^(a[250] & b[162])^(a[249] & b[163])^(a[248] & b[164])^(a[247] & b[165])^(a[246] & b[166])^(a[245] & b[167])^(a[244] & b[168])^(a[243] & b[169])^(a[242] & b[170])^(a[241] & b[171])^(a[240] & b[172])^(a[239] & b[173])^(a[238] & b[174])^(a[237] & b[175])^(a[236] & b[176])^(a[235] & b[177])^(a[234] & b[178])^(a[233] & b[179])^(a[232] & b[180])^(a[231] & b[181])^(a[230] & b[182])^(a[229] & b[183])^(a[228] & b[184])^(a[227] & b[185])^(a[226] & b[186])^(a[225] & b[187])^(a[224] & b[188])^(a[223] & b[189])^(a[222] & b[190])^(a[221] & b[191])^(a[220] & b[192])^(a[219] & b[193])^(a[218] & b[194])^(a[217] & b[195])^(a[216] & b[196])^(a[215] & b[197])^(a[214] & b[198])^(a[213] & b[199])^(a[212] & b[200])^(a[211] & b[201])^(a[210] & b[202])^(a[209] & b[203])^(a[208] & b[204])^(a[207] & b[205])^(a[206] & b[206])^(a[205] & b[207])^(a[204] & b[208])^(a[203] & b[209])^(a[202] & b[210])^(a[201] & b[211])^(a[200] & b[212])^(a[199] & b[213])^(a[198] & b[214])^(a[197] & b[215])^(a[196] & b[216])^(a[195] & b[217])^(a[194] & b[218])^(a[193] & b[219])^(a[192] & b[220])^(a[191] & b[221])^(a[190] & b[222])^(a[189] & b[223])^(a[188] & b[224])^(a[187] & b[225])^(a[186] & b[226])^(a[185] & b[227])^(a[184] & b[228])^(a[183] & b[229])^(a[182] & b[230])^(a[181] & b[231])^(a[180] & b[232])^(a[179] & b[233])^(a[178] & b[234])^(a[177] & b[235])^(a[176] & b[236])^(a[175] & b[237])^(a[174] & b[238])^(a[173] & b[239])^(a[172] & b[240])^(a[171] & b[241])^(a[170] & b[242])^(a[169] & b[243])^(a[168] & b[244])^(a[167] & b[245])^(a[166] & b[246])^(a[165] & b[247])^(a[164] & b[248])^(a[163] & b[249])^(a[162] & b[250])^(a[161] & b[251])^(a[160] & b[252])^(a[159] & b[253])^(a[158] & b[254])^(a[157] & b[255])^(a[156] & b[256])^(a[155] & b[257])^(a[154] & b[258])^(a[153] & b[259])^(a[152] & b[260])^(a[151] & b[261])^(a[150] & b[262])^(a[149] & b[263])^(a[148] & b[264])^(a[147] & b[265])^(a[146] & b[266])^(a[145] & b[267])^(a[144] & b[268])^(a[143] & b[269])^(a[142] & b[270])^(a[141] & b[271])^(a[140] & b[272])^(a[139] & b[273])^(a[138] & b[274])^(a[137] & b[275])^(a[136] & b[276])^(a[135] & b[277])^(a[134] & b[278])^(a[133] & b[279])^(a[132] & b[280])^(a[131] & b[281])^(a[130] & b[282])^(a[129] & b[283])^(a[128] & b[284])^(a[127] & b[285])^(a[126] & b[286])^(a[125] & b[287])^(a[124] & b[288])^(a[123] & b[289])^(a[122] & b[290])^(a[121] & b[291])^(a[120] & b[292])^(a[119] & b[293])^(a[118] & b[294])^(a[117] & b[295])^(a[116] & b[296])^(a[115] & b[297])^(a[114] & b[298])^(a[113] & b[299])^(a[112] & b[300])^(a[111] & b[301])^(a[110] & b[302])^(a[109] & b[303])^(a[108] & b[304])^(a[107] & b[305])^(a[106] & b[306])^(a[105] & b[307])^(a[104] & b[308])^(a[103] & b[309])^(a[102] & b[310])^(a[101] & b[311])^(a[100] & b[312])^(a[99] & b[313])^(a[98] & b[314])^(a[97] & b[315])^(a[96] & b[316])^(a[95] & b[317])^(a[94] & b[318])^(a[93] & b[319])^(a[92] & b[320])^(a[91] & b[321])^(a[90] & b[322])^(a[89] & b[323])^(a[88] & b[324])^(a[87] & b[325])^(a[86] & b[326])^(a[85] & b[327])^(a[84] & b[328])^(a[83] & b[329])^(a[82] & b[330])^(a[81] & b[331])^(a[80] & b[332])^(a[79] & b[333])^(a[78] & b[334])^(a[77] & b[335])^(a[76] & b[336])^(a[75] & b[337])^(a[74] & b[338])^(a[73] & b[339])^(a[72] & b[340])^(a[71] & b[341])^(a[70] & b[342])^(a[69] & b[343])^(a[68] & b[344])^(a[67] & b[345])^(a[66] & b[346])^(a[65] & b[347])^(a[64] & b[348])^(a[63] & b[349])^(a[62] & b[350])^(a[61] & b[351])^(a[60] & b[352])^(a[59] & b[353])^(a[58] & b[354])^(a[57] & b[355])^(a[56] & b[356])^(a[55] & b[357])^(a[54] & b[358])^(a[53] & b[359])^(a[52] & b[360])^(a[51] & b[361])^(a[50] & b[362])^(a[49] & b[363])^(a[48] & b[364])^(a[47] & b[365])^(a[46] & b[366])^(a[45] & b[367])^(a[44] & b[368])^(a[43] & b[369])^(a[42] & b[370])^(a[41] & b[371])^(a[40] & b[372])^(a[39] & b[373])^(a[38] & b[374])^(a[37] & b[375])^(a[36] & b[376])^(a[35] & b[377])^(a[34] & b[378])^(a[33] & b[379])^(a[32] & b[380])^(a[31] & b[381])^(a[30] & b[382])^(a[29] & b[383])^(a[28] & b[384])^(a[27] & b[385])^(a[26] & b[386])^(a[25] & b[387])^(a[24] & b[388])^(a[23] & b[389])^(a[22] & b[390])^(a[21] & b[391])^(a[20] & b[392])^(a[19] & b[393])^(a[18] & b[394])^(a[17] & b[395])^(a[16] & b[396])^(a[15] & b[397])^(a[14] & b[398])^(a[13] & b[399])^(a[12] & b[400])^(a[11] & b[401])^(a[10] & b[402])^(a[9] & b[403])^(a[8] & b[404])^(a[7] & b[405])^(a[6] & b[406])^(a[5] & b[407])^(a[4] & b[408]);
assign y[413] = (a[408] & b[5])^(a[407] & b[6])^(a[406] & b[7])^(a[405] & b[8])^(a[404] & b[9])^(a[403] & b[10])^(a[402] & b[11])^(a[401] & b[12])^(a[400] & b[13])^(a[399] & b[14])^(a[398] & b[15])^(a[397] & b[16])^(a[396] & b[17])^(a[395] & b[18])^(a[394] & b[19])^(a[393] & b[20])^(a[392] & b[21])^(a[391] & b[22])^(a[390] & b[23])^(a[389] & b[24])^(a[388] & b[25])^(a[387] & b[26])^(a[386] & b[27])^(a[385] & b[28])^(a[384] & b[29])^(a[383] & b[30])^(a[382] & b[31])^(a[381] & b[32])^(a[380] & b[33])^(a[379] & b[34])^(a[378] & b[35])^(a[377] & b[36])^(a[376] & b[37])^(a[375] & b[38])^(a[374] & b[39])^(a[373] & b[40])^(a[372] & b[41])^(a[371] & b[42])^(a[370] & b[43])^(a[369] & b[44])^(a[368] & b[45])^(a[367] & b[46])^(a[366] & b[47])^(a[365] & b[48])^(a[364] & b[49])^(a[363] & b[50])^(a[362] & b[51])^(a[361] & b[52])^(a[360] & b[53])^(a[359] & b[54])^(a[358] & b[55])^(a[357] & b[56])^(a[356] & b[57])^(a[355] & b[58])^(a[354] & b[59])^(a[353] & b[60])^(a[352] & b[61])^(a[351] & b[62])^(a[350] & b[63])^(a[349] & b[64])^(a[348] & b[65])^(a[347] & b[66])^(a[346] & b[67])^(a[345] & b[68])^(a[344] & b[69])^(a[343] & b[70])^(a[342] & b[71])^(a[341] & b[72])^(a[340] & b[73])^(a[339] & b[74])^(a[338] & b[75])^(a[337] & b[76])^(a[336] & b[77])^(a[335] & b[78])^(a[334] & b[79])^(a[333] & b[80])^(a[332] & b[81])^(a[331] & b[82])^(a[330] & b[83])^(a[329] & b[84])^(a[328] & b[85])^(a[327] & b[86])^(a[326] & b[87])^(a[325] & b[88])^(a[324] & b[89])^(a[323] & b[90])^(a[322] & b[91])^(a[321] & b[92])^(a[320] & b[93])^(a[319] & b[94])^(a[318] & b[95])^(a[317] & b[96])^(a[316] & b[97])^(a[315] & b[98])^(a[314] & b[99])^(a[313] & b[100])^(a[312] & b[101])^(a[311] & b[102])^(a[310] & b[103])^(a[309] & b[104])^(a[308] & b[105])^(a[307] & b[106])^(a[306] & b[107])^(a[305] & b[108])^(a[304] & b[109])^(a[303] & b[110])^(a[302] & b[111])^(a[301] & b[112])^(a[300] & b[113])^(a[299] & b[114])^(a[298] & b[115])^(a[297] & b[116])^(a[296] & b[117])^(a[295] & b[118])^(a[294] & b[119])^(a[293] & b[120])^(a[292] & b[121])^(a[291] & b[122])^(a[290] & b[123])^(a[289] & b[124])^(a[288] & b[125])^(a[287] & b[126])^(a[286] & b[127])^(a[285] & b[128])^(a[284] & b[129])^(a[283] & b[130])^(a[282] & b[131])^(a[281] & b[132])^(a[280] & b[133])^(a[279] & b[134])^(a[278] & b[135])^(a[277] & b[136])^(a[276] & b[137])^(a[275] & b[138])^(a[274] & b[139])^(a[273] & b[140])^(a[272] & b[141])^(a[271] & b[142])^(a[270] & b[143])^(a[269] & b[144])^(a[268] & b[145])^(a[267] & b[146])^(a[266] & b[147])^(a[265] & b[148])^(a[264] & b[149])^(a[263] & b[150])^(a[262] & b[151])^(a[261] & b[152])^(a[260] & b[153])^(a[259] & b[154])^(a[258] & b[155])^(a[257] & b[156])^(a[256] & b[157])^(a[255] & b[158])^(a[254] & b[159])^(a[253] & b[160])^(a[252] & b[161])^(a[251] & b[162])^(a[250] & b[163])^(a[249] & b[164])^(a[248] & b[165])^(a[247] & b[166])^(a[246] & b[167])^(a[245] & b[168])^(a[244] & b[169])^(a[243] & b[170])^(a[242] & b[171])^(a[241] & b[172])^(a[240] & b[173])^(a[239] & b[174])^(a[238] & b[175])^(a[237] & b[176])^(a[236] & b[177])^(a[235] & b[178])^(a[234] & b[179])^(a[233] & b[180])^(a[232] & b[181])^(a[231] & b[182])^(a[230] & b[183])^(a[229] & b[184])^(a[228] & b[185])^(a[227] & b[186])^(a[226] & b[187])^(a[225] & b[188])^(a[224] & b[189])^(a[223] & b[190])^(a[222] & b[191])^(a[221] & b[192])^(a[220] & b[193])^(a[219] & b[194])^(a[218] & b[195])^(a[217] & b[196])^(a[216] & b[197])^(a[215] & b[198])^(a[214] & b[199])^(a[213] & b[200])^(a[212] & b[201])^(a[211] & b[202])^(a[210] & b[203])^(a[209] & b[204])^(a[208] & b[205])^(a[207] & b[206])^(a[206] & b[207])^(a[205] & b[208])^(a[204] & b[209])^(a[203] & b[210])^(a[202] & b[211])^(a[201] & b[212])^(a[200] & b[213])^(a[199] & b[214])^(a[198] & b[215])^(a[197] & b[216])^(a[196] & b[217])^(a[195] & b[218])^(a[194] & b[219])^(a[193] & b[220])^(a[192] & b[221])^(a[191] & b[222])^(a[190] & b[223])^(a[189] & b[224])^(a[188] & b[225])^(a[187] & b[226])^(a[186] & b[227])^(a[185] & b[228])^(a[184] & b[229])^(a[183] & b[230])^(a[182] & b[231])^(a[181] & b[232])^(a[180] & b[233])^(a[179] & b[234])^(a[178] & b[235])^(a[177] & b[236])^(a[176] & b[237])^(a[175] & b[238])^(a[174] & b[239])^(a[173] & b[240])^(a[172] & b[241])^(a[171] & b[242])^(a[170] & b[243])^(a[169] & b[244])^(a[168] & b[245])^(a[167] & b[246])^(a[166] & b[247])^(a[165] & b[248])^(a[164] & b[249])^(a[163] & b[250])^(a[162] & b[251])^(a[161] & b[252])^(a[160] & b[253])^(a[159] & b[254])^(a[158] & b[255])^(a[157] & b[256])^(a[156] & b[257])^(a[155] & b[258])^(a[154] & b[259])^(a[153] & b[260])^(a[152] & b[261])^(a[151] & b[262])^(a[150] & b[263])^(a[149] & b[264])^(a[148] & b[265])^(a[147] & b[266])^(a[146] & b[267])^(a[145] & b[268])^(a[144] & b[269])^(a[143] & b[270])^(a[142] & b[271])^(a[141] & b[272])^(a[140] & b[273])^(a[139] & b[274])^(a[138] & b[275])^(a[137] & b[276])^(a[136] & b[277])^(a[135] & b[278])^(a[134] & b[279])^(a[133] & b[280])^(a[132] & b[281])^(a[131] & b[282])^(a[130] & b[283])^(a[129] & b[284])^(a[128] & b[285])^(a[127] & b[286])^(a[126] & b[287])^(a[125] & b[288])^(a[124] & b[289])^(a[123] & b[290])^(a[122] & b[291])^(a[121] & b[292])^(a[120] & b[293])^(a[119] & b[294])^(a[118] & b[295])^(a[117] & b[296])^(a[116] & b[297])^(a[115] & b[298])^(a[114] & b[299])^(a[113] & b[300])^(a[112] & b[301])^(a[111] & b[302])^(a[110] & b[303])^(a[109] & b[304])^(a[108] & b[305])^(a[107] & b[306])^(a[106] & b[307])^(a[105] & b[308])^(a[104] & b[309])^(a[103] & b[310])^(a[102] & b[311])^(a[101] & b[312])^(a[100] & b[313])^(a[99] & b[314])^(a[98] & b[315])^(a[97] & b[316])^(a[96] & b[317])^(a[95] & b[318])^(a[94] & b[319])^(a[93] & b[320])^(a[92] & b[321])^(a[91] & b[322])^(a[90] & b[323])^(a[89] & b[324])^(a[88] & b[325])^(a[87] & b[326])^(a[86] & b[327])^(a[85] & b[328])^(a[84] & b[329])^(a[83] & b[330])^(a[82] & b[331])^(a[81] & b[332])^(a[80] & b[333])^(a[79] & b[334])^(a[78] & b[335])^(a[77] & b[336])^(a[76] & b[337])^(a[75] & b[338])^(a[74] & b[339])^(a[73] & b[340])^(a[72] & b[341])^(a[71] & b[342])^(a[70] & b[343])^(a[69] & b[344])^(a[68] & b[345])^(a[67] & b[346])^(a[66] & b[347])^(a[65] & b[348])^(a[64] & b[349])^(a[63] & b[350])^(a[62] & b[351])^(a[61] & b[352])^(a[60] & b[353])^(a[59] & b[354])^(a[58] & b[355])^(a[57] & b[356])^(a[56] & b[357])^(a[55] & b[358])^(a[54] & b[359])^(a[53] & b[360])^(a[52] & b[361])^(a[51] & b[362])^(a[50] & b[363])^(a[49] & b[364])^(a[48] & b[365])^(a[47] & b[366])^(a[46] & b[367])^(a[45] & b[368])^(a[44] & b[369])^(a[43] & b[370])^(a[42] & b[371])^(a[41] & b[372])^(a[40] & b[373])^(a[39] & b[374])^(a[38] & b[375])^(a[37] & b[376])^(a[36] & b[377])^(a[35] & b[378])^(a[34] & b[379])^(a[33] & b[380])^(a[32] & b[381])^(a[31] & b[382])^(a[30] & b[383])^(a[29] & b[384])^(a[28] & b[385])^(a[27] & b[386])^(a[26] & b[387])^(a[25] & b[388])^(a[24] & b[389])^(a[23] & b[390])^(a[22] & b[391])^(a[21] & b[392])^(a[20] & b[393])^(a[19] & b[394])^(a[18] & b[395])^(a[17] & b[396])^(a[16] & b[397])^(a[15] & b[398])^(a[14] & b[399])^(a[13] & b[400])^(a[12] & b[401])^(a[11] & b[402])^(a[10] & b[403])^(a[9] & b[404])^(a[8] & b[405])^(a[7] & b[406])^(a[6] & b[407])^(a[5] & b[408]);
assign y[414] = (a[408] & b[6])^(a[407] & b[7])^(a[406] & b[8])^(a[405] & b[9])^(a[404] & b[10])^(a[403] & b[11])^(a[402] & b[12])^(a[401] & b[13])^(a[400] & b[14])^(a[399] & b[15])^(a[398] & b[16])^(a[397] & b[17])^(a[396] & b[18])^(a[395] & b[19])^(a[394] & b[20])^(a[393] & b[21])^(a[392] & b[22])^(a[391] & b[23])^(a[390] & b[24])^(a[389] & b[25])^(a[388] & b[26])^(a[387] & b[27])^(a[386] & b[28])^(a[385] & b[29])^(a[384] & b[30])^(a[383] & b[31])^(a[382] & b[32])^(a[381] & b[33])^(a[380] & b[34])^(a[379] & b[35])^(a[378] & b[36])^(a[377] & b[37])^(a[376] & b[38])^(a[375] & b[39])^(a[374] & b[40])^(a[373] & b[41])^(a[372] & b[42])^(a[371] & b[43])^(a[370] & b[44])^(a[369] & b[45])^(a[368] & b[46])^(a[367] & b[47])^(a[366] & b[48])^(a[365] & b[49])^(a[364] & b[50])^(a[363] & b[51])^(a[362] & b[52])^(a[361] & b[53])^(a[360] & b[54])^(a[359] & b[55])^(a[358] & b[56])^(a[357] & b[57])^(a[356] & b[58])^(a[355] & b[59])^(a[354] & b[60])^(a[353] & b[61])^(a[352] & b[62])^(a[351] & b[63])^(a[350] & b[64])^(a[349] & b[65])^(a[348] & b[66])^(a[347] & b[67])^(a[346] & b[68])^(a[345] & b[69])^(a[344] & b[70])^(a[343] & b[71])^(a[342] & b[72])^(a[341] & b[73])^(a[340] & b[74])^(a[339] & b[75])^(a[338] & b[76])^(a[337] & b[77])^(a[336] & b[78])^(a[335] & b[79])^(a[334] & b[80])^(a[333] & b[81])^(a[332] & b[82])^(a[331] & b[83])^(a[330] & b[84])^(a[329] & b[85])^(a[328] & b[86])^(a[327] & b[87])^(a[326] & b[88])^(a[325] & b[89])^(a[324] & b[90])^(a[323] & b[91])^(a[322] & b[92])^(a[321] & b[93])^(a[320] & b[94])^(a[319] & b[95])^(a[318] & b[96])^(a[317] & b[97])^(a[316] & b[98])^(a[315] & b[99])^(a[314] & b[100])^(a[313] & b[101])^(a[312] & b[102])^(a[311] & b[103])^(a[310] & b[104])^(a[309] & b[105])^(a[308] & b[106])^(a[307] & b[107])^(a[306] & b[108])^(a[305] & b[109])^(a[304] & b[110])^(a[303] & b[111])^(a[302] & b[112])^(a[301] & b[113])^(a[300] & b[114])^(a[299] & b[115])^(a[298] & b[116])^(a[297] & b[117])^(a[296] & b[118])^(a[295] & b[119])^(a[294] & b[120])^(a[293] & b[121])^(a[292] & b[122])^(a[291] & b[123])^(a[290] & b[124])^(a[289] & b[125])^(a[288] & b[126])^(a[287] & b[127])^(a[286] & b[128])^(a[285] & b[129])^(a[284] & b[130])^(a[283] & b[131])^(a[282] & b[132])^(a[281] & b[133])^(a[280] & b[134])^(a[279] & b[135])^(a[278] & b[136])^(a[277] & b[137])^(a[276] & b[138])^(a[275] & b[139])^(a[274] & b[140])^(a[273] & b[141])^(a[272] & b[142])^(a[271] & b[143])^(a[270] & b[144])^(a[269] & b[145])^(a[268] & b[146])^(a[267] & b[147])^(a[266] & b[148])^(a[265] & b[149])^(a[264] & b[150])^(a[263] & b[151])^(a[262] & b[152])^(a[261] & b[153])^(a[260] & b[154])^(a[259] & b[155])^(a[258] & b[156])^(a[257] & b[157])^(a[256] & b[158])^(a[255] & b[159])^(a[254] & b[160])^(a[253] & b[161])^(a[252] & b[162])^(a[251] & b[163])^(a[250] & b[164])^(a[249] & b[165])^(a[248] & b[166])^(a[247] & b[167])^(a[246] & b[168])^(a[245] & b[169])^(a[244] & b[170])^(a[243] & b[171])^(a[242] & b[172])^(a[241] & b[173])^(a[240] & b[174])^(a[239] & b[175])^(a[238] & b[176])^(a[237] & b[177])^(a[236] & b[178])^(a[235] & b[179])^(a[234] & b[180])^(a[233] & b[181])^(a[232] & b[182])^(a[231] & b[183])^(a[230] & b[184])^(a[229] & b[185])^(a[228] & b[186])^(a[227] & b[187])^(a[226] & b[188])^(a[225] & b[189])^(a[224] & b[190])^(a[223] & b[191])^(a[222] & b[192])^(a[221] & b[193])^(a[220] & b[194])^(a[219] & b[195])^(a[218] & b[196])^(a[217] & b[197])^(a[216] & b[198])^(a[215] & b[199])^(a[214] & b[200])^(a[213] & b[201])^(a[212] & b[202])^(a[211] & b[203])^(a[210] & b[204])^(a[209] & b[205])^(a[208] & b[206])^(a[207] & b[207])^(a[206] & b[208])^(a[205] & b[209])^(a[204] & b[210])^(a[203] & b[211])^(a[202] & b[212])^(a[201] & b[213])^(a[200] & b[214])^(a[199] & b[215])^(a[198] & b[216])^(a[197] & b[217])^(a[196] & b[218])^(a[195] & b[219])^(a[194] & b[220])^(a[193] & b[221])^(a[192] & b[222])^(a[191] & b[223])^(a[190] & b[224])^(a[189] & b[225])^(a[188] & b[226])^(a[187] & b[227])^(a[186] & b[228])^(a[185] & b[229])^(a[184] & b[230])^(a[183] & b[231])^(a[182] & b[232])^(a[181] & b[233])^(a[180] & b[234])^(a[179] & b[235])^(a[178] & b[236])^(a[177] & b[237])^(a[176] & b[238])^(a[175] & b[239])^(a[174] & b[240])^(a[173] & b[241])^(a[172] & b[242])^(a[171] & b[243])^(a[170] & b[244])^(a[169] & b[245])^(a[168] & b[246])^(a[167] & b[247])^(a[166] & b[248])^(a[165] & b[249])^(a[164] & b[250])^(a[163] & b[251])^(a[162] & b[252])^(a[161] & b[253])^(a[160] & b[254])^(a[159] & b[255])^(a[158] & b[256])^(a[157] & b[257])^(a[156] & b[258])^(a[155] & b[259])^(a[154] & b[260])^(a[153] & b[261])^(a[152] & b[262])^(a[151] & b[263])^(a[150] & b[264])^(a[149] & b[265])^(a[148] & b[266])^(a[147] & b[267])^(a[146] & b[268])^(a[145] & b[269])^(a[144] & b[270])^(a[143] & b[271])^(a[142] & b[272])^(a[141] & b[273])^(a[140] & b[274])^(a[139] & b[275])^(a[138] & b[276])^(a[137] & b[277])^(a[136] & b[278])^(a[135] & b[279])^(a[134] & b[280])^(a[133] & b[281])^(a[132] & b[282])^(a[131] & b[283])^(a[130] & b[284])^(a[129] & b[285])^(a[128] & b[286])^(a[127] & b[287])^(a[126] & b[288])^(a[125] & b[289])^(a[124] & b[290])^(a[123] & b[291])^(a[122] & b[292])^(a[121] & b[293])^(a[120] & b[294])^(a[119] & b[295])^(a[118] & b[296])^(a[117] & b[297])^(a[116] & b[298])^(a[115] & b[299])^(a[114] & b[300])^(a[113] & b[301])^(a[112] & b[302])^(a[111] & b[303])^(a[110] & b[304])^(a[109] & b[305])^(a[108] & b[306])^(a[107] & b[307])^(a[106] & b[308])^(a[105] & b[309])^(a[104] & b[310])^(a[103] & b[311])^(a[102] & b[312])^(a[101] & b[313])^(a[100] & b[314])^(a[99] & b[315])^(a[98] & b[316])^(a[97] & b[317])^(a[96] & b[318])^(a[95] & b[319])^(a[94] & b[320])^(a[93] & b[321])^(a[92] & b[322])^(a[91] & b[323])^(a[90] & b[324])^(a[89] & b[325])^(a[88] & b[326])^(a[87] & b[327])^(a[86] & b[328])^(a[85] & b[329])^(a[84] & b[330])^(a[83] & b[331])^(a[82] & b[332])^(a[81] & b[333])^(a[80] & b[334])^(a[79] & b[335])^(a[78] & b[336])^(a[77] & b[337])^(a[76] & b[338])^(a[75] & b[339])^(a[74] & b[340])^(a[73] & b[341])^(a[72] & b[342])^(a[71] & b[343])^(a[70] & b[344])^(a[69] & b[345])^(a[68] & b[346])^(a[67] & b[347])^(a[66] & b[348])^(a[65] & b[349])^(a[64] & b[350])^(a[63] & b[351])^(a[62] & b[352])^(a[61] & b[353])^(a[60] & b[354])^(a[59] & b[355])^(a[58] & b[356])^(a[57] & b[357])^(a[56] & b[358])^(a[55] & b[359])^(a[54] & b[360])^(a[53] & b[361])^(a[52] & b[362])^(a[51] & b[363])^(a[50] & b[364])^(a[49] & b[365])^(a[48] & b[366])^(a[47] & b[367])^(a[46] & b[368])^(a[45] & b[369])^(a[44] & b[370])^(a[43] & b[371])^(a[42] & b[372])^(a[41] & b[373])^(a[40] & b[374])^(a[39] & b[375])^(a[38] & b[376])^(a[37] & b[377])^(a[36] & b[378])^(a[35] & b[379])^(a[34] & b[380])^(a[33] & b[381])^(a[32] & b[382])^(a[31] & b[383])^(a[30] & b[384])^(a[29] & b[385])^(a[28] & b[386])^(a[27] & b[387])^(a[26] & b[388])^(a[25] & b[389])^(a[24] & b[390])^(a[23] & b[391])^(a[22] & b[392])^(a[21] & b[393])^(a[20] & b[394])^(a[19] & b[395])^(a[18] & b[396])^(a[17] & b[397])^(a[16] & b[398])^(a[15] & b[399])^(a[14] & b[400])^(a[13] & b[401])^(a[12] & b[402])^(a[11] & b[403])^(a[10] & b[404])^(a[9] & b[405])^(a[8] & b[406])^(a[7] & b[407])^(a[6] & b[408]);
assign y[415] = (a[408] & b[7])^(a[407] & b[8])^(a[406] & b[9])^(a[405] & b[10])^(a[404] & b[11])^(a[403] & b[12])^(a[402] & b[13])^(a[401] & b[14])^(a[400] & b[15])^(a[399] & b[16])^(a[398] & b[17])^(a[397] & b[18])^(a[396] & b[19])^(a[395] & b[20])^(a[394] & b[21])^(a[393] & b[22])^(a[392] & b[23])^(a[391] & b[24])^(a[390] & b[25])^(a[389] & b[26])^(a[388] & b[27])^(a[387] & b[28])^(a[386] & b[29])^(a[385] & b[30])^(a[384] & b[31])^(a[383] & b[32])^(a[382] & b[33])^(a[381] & b[34])^(a[380] & b[35])^(a[379] & b[36])^(a[378] & b[37])^(a[377] & b[38])^(a[376] & b[39])^(a[375] & b[40])^(a[374] & b[41])^(a[373] & b[42])^(a[372] & b[43])^(a[371] & b[44])^(a[370] & b[45])^(a[369] & b[46])^(a[368] & b[47])^(a[367] & b[48])^(a[366] & b[49])^(a[365] & b[50])^(a[364] & b[51])^(a[363] & b[52])^(a[362] & b[53])^(a[361] & b[54])^(a[360] & b[55])^(a[359] & b[56])^(a[358] & b[57])^(a[357] & b[58])^(a[356] & b[59])^(a[355] & b[60])^(a[354] & b[61])^(a[353] & b[62])^(a[352] & b[63])^(a[351] & b[64])^(a[350] & b[65])^(a[349] & b[66])^(a[348] & b[67])^(a[347] & b[68])^(a[346] & b[69])^(a[345] & b[70])^(a[344] & b[71])^(a[343] & b[72])^(a[342] & b[73])^(a[341] & b[74])^(a[340] & b[75])^(a[339] & b[76])^(a[338] & b[77])^(a[337] & b[78])^(a[336] & b[79])^(a[335] & b[80])^(a[334] & b[81])^(a[333] & b[82])^(a[332] & b[83])^(a[331] & b[84])^(a[330] & b[85])^(a[329] & b[86])^(a[328] & b[87])^(a[327] & b[88])^(a[326] & b[89])^(a[325] & b[90])^(a[324] & b[91])^(a[323] & b[92])^(a[322] & b[93])^(a[321] & b[94])^(a[320] & b[95])^(a[319] & b[96])^(a[318] & b[97])^(a[317] & b[98])^(a[316] & b[99])^(a[315] & b[100])^(a[314] & b[101])^(a[313] & b[102])^(a[312] & b[103])^(a[311] & b[104])^(a[310] & b[105])^(a[309] & b[106])^(a[308] & b[107])^(a[307] & b[108])^(a[306] & b[109])^(a[305] & b[110])^(a[304] & b[111])^(a[303] & b[112])^(a[302] & b[113])^(a[301] & b[114])^(a[300] & b[115])^(a[299] & b[116])^(a[298] & b[117])^(a[297] & b[118])^(a[296] & b[119])^(a[295] & b[120])^(a[294] & b[121])^(a[293] & b[122])^(a[292] & b[123])^(a[291] & b[124])^(a[290] & b[125])^(a[289] & b[126])^(a[288] & b[127])^(a[287] & b[128])^(a[286] & b[129])^(a[285] & b[130])^(a[284] & b[131])^(a[283] & b[132])^(a[282] & b[133])^(a[281] & b[134])^(a[280] & b[135])^(a[279] & b[136])^(a[278] & b[137])^(a[277] & b[138])^(a[276] & b[139])^(a[275] & b[140])^(a[274] & b[141])^(a[273] & b[142])^(a[272] & b[143])^(a[271] & b[144])^(a[270] & b[145])^(a[269] & b[146])^(a[268] & b[147])^(a[267] & b[148])^(a[266] & b[149])^(a[265] & b[150])^(a[264] & b[151])^(a[263] & b[152])^(a[262] & b[153])^(a[261] & b[154])^(a[260] & b[155])^(a[259] & b[156])^(a[258] & b[157])^(a[257] & b[158])^(a[256] & b[159])^(a[255] & b[160])^(a[254] & b[161])^(a[253] & b[162])^(a[252] & b[163])^(a[251] & b[164])^(a[250] & b[165])^(a[249] & b[166])^(a[248] & b[167])^(a[247] & b[168])^(a[246] & b[169])^(a[245] & b[170])^(a[244] & b[171])^(a[243] & b[172])^(a[242] & b[173])^(a[241] & b[174])^(a[240] & b[175])^(a[239] & b[176])^(a[238] & b[177])^(a[237] & b[178])^(a[236] & b[179])^(a[235] & b[180])^(a[234] & b[181])^(a[233] & b[182])^(a[232] & b[183])^(a[231] & b[184])^(a[230] & b[185])^(a[229] & b[186])^(a[228] & b[187])^(a[227] & b[188])^(a[226] & b[189])^(a[225] & b[190])^(a[224] & b[191])^(a[223] & b[192])^(a[222] & b[193])^(a[221] & b[194])^(a[220] & b[195])^(a[219] & b[196])^(a[218] & b[197])^(a[217] & b[198])^(a[216] & b[199])^(a[215] & b[200])^(a[214] & b[201])^(a[213] & b[202])^(a[212] & b[203])^(a[211] & b[204])^(a[210] & b[205])^(a[209] & b[206])^(a[208] & b[207])^(a[207] & b[208])^(a[206] & b[209])^(a[205] & b[210])^(a[204] & b[211])^(a[203] & b[212])^(a[202] & b[213])^(a[201] & b[214])^(a[200] & b[215])^(a[199] & b[216])^(a[198] & b[217])^(a[197] & b[218])^(a[196] & b[219])^(a[195] & b[220])^(a[194] & b[221])^(a[193] & b[222])^(a[192] & b[223])^(a[191] & b[224])^(a[190] & b[225])^(a[189] & b[226])^(a[188] & b[227])^(a[187] & b[228])^(a[186] & b[229])^(a[185] & b[230])^(a[184] & b[231])^(a[183] & b[232])^(a[182] & b[233])^(a[181] & b[234])^(a[180] & b[235])^(a[179] & b[236])^(a[178] & b[237])^(a[177] & b[238])^(a[176] & b[239])^(a[175] & b[240])^(a[174] & b[241])^(a[173] & b[242])^(a[172] & b[243])^(a[171] & b[244])^(a[170] & b[245])^(a[169] & b[246])^(a[168] & b[247])^(a[167] & b[248])^(a[166] & b[249])^(a[165] & b[250])^(a[164] & b[251])^(a[163] & b[252])^(a[162] & b[253])^(a[161] & b[254])^(a[160] & b[255])^(a[159] & b[256])^(a[158] & b[257])^(a[157] & b[258])^(a[156] & b[259])^(a[155] & b[260])^(a[154] & b[261])^(a[153] & b[262])^(a[152] & b[263])^(a[151] & b[264])^(a[150] & b[265])^(a[149] & b[266])^(a[148] & b[267])^(a[147] & b[268])^(a[146] & b[269])^(a[145] & b[270])^(a[144] & b[271])^(a[143] & b[272])^(a[142] & b[273])^(a[141] & b[274])^(a[140] & b[275])^(a[139] & b[276])^(a[138] & b[277])^(a[137] & b[278])^(a[136] & b[279])^(a[135] & b[280])^(a[134] & b[281])^(a[133] & b[282])^(a[132] & b[283])^(a[131] & b[284])^(a[130] & b[285])^(a[129] & b[286])^(a[128] & b[287])^(a[127] & b[288])^(a[126] & b[289])^(a[125] & b[290])^(a[124] & b[291])^(a[123] & b[292])^(a[122] & b[293])^(a[121] & b[294])^(a[120] & b[295])^(a[119] & b[296])^(a[118] & b[297])^(a[117] & b[298])^(a[116] & b[299])^(a[115] & b[300])^(a[114] & b[301])^(a[113] & b[302])^(a[112] & b[303])^(a[111] & b[304])^(a[110] & b[305])^(a[109] & b[306])^(a[108] & b[307])^(a[107] & b[308])^(a[106] & b[309])^(a[105] & b[310])^(a[104] & b[311])^(a[103] & b[312])^(a[102] & b[313])^(a[101] & b[314])^(a[100] & b[315])^(a[99] & b[316])^(a[98] & b[317])^(a[97] & b[318])^(a[96] & b[319])^(a[95] & b[320])^(a[94] & b[321])^(a[93] & b[322])^(a[92] & b[323])^(a[91] & b[324])^(a[90] & b[325])^(a[89] & b[326])^(a[88] & b[327])^(a[87] & b[328])^(a[86] & b[329])^(a[85] & b[330])^(a[84] & b[331])^(a[83] & b[332])^(a[82] & b[333])^(a[81] & b[334])^(a[80] & b[335])^(a[79] & b[336])^(a[78] & b[337])^(a[77] & b[338])^(a[76] & b[339])^(a[75] & b[340])^(a[74] & b[341])^(a[73] & b[342])^(a[72] & b[343])^(a[71] & b[344])^(a[70] & b[345])^(a[69] & b[346])^(a[68] & b[347])^(a[67] & b[348])^(a[66] & b[349])^(a[65] & b[350])^(a[64] & b[351])^(a[63] & b[352])^(a[62] & b[353])^(a[61] & b[354])^(a[60] & b[355])^(a[59] & b[356])^(a[58] & b[357])^(a[57] & b[358])^(a[56] & b[359])^(a[55] & b[360])^(a[54] & b[361])^(a[53] & b[362])^(a[52] & b[363])^(a[51] & b[364])^(a[50] & b[365])^(a[49] & b[366])^(a[48] & b[367])^(a[47] & b[368])^(a[46] & b[369])^(a[45] & b[370])^(a[44] & b[371])^(a[43] & b[372])^(a[42] & b[373])^(a[41] & b[374])^(a[40] & b[375])^(a[39] & b[376])^(a[38] & b[377])^(a[37] & b[378])^(a[36] & b[379])^(a[35] & b[380])^(a[34] & b[381])^(a[33] & b[382])^(a[32] & b[383])^(a[31] & b[384])^(a[30] & b[385])^(a[29] & b[386])^(a[28] & b[387])^(a[27] & b[388])^(a[26] & b[389])^(a[25] & b[390])^(a[24] & b[391])^(a[23] & b[392])^(a[22] & b[393])^(a[21] & b[394])^(a[20] & b[395])^(a[19] & b[396])^(a[18] & b[397])^(a[17] & b[398])^(a[16] & b[399])^(a[15] & b[400])^(a[14] & b[401])^(a[13] & b[402])^(a[12] & b[403])^(a[11] & b[404])^(a[10] & b[405])^(a[9] & b[406])^(a[8] & b[407])^(a[7] & b[408]);
assign y[416] = (a[408] & b[8])^(a[407] & b[9])^(a[406] & b[10])^(a[405] & b[11])^(a[404] & b[12])^(a[403] & b[13])^(a[402] & b[14])^(a[401] & b[15])^(a[400] & b[16])^(a[399] & b[17])^(a[398] & b[18])^(a[397] & b[19])^(a[396] & b[20])^(a[395] & b[21])^(a[394] & b[22])^(a[393] & b[23])^(a[392] & b[24])^(a[391] & b[25])^(a[390] & b[26])^(a[389] & b[27])^(a[388] & b[28])^(a[387] & b[29])^(a[386] & b[30])^(a[385] & b[31])^(a[384] & b[32])^(a[383] & b[33])^(a[382] & b[34])^(a[381] & b[35])^(a[380] & b[36])^(a[379] & b[37])^(a[378] & b[38])^(a[377] & b[39])^(a[376] & b[40])^(a[375] & b[41])^(a[374] & b[42])^(a[373] & b[43])^(a[372] & b[44])^(a[371] & b[45])^(a[370] & b[46])^(a[369] & b[47])^(a[368] & b[48])^(a[367] & b[49])^(a[366] & b[50])^(a[365] & b[51])^(a[364] & b[52])^(a[363] & b[53])^(a[362] & b[54])^(a[361] & b[55])^(a[360] & b[56])^(a[359] & b[57])^(a[358] & b[58])^(a[357] & b[59])^(a[356] & b[60])^(a[355] & b[61])^(a[354] & b[62])^(a[353] & b[63])^(a[352] & b[64])^(a[351] & b[65])^(a[350] & b[66])^(a[349] & b[67])^(a[348] & b[68])^(a[347] & b[69])^(a[346] & b[70])^(a[345] & b[71])^(a[344] & b[72])^(a[343] & b[73])^(a[342] & b[74])^(a[341] & b[75])^(a[340] & b[76])^(a[339] & b[77])^(a[338] & b[78])^(a[337] & b[79])^(a[336] & b[80])^(a[335] & b[81])^(a[334] & b[82])^(a[333] & b[83])^(a[332] & b[84])^(a[331] & b[85])^(a[330] & b[86])^(a[329] & b[87])^(a[328] & b[88])^(a[327] & b[89])^(a[326] & b[90])^(a[325] & b[91])^(a[324] & b[92])^(a[323] & b[93])^(a[322] & b[94])^(a[321] & b[95])^(a[320] & b[96])^(a[319] & b[97])^(a[318] & b[98])^(a[317] & b[99])^(a[316] & b[100])^(a[315] & b[101])^(a[314] & b[102])^(a[313] & b[103])^(a[312] & b[104])^(a[311] & b[105])^(a[310] & b[106])^(a[309] & b[107])^(a[308] & b[108])^(a[307] & b[109])^(a[306] & b[110])^(a[305] & b[111])^(a[304] & b[112])^(a[303] & b[113])^(a[302] & b[114])^(a[301] & b[115])^(a[300] & b[116])^(a[299] & b[117])^(a[298] & b[118])^(a[297] & b[119])^(a[296] & b[120])^(a[295] & b[121])^(a[294] & b[122])^(a[293] & b[123])^(a[292] & b[124])^(a[291] & b[125])^(a[290] & b[126])^(a[289] & b[127])^(a[288] & b[128])^(a[287] & b[129])^(a[286] & b[130])^(a[285] & b[131])^(a[284] & b[132])^(a[283] & b[133])^(a[282] & b[134])^(a[281] & b[135])^(a[280] & b[136])^(a[279] & b[137])^(a[278] & b[138])^(a[277] & b[139])^(a[276] & b[140])^(a[275] & b[141])^(a[274] & b[142])^(a[273] & b[143])^(a[272] & b[144])^(a[271] & b[145])^(a[270] & b[146])^(a[269] & b[147])^(a[268] & b[148])^(a[267] & b[149])^(a[266] & b[150])^(a[265] & b[151])^(a[264] & b[152])^(a[263] & b[153])^(a[262] & b[154])^(a[261] & b[155])^(a[260] & b[156])^(a[259] & b[157])^(a[258] & b[158])^(a[257] & b[159])^(a[256] & b[160])^(a[255] & b[161])^(a[254] & b[162])^(a[253] & b[163])^(a[252] & b[164])^(a[251] & b[165])^(a[250] & b[166])^(a[249] & b[167])^(a[248] & b[168])^(a[247] & b[169])^(a[246] & b[170])^(a[245] & b[171])^(a[244] & b[172])^(a[243] & b[173])^(a[242] & b[174])^(a[241] & b[175])^(a[240] & b[176])^(a[239] & b[177])^(a[238] & b[178])^(a[237] & b[179])^(a[236] & b[180])^(a[235] & b[181])^(a[234] & b[182])^(a[233] & b[183])^(a[232] & b[184])^(a[231] & b[185])^(a[230] & b[186])^(a[229] & b[187])^(a[228] & b[188])^(a[227] & b[189])^(a[226] & b[190])^(a[225] & b[191])^(a[224] & b[192])^(a[223] & b[193])^(a[222] & b[194])^(a[221] & b[195])^(a[220] & b[196])^(a[219] & b[197])^(a[218] & b[198])^(a[217] & b[199])^(a[216] & b[200])^(a[215] & b[201])^(a[214] & b[202])^(a[213] & b[203])^(a[212] & b[204])^(a[211] & b[205])^(a[210] & b[206])^(a[209] & b[207])^(a[208] & b[208])^(a[207] & b[209])^(a[206] & b[210])^(a[205] & b[211])^(a[204] & b[212])^(a[203] & b[213])^(a[202] & b[214])^(a[201] & b[215])^(a[200] & b[216])^(a[199] & b[217])^(a[198] & b[218])^(a[197] & b[219])^(a[196] & b[220])^(a[195] & b[221])^(a[194] & b[222])^(a[193] & b[223])^(a[192] & b[224])^(a[191] & b[225])^(a[190] & b[226])^(a[189] & b[227])^(a[188] & b[228])^(a[187] & b[229])^(a[186] & b[230])^(a[185] & b[231])^(a[184] & b[232])^(a[183] & b[233])^(a[182] & b[234])^(a[181] & b[235])^(a[180] & b[236])^(a[179] & b[237])^(a[178] & b[238])^(a[177] & b[239])^(a[176] & b[240])^(a[175] & b[241])^(a[174] & b[242])^(a[173] & b[243])^(a[172] & b[244])^(a[171] & b[245])^(a[170] & b[246])^(a[169] & b[247])^(a[168] & b[248])^(a[167] & b[249])^(a[166] & b[250])^(a[165] & b[251])^(a[164] & b[252])^(a[163] & b[253])^(a[162] & b[254])^(a[161] & b[255])^(a[160] & b[256])^(a[159] & b[257])^(a[158] & b[258])^(a[157] & b[259])^(a[156] & b[260])^(a[155] & b[261])^(a[154] & b[262])^(a[153] & b[263])^(a[152] & b[264])^(a[151] & b[265])^(a[150] & b[266])^(a[149] & b[267])^(a[148] & b[268])^(a[147] & b[269])^(a[146] & b[270])^(a[145] & b[271])^(a[144] & b[272])^(a[143] & b[273])^(a[142] & b[274])^(a[141] & b[275])^(a[140] & b[276])^(a[139] & b[277])^(a[138] & b[278])^(a[137] & b[279])^(a[136] & b[280])^(a[135] & b[281])^(a[134] & b[282])^(a[133] & b[283])^(a[132] & b[284])^(a[131] & b[285])^(a[130] & b[286])^(a[129] & b[287])^(a[128] & b[288])^(a[127] & b[289])^(a[126] & b[290])^(a[125] & b[291])^(a[124] & b[292])^(a[123] & b[293])^(a[122] & b[294])^(a[121] & b[295])^(a[120] & b[296])^(a[119] & b[297])^(a[118] & b[298])^(a[117] & b[299])^(a[116] & b[300])^(a[115] & b[301])^(a[114] & b[302])^(a[113] & b[303])^(a[112] & b[304])^(a[111] & b[305])^(a[110] & b[306])^(a[109] & b[307])^(a[108] & b[308])^(a[107] & b[309])^(a[106] & b[310])^(a[105] & b[311])^(a[104] & b[312])^(a[103] & b[313])^(a[102] & b[314])^(a[101] & b[315])^(a[100] & b[316])^(a[99] & b[317])^(a[98] & b[318])^(a[97] & b[319])^(a[96] & b[320])^(a[95] & b[321])^(a[94] & b[322])^(a[93] & b[323])^(a[92] & b[324])^(a[91] & b[325])^(a[90] & b[326])^(a[89] & b[327])^(a[88] & b[328])^(a[87] & b[329])^(a[86] & b[330])^(a[85] & b[331])^(a[84] & b[332])^(a[83] & b[333])^(a[82] & b[334])^(a[81] & b[335])^(a[80] & b[336])^(a[79] & b[337])^(a[78] & b[338])^(a[77] & b[339])^(a[76] & b[340])^(a[75] & b[341])^(a[74] & b[342])^(a[73] & b[343])^(a[72] & b[344])^(a[71] & b[345])^(a[70] & b[346])^(a[69] & b[347])^(a[68] & b[348])^(a[67] & b[349])^(a[66] & b[350])^(a[65] & b[351])^(a[64] & b[352])^(a[63] & b[353])^(a[62] & b[354])^(a[61] & b[355])^(a[60] & b[356])^(a[59] & b[357])^(a[58] & b[358])^(a[57] & b[359])^(a[56] & b[360])^(a[55] & b[361])^(a[54] & b[362])^(a[53] & b[363])^(a[52] & b[364])^(a[51] & b[365])^(a[50] & b[366])^(a[49] & b[367])^(a[48] & b[368])^(a[47] & b[369])^(a[46] & b[370])^(a[45] & b[371])^(a[44] & b[372])^(a[43] & b[373])^(a[42] & b[374])^(a[41] & b[375])^(a[40] & b[376])^(a[39] & b[377])^(a[38] & b[378])^(a[37] & b[379])^(a[36] & b[380])^(a[35] & b[381])^(a[34] & b[382])^(a[33] & b[383])^(a[32] & b[384])^(a[31] & b[385])^(a[30] & b[386])^(a[29] & b[387])^(a[28] & b[388])^(a[27] & b[389])^(a[26] & b[390])^(a[25] & b[391])^(a[24] & b[392])^(a[23] & b[393])^(a[22] & b[394])^(a[21] & b[395])^(a[20] & b[396])^(a[19] & b[397])^(a[18] & b[398])^(a[17] & b[399])^(a[16] & b[400])^(a[15] & b[401])^(a[14] & b[402])^(a[13] & b[403])^(a[12] & b[404])^(a[11] & b[405])^(a[10] & b[406])^(a[9] & b[407])^(a[8] & b[408]);
assign y[417] = (a[408] & b[9])^(a[407] & b[10])^(a[406] & b[11])^(a[405] & b[12])^(a[404] & b[13])^(a[403] & b[14])^(a[402] & b[15])^(a[401] & b[16])^(a[400] & b[17])^(a[399] & b[18])^(a[398] & b[19])^(a[397] & b[20])^(a[396] & b[21])^(a[395] & b[22])^(a[394] & b[23])^(a[393] & b[24])^(a[392] & b[25])^(a[391] & b[26])^(a[390] & b[27])^(a[389] & b[28])^(a[388] & b[29])^(a[387] & b[30])^(a[386] & b[31])^(a[385] & b[32])^(a[384] & b[33])^(a[383] & b[34])^(a[382] & b[35])^(a[381] & b[36])^(a[380] & b[37])^(a[379] & b[38])^(a[378] & b[39])^(a[377] & b[40])^(a[376] & b[41])^(a[375] & b[42])^(a[374] & b[43])^(a[373] & b[44])^(a[372] & b[45])^(a[371] & b[46])^(a[370] & b[47])^(a[369] & b[48])^(a[368] & b[49])^(a[367] & b[50])^(a[366] & b[51])^(a[365] & b[52])^(a[364] & b[53])^(a[363] & b[54])^(a[362] & b[55])^(a[361] & b[56])^(a[360] & b[57])^(a[359] & b[58])^(a[358] & b[59])^(a[357] & b[60])^(a[356] & b[61])^(a[355] & b[62])^(a[354] & b[63])^(a[353] & b[64])^(a[352] & b[65])^(a[351] & b[66])^(a[350] & b[67])^(a[349] & b[68])^(a[348] & b[69])^(a[347] & b[70])^(a[346] & b[71])^(a[345] & b[72])^(a[344] & b[73])^(a[343] & b[74])^(a[342] & b[75])^(a[341] & b[76])^(a[340] & b[77])^(a[339] & b[78])^(a[338] & b[79])^(a[337] & b[80])^(a[336] & b[81])^(a[335] & b[82])^(a[334] & b[83])^(a[333] & b[84])^(a[332] & b[85])^(a[331] & b[86])^(a[330] & b[87])^(a[329] & b[88])^(a[328] & b[89])^(a[327] & b[90])^(a[326] & b[91])^(a[325] & b[92])^(a[324] & b[93])^(a[323] & b[94])^(a[322] & b[95])^(a[321] & b[96])^(a[320] & b[97])^(a[319] & b[98])^(a[318] & b[99])^(a[317] & b[100])^(a[316] & b[101])^(a[315] & b[102])^(a[314] & b[103])^(a[313] & b[104])^(a[312] & b[105])^(a[311] & b[106])^(a[310] & b[107])^(a[309] & b[108])^(a[308] & b[109])^(a[307] & b[110])^(a[306] & b[111])^(a[305] & b[112])^(a[304] & b[113])^(a[303] & b[114])^(a[302] & b[115])^(a[301] & b[116])^(a[300] & b[117])^(a[299] & b[118])^(a[298] & b[119])^(a[297] & b[120])^(a[296] & b[121])^(a[295] & b[122])^(a[294] & b[123])^(a[293] & b[124])^(a[292] & b[125])^(a[291] & b[126])^(a[290] & b[127])^(a[289] & b[128])^(a[288] & b[129])^(a[287] & b[130])^(a[286] & b[131])^(a[285] & b[132])^(a[284] & b[133])^(a[283] & b[134])^(a[282] & b[135])^(a[281] & b[136])^(a[280] & b[137])^(a[279] & b[138])^(a[278] & b[139])^(a[277] & b[140])^(a[276] & b[141])^(a[275] & b[142])^(a[274] & b[143])^(a[273] & b[144])^(a[272] & b[145])^(a[271] & b[146])^(a[270] & b[147])^(a[269] & b[148])^(a[268] & b[149])^(a[267] & b[150])^(a[266] & b[151])^(a[265] & b[152])^(a[264] & b[153])^(a[263] & b[154])^(a[262] & b[155])^(a[261] & b[156])^(a[260] & b[157])^(a[259] & b[158])^(a[258] & b[159])^(a[257] & b[160])^(a[256] & b[161])^(a[255] & b[162])^(a[254] & b[163])^(a[253] & b[164])^(a[252] & b[165])^(a[251] & b[166])^(a[250] & b[167])^(a[249] & b[168])^(a[248] & b[169])^(a[247] & b[170])^(a[246] & b[171])^(a[245] & b[172])^(a[244] & b[173])^(a[243] & b[174])^(a[242] & b[175])^(a[241] & b[176])^(a[240] & b[177])^(a[239] & b[178])^(a[238] & b[179])^(a[237] & b[180])^(a[236] & b[181])^(a[235] & b[182])^(a[234] & b[183])^(a[233] & b[184])^(a[232] & b[185])^(a[231] & b[186])^(a[230] & b[187])^(a[229] & b[188])^(a[228] & b[189])^(a[227] & b[190])^(a[226] & b[191])^(a[225] & b[192])^(a[224] & b[193])^(a[223] & b[194])^(a[222] & b[195])^(a[221] & b[196])^(a[220] & b[197])^(a[219] & b[198])^(a[218] & b[199])^(a[217] & b[200])^(a[216] & b[201])^(a[215] & b[202])^(a[214] & b[203])^(a[213] & b[204])^(a[212] & b[205])^(a[211] & b[206])^(a[210] & b[207])^(a[209] & b[208])^(a[208] & b[209])^(a[207] & b[210])^(a[206] & b[211])^(a[205] & b[212])^(a[204] & b[213])^(a[203] & b[214])^(a[202] & b[215])^(a[201] & b[216])^(a[200] & b[217])^(a[199] & b[218])^(a[198] & b[219])^(a[197] & b[220])^(a[196] & b[221])^(a[195] & b[222])^(a[194] & b[223])^(a[193] & b[224])^(a[192] & b[225])^(a[191] & b[226])^(a[190] & b[227])^(a[189] & b[228])^(a[188] & b[229])^(a[187] & b[230])^(a[186] & b[231])^(a[185] & b[232])^(a[184] & b[233])^(a[183] & b[234])^(a[182] & b[235])^(a[181] & b[236])^(a[180] & b[237])^(a[179] & b[238])^(a[178] & b[239])^(a[177] & b[240])^(a[176] & b[241])^(a[175] & b[242])^(a[174] & b[243])^(a[173] & b[244])^(a[172] & b[245])^(a[171] & b[246])^(a[170] & b[247])^(a[169] & b[248])^(a[168] & b[249])^(a[167] & b[250])^(a[166] & b[251])^(a[165] & b[252])^(a[164] & b[253])^(a[163] & b[254])^(a[162] & b[255])^(a[161] & b[256])^(a[160] & b[257])^(a[159] & b[258])^(a[158] & b[259])^(a[157] & b[260])^(a[156] & b[261])^(a[155] & b[262])^(a[154] & b[263])^(a[153] & b[264])^(a[152] & b[265])^(a[151] & b[266])^(a[150] & b[267])^(a[149] & b[268])^(a[148] & b[269])^(a[147] & b[270])^(a[146] & b[271])^(a[145] & b[272])^(a[144] & b[273])^(a[143] & b[274])^(a[142] & b[275])^(a[141] & b[276])^(a[140] & b[277])^(a[139] & b[278])^(a[138] & b[279])^(a[137] & b[280])^(a[136] & b[281])^(a[135] & b[282])^(a[134] & b[283])^(a[133] & b[284])^(a[132] & b[285])^(a[131] & b[286])^(a[130] & b[287])^(a[129] & b[288])^(a[128] & b[289])^(a[127] & b[290])^(a[126] & b[291])^(a[125] & b[292])^(a[124] & b[293])^(a[123] & b[294])^(a[122] & b[295])^(a[121] & b[296])^(a[120] & b[297])^(a[119] & b[298])^(a[118] & b[299])^(a[117] & b[300])^(a[116] & b[301])^(a[115] & b[302])^(a[114] & b[303])^(a[113] & b[304])^(a[112] & b[305])^(a[111] & b[306])^(a[110] & b[307])^(a[109] & b[308])^(a[108] & b[309])^(a[107] & b[310])^(a[106] & b[311])^(a[105] & b[312])^(a[104] & b[313])^(a[103] & b[314])^(a[102] & b[315])^(a[101] & b[316])^(a[100] & b[317])^(a[99] & b[318])^(a[98] & b[319])^(a[97] & b[320])^(a[96] & b[321])^(a[95] & b[322])^(a[94] & b[323])^(a[93] & b[324])^(a[92] & b[325])^(a[91] & b[326])^(a[90] & b[327])^(a[89] & b[328])^(a[88] & b[329])^(a[87] & b[330])^(a[86] & b[331])^(a[85] & b[332])^(a[84] & b[333])^(a[83] & b[334])^(a[82] & b[335])^(a[81] & b[336])^(a[80] & b[337])^(a[79] & b[338])^(a[78] & b[339])^(a[77] & b[340])^(a[76] & b[341])^(a[75] & b[342])^(a[74] & b[343])^(a[73] & b[344])^(a[72] & b[345])^(a[71] & b[346])^(a[70] & b[347])^(a[69] & b[348])^(a[68] & b[349])^(a[67] & b[350])^(a[66] & b[351])^(a[65] & b[352])^(a[64] & b[353])^(a[63] & b[354])^(a[62] & b[355])^(a[61] & b[356])^(a[60] & b[357])^(a[59] & b[358])^(a[58] & b[359])^(a[57] & b[360])^(a[56] & b[361])^(a[55] & b[362])^(a[54] & b[363])^(a[53] & b[364])^(a[52] & b[365])^(a[51] & b[366])^(a[50] & b[367])^(a[49] & b[368])^(a[48] & b[369])^(a[47] & b[370])^(a[46] & b[371])^(a[45] & b[372])^(a[44] & b[373])^(a[43] & b[374])^(a[42] & b[375])^(a[41] & b[376])^(a[40] & b[377])^(a[39] & b[378])^(a[38] & b[379])^(a[37] & b[380])^(a[36] & b[381])^(a[35] & b[382])^(a[34] & b[383])^(a[33] & b[384])^(a[32] & b[385])^(a[31] & b[386])^(a[30] & b[387])^(a[29] & b[388])^(a[28] & b[389])^(a[27] & b[390])^(a[26] & b[391])^(a[25] & b[392])^(a[24] & b[393])^(a[23] & b[394])^(a[22] & b[395])^(a[21] & b[396])^(a[20] & b[397])^(a[19] & b[398])^(a[18] & b[399])^(a[17] & b[400])^(a[16] & b[401])^(a[15] & b[402])^(a[14] & b[403])^(a[13] & b[404])^(a[12] & b[405])^(a[11] & b[406])^(a[10] & b[407])^(a[9] & b[408]);
assign y[418] = (a[408] & b[10])^(a[407] & b[11])^(a[406] & b[12])^(a[405] & b[13])^(a[404] & b[14])^(a[403] & b[15])^(a[402] & b[16])^(a[401] & b[17])^(a[400] & b[18])^(a[399] & b[19])^(a[398] & b[20])^(a[397] & b[21])^(a[396] & b[22])^(a[395] & b[23])^(a[394] & b[24])^(a[393] & b[25])^(a[392] & b[26])^(a[391] & b[27])^(a[390] & b[28])^(a[389] & b[29])^(a[388] & b[30])^(a[387] & b[31])^(a[386] & b[32])^(a[385] & b[33])^(a[384] & b[34])^(a[383] & b[35])^(a[382] & b[36])^(a[381] & b[37])^(a[380] & b[38])^(a[379] & b[39])^(a[378] & b[40])^(a[377] & b[41])^(a[376] & b[42])^(a[375] & b[43])^(a[374] & b[44])^(a[373] & b[45])^(a[372] & b[46])^(a[371] & b[47])^(a[370] & b[48])^(a[369] & b[49])^(a[368] & b[50])^(a[367] & b[51])^(a[366] & b[52])^(a[365] & b[53])^(a[364] & b[54])^(a[363] & b[55])^(a[362] & b[56])^(a[361] & b[57])^(a[360] & b[58])^(a[359] & b[59])^(a[358] & b[60])^(a[357] & b[61])^(a[356] & b[62])^(a[355] & b[63])^(a[354] & b[64])^(a[353] & b[65])^(a[352] & b[66])^(a[351] & b[67])^(a[350] & b[68])^(a[349] & b[69])^(a[348] & b[70])^(a[347] & b[71])^(a[346] & b[72])^(a[345] & b[73])^(a[344] & b[74])^(a[343] & b[75])^(a[342] & b[76])^(a[341] & b[77])^(a[340] & b[78])^(a[339] & b[79])^(a[338] & b[80])^(a[337] & b[81])^(a[336] & b[82])^(a[335] & b[83])^(a[334] & b[84])^(a[333] & b[85])^(a[332] & b[86])^(a[331] & b[87])^(a[330] & b[88])^(a[329] & b[89])^(a[328] & b[90])^(a[327] & b[91])^(a[326] & b[92])^(a[325] & b[93])^(a[324] & b[94])^(a[323] & b[95])^(a[322] & b[96])^(a[321] & b[97])^(a[320] & b[98])^(a[319] & b[99])^(a[318] & b[100])^(a[317] & b[101])^(a[316] & b[102])^(a[315] & b[103])^(a[314] & b[104])^(a[313] & b[105])^(a[312] & b[106])^(a[311] & b[107])^(a[310] & b[108])^(a[309] & b[109])^(a[308] & b[110])^(a[307] & b[111])^(a[306] & b[112])^(a[305] & b[113])^(a[304] & b[114])^(a[303] & b[115])^(a[302] & b[116])^(a[301] & b[117])^(a[300] & b[118])^(a[299] & b[119])^(a[298] & b[120])^(a[297] & b[121])^(a[296] & b[122])^(a[295] & b[123])^(a[294] & b[124])^(a[293] & b[125])^(a[292] & b[126])^(a[291] & b[127])^(a[290] & b[128])^(a[289] & b[129])^(a[288] & b[130])^(a[287] & b[131])^(a[286] & b[132])^(a[285] & b[133])^(a[284] & b[134])^(a[283] & b[135])^(a[282] & b[136])^(a[281] & b[137])^(a[280] & b[138])^(a[279] & b[139])^(a[278] & b[140])^(a[277] & b[141])^(a[276] & b[142])^(a[275] & b[143])^(a[274] & b[144])^(a[273] & b[145])^(a[272] & b[146])^(a[271] & b[147])^(a[270] & b[148])^(a[269] & b[149])^(a[268] & b[150])^(a[267] & b[151])^(a[266] & b[152])^(a[265] & b[153])^(a[264] & b[154])^(a[263] & b[155])^(a[262] & b[156])^(a[261] & b[157])^(a[260] & b[158])^(a[259] & b[159])^(a[258] & b[160])^(a[257] & b[161])^(a[256] & b[162])^(a[255] & b[163])^(a[254] & b[164])^(a[253] & b[165])^(a[252] & b[166])^(a[251] & b[167])^(a[250] & b[168])^(a[249] & b[169])^(a[248] & b[170])^(a[247] & b[171])^(a[246] & b[172])^(a[245] & b[173])^(a[244] & b[174])^(a[243] & b[175])^(a[242] & b[176])^(a[241] & b[177])^(a[240] & b[178])^(a[239] & b[179])^(a[238] & b[180])^(a[237] & b[181])^(a[236] & b[182])^(a[235] & b[183])^(a[234] & b[184])^(a[233] & b[185])^(a[232] & b[186])^(a[231] & b[187])^(a[230] & b[188])^(a[229] & b[189])^(a[228] & b[190])^(a[227] & b[191])^(a[226] & b[192])^(a[225] & b[193])^(a[224] & b[194])^(a[223] & b[195])^(a[222] & b[196])^(a[221] & b[197])^(a[220] & b[198])^(a[219] & b[199])^(a[218] & b[200])^(a[217] & b[201])^(a[216] & b[202])^(a[215] & b[203])^(a[214] & b[204])^(a[213] & b[205])^(a[212] & b[206])^(a[211] & b[207])^(a[210] & b[208])^(a[209] & b[209])^(a[208] & b[210])^(a[207] & b[211])^(a[206] & b[212])^(a[205] & b[213])^(a[204] & b[214])^(a[203] & b[215])^(a[202] & b[216])^(a[201] & b[217])^(a[200] & b[218])^(a[199] & b[219])^(a[198] & b[220])^(a[197] & b[221])^(a[196] & b[222])^(a[195] & b[223])^(a[194] & b[224])^(a[193] & b[225])^(a[192] & b[226])^(a[191] & b[227])^(a[190] & b[228])^(a[189] & b[229])^(a[188] & b[230])^(a[187] & b[231])^(a[186] & b[232])^(a[185] & b[233])^(a[184] & b[234])^(a[183] & b[235])^(a[182] & b[236])^(a[181] & b[237])^(a[180] & b[238])^(a[179] & b[239])^(a[178] & b[240])^(a[177] & b[241])^(a[176] & b[242])^(a[175] & b[243])^(a[174] & b[244])^(a[173] & b[245])^(a[172] & b[246])^(a[171] & b[247])^(a[170] & b[248])^(a[169] & b[249])^(a[168] & b[250])^(a[167] & b[251])^(a[166] & b[252])^(a[165] & b[253])^(a[164] & b[254])^(a[163] & b[255])^(a[162] & b[256])^(a[161] & b[257])^(a[160] & b[258])^(a[159] & b[259])^(a[158] & b[260])^(a[157] & b[261])^(a[156] & b[262])^(a[155] & b[263])^(a[154] & b[264])^(a[153] & b[265])^(a[152] & b[266])^(a[151] & b[267])^(a[150] & b[268])^(a[149] & b[269])^(a[148] & b[270])^(a[147] & b[271])^(a[146] & b[272])^(a[145] & b[273])^(a[144] & b[274])^(a[143] & b[275])^(a[142] & b[276])^(a[141] & b[277])^(a[140] & b[278])^(a[139] & b[279])^(a[138] & b[280])^(a[137] & b[281])^(a[136] & b[282])^(a[135] & b[283])^(a[134] & b[284])^(a[133] & b[285])^(a[132] & b[286])^(a[131] & b[287])^(a[130] & b[288])^(a[129] & b[289])^(a[128] & b[290])^(a[127] & b[291])^(a[126] & b[292])^(a[125] & b[293])^(a[124] & b[294])^(a[123] & b[295])^(a[122] & b[296])^(a[121] & b[297])^(a[120] & b[298])^(a[119] & b[299])^(a[118] & b[300])^(a[117] & b[301])^(a[116] & b[302])^(a[115] & b[303])^(a[114] & b[304])^(a[113] & b[305])^(a[112] & b[306])^(a[111] & b[307])^(a[110] & b[308])^(a[109] & b[309])^(a[108] & b[310])^(a[107] & b[311])^(a[106] & b[312])^(a[105] & b[313])^(a[104] & b[314])^(a[103] & b[315])^(a[102] & b[316])^(a[101] & b[317])^(a[100] & b[318])^(a[99] & b[319])^(a[98] & b[320])^(a[97] & b[321])^(a[96] & b[322])^(a[95] & b[323])^(a[94] & b[324])^(a[93] & b[325])^(a[92] & b[326])^(a[91] & b[327])^(a[90] & b[328])^(a[89] & b[329])^(a[88] & b[330])^(a[87] & b[331])^(a[86] & b[332])^(a[85] & b[333])^(a[84] & b[334])^(a[83] & b[335])^(a[82] & b[336])^(a[81] & b[337])^(a[80] & b[338])^(a[79] & b[339])^(a[78] & b[340])^(a[77] & b[341])^(a[76] & b[342])^(a[75] & b[343])^(a[74] & b[344])^(a[73] & b[345])^(a[72] & b[346])^(a[71] & b[347])^(a[70] & b[348])^(a[69] & b[349])^(a[68] & b[350])^(a[67] & b[351])^(a[66] & b[352])^(a[65] & b[353])^(a[64] & b[354])^(a[63] & b[355])^(a[62] & b[356])^(a[61] & b[357])^(a[60] & b[358])^(a[59] & b[359])^(a[58] & b[360])^(a[57] & b[361])^(a[56] & b[362])^(a[55] & b[363])^(a[54] & b[364])^(a[53] & b[365])^(a[52] & b[366])^(a[51] & b[367])^(a[50] & b[368])^(a[49] & b[369])^(a[48] & b[370])^(a[47] & b[371])^(a[46] & b[372])^(a[45] & b[373])^(a[44] & b[374])^(a[43] & b[375])^(a[42] & b[376])^(a[41] & b[377])^(a[40] & b[378])^(a[39] & b[379])^(a[38] & b[380])^(a[37] & b[381])^(a[36] & b[382])^(a[35] & b[383])^(a[34] & b[384])^(a[33] & b[385])^(a[32] & b[386])^(a[31] & b[387])^(a[30] & b[388])^(a[29] & b[389])^(a[28] & b[390])^(a[27] & b[391])^(a[26] & b[392])^(a[25] & b[393])^(a[24] & b[394])^(a[23] & b[395])^(a[22] & b[396])^(a[21] & b[397])^(a[20] & b[398])^(a[19] & b[399])^(a[18] & b[400])^(a[17] & b[401])^(a[16] & b[402])^(a[15] & b[403])^(a[14] & b[404])^(a[13] & b[405])^(a[12] & b[406])^(a[11] & b[407])^(a[10] & b[408]);
assign y[419] = (a[408] & b[11])^(a[407] & b[12])^(a[406] & b[13])^(a[405] & b[14])^(a[404] & b[15])^(a[403] & b[16])^(a[402] & b[17])^(a[401] & b[18])^(a[400] & b[19])^(a[399] & b[20])^(a[398] & b[21])^(a[397] & b[22])^(a[396] & b[23])^(a[395] & b[24])^(a[394] & b[25])^(a[393] & b[26])^(a[392] & b[27])^(a[391] & b[28])^(a[390] & b[29])^(a[389] & b[30])^(a[388] & b[31])^(a[387] & b[32])^(a[386] & b[33])^(a[385] & b[34])^(a[384] & b[35])^(a[383] & b[36])^(a[382] & b[37])^(a[381] & b[38])^(a[380] & b[39])^(a[379] & b[40])^(a[378] & b[41])^(a[377] & b[42])^(a[376] & b[43])^(a[375] & b[44])^(a[374] & b[45])^(a[373] & b[46])^(a[372] & b[47])^(a[371] & b[48])^(a[370] & b[49])^(a[369] & b[50])^(a[368] & b[51])^(a[367] & b[52])^(a[366] & b[53])^(a[365] & b[54])^(a[364] & b[55])^(a[363] & b[56])^(a[362] & b[57])^(a[361] & b[58])^(a[360] & b[59])^(a[359] & b[60])^(a[358] & b[61])^(a[357] & b[62])^(a[356] & b[63])^(a[355] & b[64])^(a[354] & b[65])^(a[353] & b[66])^(a[352] & b[67])^(a[351] & b[68])^(a[350] & b[69])^(a[349] & b[70])^(a[348] & b[71])^(a[347] & b[72])^(a[346] & b[73])^(a[345] & b[74])^(a[344] & b[75])^(a[343] & b[76])^(a[342] & b[77])^(a[341] & b[78])^(a[340] & b[79])^(a[339] & b[80])^(a[338] & b[81])^(a[337] & b[82])^(a[336] & b[83])^(a[335] & b[84])^(a[334] & b[85])^(a[333] & b[86])^(a[332] & b[87])^(a[331] & b[88])^(a[330] & b[89])^(a[329] & b[90])^(a[328] & b[91])^(a[327] & b[92])^(a[326] & b[93])^(a[325] & b[94])^(a[324] & b[95])^(a[323] & b[96])^(a[322] & b[97])^(a[321] & b[98])^(a[320] & b[99])^(a[319] & b[100])^(a[318] & b[101])^(a[317] & b[102])^(a[316] & b[103])^(a[315] & b[104])^(a[314] & b[105])^(a[313] & b[106])^(a[312] & b[107])^(a[311] & b[108])^(a[310] & b[109])^(a[309] & b[110])^(a[308] & b[111])^(a[307] & b[112])^(a[306] & b[113])^(a[305] & b[114])^(a[304] & b[115])^(a[303] & b[116])^(a[302] & b[117])^(a[301] & b[118])^(a[300] & b[119])^(a[299] & b[120])^(a[298] & b[121])^(a[297] & b[122])^(a[296] & b[123])^(a[295] & b[124])^(a[294] & b[125])^(a[293] & b[126])^(a[292] & b[127])^(a[291] & b[128])^(a[290] & b[129])^(a[289] & b[130])^(a[288] & b[131])^(a[287] & b[132])^(a[286] & b[133])^(a[285] & b[134])^(a[284] & b[135])^(a[283] & b[136])^(a[282] & b[137])^(a[281] & b[138])^(a[280] & b[139])^(a[279] & b[140])^(a[278] & b[141])^(a[277] & b[142])^(a[276] & b[143])^(a[275] & b[144])^(a[274] & b[145])^(a[273] & b[146])^(a[272] & b[147])^(a[271] & b[148])^(a[270] & b[149])^(a[269] & b[150])^(a[268] & b[151])^(a[267] & b[152])^(a[266] & b[153])^(a[265] & b[154])^(a[264] & b[155])^(a[263] & b[156])^(a[262] & b[157])^(a[261] & b[158])^(a[260] & b[159])^(a[259] & b[160])^(a[258] & b[161])^(a[257] & b[162])^(a[256] & b[163])^(a[255] & b[164])^(a[254] & b[165])^(a[253] & b[166])^(a[252] & b[167])^(a[251] & b[168])^(a[250] & b[169])^(a[249] & b[170])^(a[248] & b[171])^(a[247] & b[172])^(a[246] & b[173])^(a[245] & b[174])^(a[244] & b[175])^(a[243] & b[176])^(a[242] & b[177])^(a[241] & b[178])^(a[240] & b[179])^(a[239] & b[180])^(a[238] & b[181])^(a[237] & b[182])^(a[236] & b[183])^(a[235] & b[184])^(a[234] & b[185])^(a[233] & b[186])^(a[232] & b[187])^(a[231] & b[188])^(a[230] & b[189])^(a[229] & b[190])^(a[228] & b[191])^(a[227] & b[192])^(a[226] & b[193])^(a[225] & b[194])^(a[224] & b[195])^(a[223] & b[196])^(a[222] & b[197])^(a[221] & b[198])^(a[220] & b[199])^(a[219] & b[200])^(a[218] & b[201])^(a[217] & b[202])^(a[216] & b[203])^(a[215] & b[204])^(a[214] & b[205])^(a[213] & b[206])^(a[212] & b[207])^(a[211] & b[208])^(a[210] & b[209])^(a[209] & b[210])^(a[208] & b[211])^(a[207] & b[212])^(a[206] & b[213])^(a[205] & b[214])^(a[204] & b[215])^(a[203] & b[216])^(a[202] & b[217])^(a[201] & b[218])^(a[200] & b[219])^(a[199] & b[220])^(a[198] & b[221])^(a[197] & b[222])^(a[196] & b[223])^(a[195] & b[224])^(a[194] & b[225])^(a[193] & b[226])^(a[192] & b[227])^(a[191] & b[228])^(a[190] & b[229])^(a[189] & b[230])^(a[188] & b[231])^(a[187] & b[232])^(a[186] & b[233])^(a[185] & b[234])^(a[184] & b[235])^(a[183] & b[236])^(a[182] & b[237])^(a[181] & b[238])^(a[180] & b[239])^(a[179] & b[240])^(a[178] & b[241])^(a[177] & b[242])^(a[176] & b[243])^(a[175] & b[244])^(a[174] & b[245])^(a[173] & b[246])^(a[172] & b[247])^(a[171] & b[248])^(a[170] & b[249])^(a[169] & b[250])^(a[168] & b[251])^(a[167] & b[252])^(a[166] & b[253])^(a[165] & b[254])^(a[164] & b[255])^(a[163] & b[256])^(a[162] & b[257])^(a[161] & b[258])^(a[160] & b[259])^(a[159] & b[260])^(a[158] & b[261])^(a[157] & b[262])^(a[156] & b[263])^(a[155] & b[264])^(a[154] & b[265])^(a[153] & b[266])^(a[152] & b[267])^(a[151] & b[268])^(a[150] & b[269])^(a[149] & b[270])^(a[148] & b[271])^(a[147] & b[272])^(a[146] & b[273])^(a[145] & b[274])^(a[144] & b[275])^(a[143] & b[276])^(a[142] & b[277])^(a[141] & b[278])^(a[140] & b[279])^(a[139] & b[280])^(a[138] & b[281])^(a[137] & b[282])^(a[136] & b[283])^(a[135] & b[284])^(a[134] & b[285])^(a[133] & b[286])^(a[132] & b[287])^(a[131] & b[288])^(a[130] & b[289])^(a[129] & b[290])^(a[128] & b[291])^(a[127] & b[292])^(a[126] & b[293])^(a[125] & b[294])^(a[124] & b[295])^(a[123] & b[296])^(a[122] & b[297])^(a[121] & b[298])^(a[120] & b[299])^(a[119] & b[300])^(a[118] & b[301])^(a[117] & b[302])^(a[116] & b[303])^(a[115] & b[304])^(a[114] & b[305])^(a[113] & b[306])^(a[112] & b[307])^(a[111] & b[308])^(a[110] & b[309])^(a[109] & b[310])^(a[108] & b[311])^(a[107] & b[312])^(a[106] & b[313])^(a[105] & b[314])^(a[104] & b[315])^(a[103] & b[316])^(a[102] & b[317])^(a[101] & b[318])^(a[100] & b[319])^(a[99] & b[320])^(a[98] & b[321])^(a[97] & b[322])^(a[96] & b[323])^(a[95] & b[324])^(a[94] & b[325])^(a[93] & b[326])^(a[92] & b[327])^(a[91] & b[328])^(a[90] & b[329])^(a[89] & b[330])^(a[88] & b[331])^(a[87] & b[332])^(a[86] & b[333])^(a[85] & b[334])^(a[84] & b[335])^(a[83] & b[336])^(a[82] & b[337])^(a[81] & b[338])^(a[80] & b[339])^(a[79] & b[340])^(a[78] & b[341])^(a[77] & b[342])^(a[76] & b[343])^(a[75] & b[344])^(a[74] & b[345])^(a[73] & b[346])^(a[72] & b[347])^(a[71] & b[348])^(a[70] & b[349])^(a[69] & b[350])^(a[68] & b[351])^(a[67] & b[352])^(a[66] & b[353])^(a[65] & b[354])^(a[64] & b[355])^(a[63] & b[356])^(a[62] & b[357])^(a[61] & b[358])^(a[60] & b[359])^(a[59] & b[360])^(a[58] & b[361])^(a[57] & b[362])^(a[56] & b[363])^(a[55] & b[364])^(a[54] & b[365])^(a[53] & b[366])^(a[52] & b[367])^(a[51] & b[368])^(a[50] & b[369])^(a[49] & b[370])^(a[48] & b[371])^(a[47] & b[372])^(a[46] & b[373])^(a[45] & b[374])^(a[44] & b[375])^(a[43] & b[376])^(a[42] & b[377])^(a[41] & b[378])^(a[40] & b[379])^(a[39] & b[380])^(a[38] & b[381])^(a[37] & b[382])^(a[36] & b[383])^(a[35] & b[384])^(a[34] & b[385])^(a[33] & b[386])^(a[32] & b[387])^(a[31] & b[388])^(a[30] & b[389])^(a[29] & b[390])^(a[28] & b[391])^(a[27] & b[392])^(a[26] & b[393])^(a[25] & b[394])^(a[24] & b[395])^(a[23] & b[396])^(a[22] & b[397])^(a[21] & b[398])^(a[20] & b[399])^(a[19] & b[400])^(a[18] & b[401])^(a[17] & b[402])^(a[16] & b[403])^(a[15] & b[404])^(a[14] & b[405])^(a[13] & b[406])^(a[12] & b[407])^(a[11] & b[408]);
assign y[420] = (a[408] & b[12])^(a[407] & b[13])^(a[406] & b[14])^(a[405] & b[15])^(a[404] & b[16])^(a[403] & b[17])^(a[402] & b[18])^(a[401] & b[19])^(a[400] & b[20])^(a[399] & b[21])^(a[398] & b[22])^(a[397] & b[23])^(a[396] & b[24])^(a[395] & b[25])^(a[394] & b[26])^(a[393] & b[27])^(a[392] & b[28])^(a[391] & b[29])^(a[390] & b[30])^(a[389] & b[31])^(a[388] & b[32])^(a[387] & b[33])^(a[386] & b[34])^(a[385] & b[35])^(a[384] & b[36])^(a[383] & b[37])^(a[382] & b[38])^(a[381] & b[39])^(a[380] & b[40])^(a[379] & b[41])^(a[378] & b[42])^(a[377] & b[43])^(a[376] & b[44])^(a[375] & b[45])^(a[374] & b[46])^(a[373] & b[47])^(a[372] & b[48])^(a[371] & b[49])^(a[370] & b[50])^(a[369] & b[51])^(a[368] & b[52])^(a[367] & b[53])^(a[366] & b[54])^(a[365] & b[55])^(a[364] & b[56])^(a[363] & b[57])^(a[362] & b[58])^(a[361] & b[59])^(a[360] & b[60])^(a[359] & b[61])^(a[358] & b[62])^(a[357] & b[63])^(a[356] & b[64])^(a[355] & b[65])^(a[354] & b[66])^(a[353] & b[67])^(a[352] & b[68])^(a[351] & b[69])^(a[350] & b[70])^(a[349] & b[71])^(a[348] & b[72])^(a[347] & b[73])^(a[346] & b[74])^(a[345] & b[75])^(a[344] & b[76])^(a[343] & b[77])^(a[342] & b[78])^(a[341] & b[79])^(a[340] & b[80])^(a[339] & b[81])^(a[338] & b[82])^(a[337] & b[83])^(a[336] & b[84])^(a[335] & b[85])^(a[334] & b[86])^(a[333] & b[87])^(a[332] & b[88])^(a[331] & b[89])^(a[330] & b[90])^(a[329] & b[91])^(a[328] & b[92])^(a[327] & b[93])^(a[326] & b[94])^(a[325] & b[95])^(a[324] & b[96])^(a[323] & b[97])^(a[322] & b[98])^(a[321] & b[99])^(a[320] & b[100])^(a[319] & b[101])^(a[318] & b[102])^(a[317] & b[103])^(a[316] & b[104])^(a[315] & b[105])^(a[314] & b[106])^(a[313] & b[107])^(a[312] & b[108])^(a[311] & b[109])^(a[310] & b[110])^(a[309] & b[111])^(a[308] & b[112])^(a[307] & b[113])^(a[306] & b[114])^(a[305] & b[115])^(a[304] & b[116])^(a[303] & b[117])^(a[302] & b[118])^(a[301] & b[119])^(a[300] & b[120])^(a[299] & b[121])^(a[298] & b[122])^(a[297] & b[123])^(a[296] & b[124])^(a[295] & b[125])^(a[294] & b[126])^(a[293] & b[127])^(a[292] & b[128])^(a[291] & b[129])^(a[290] & b[130])^(a[289] & b[131])^(a[288] & b[132])^(a[287] & b[133])^(a[286] & b[134])^(a[285] & b[135])^(a[284] & b[136])^(a[283] & b[137])^(a[282] & b[138])^(a[281] & b[139])^(a[280] & b[140])^(a[279] & b[141])^(a[278] & b[142])^(a[277] & b[143])^(a[276] & b[144])^(a[275] & b[145])^(a[274] & b[146])^(a[273] & b[147])^(a[272] & b[148])^(a[271] & b[149])^(a[270] & b[150])^(a[269] & b[151])^(a[268] & b[152])^(a[267] & b[153])^(a[266] & b[154])^(a[265] & b[155])^(a[264] & b[156])^(a[263] & b[157])^(a[262] & b[158])^(a[261] & b[159])^(a[260] & b[160])^(a[259] & b[161])^(a[258] & b[162])^(a[257] & b[163])^(a[256] & b[164])^(a[255] & b[165])^(a[254] & b[166])^(a[253] & b[167])^(a[252] & b[168])^(a[251] & b[169])^(a[250] & b[170])^(a[249] & b[171])^(a[248] & b[172])^(a[247] & b[173])^(a[246] & b[174])^(a[245] & b[175])^(a[244] & b[176])^(a[243] & b[177])^(a[242] & b[178])^(a[241] & b[179])^(a[240] & b[180])^(a[239] & b[181])^(a[238] & b[182])^(a[237] & b[183])^(a[236] & b[184])^(a[235] & b[185])^(a[234] & b[186])^(a[233] & b[187])^(a[232] & b[188])^(a[231] & b[189])^(a[230] & b[190])^(a[229] & b[191])^(a[228] & b[192])^(a[227] & b[193])^(a[226] & b[194])^(a[225] & b[195])^(a[224] & b[196])^(a[223] & b[197])^(a[222] & b[198])^(a[221] & b[199])^(a[220] & b[200])^(a[219] & b[201])^(a[218] & b[202])^(a[217] & b[203])^(a[216] & b[204])^(a[215] & b[205])^(a[214] & b[206])^(a[213] & b[207])^(a[212] & b[208])^(a[211] & b[209])^(a[210] & b[210])^(a[209] & b[211])^(a[208] & b[212])^(a[207] & b[213])^(a[206] & b[214])^(a[205] & b[215])^(a[204] & b[216])^(a[203] & b[217])^(a[202] & b[218])^(a[201] & b[219])^(a[200] & b[220])^(a[199] & b[221])^(a[198] & b[222])^(a[197] & b[223])^(a[196] & b[224])^(a[195] & b[225])^(a[194] & b[226])^(a[193] & b[227])^(a[192] & b[228])^(a[191] & b[229])^(a[190] & b[230])^(a[189] & b[231])^(a[188] & b[232])^(a[187] & b[233])^(a[186] & b[234])^(a[185] & b[235])^(a[184] & b[236])^(a[183] & b[237])^(a[182] & b[238])^(a[181] & b[239])^(a[180] & b[240])^(a[179] & b[241])^(a[178] & b[242])^(a[177] & b[243])^(a[176] & b[244])^(a[175] & b[245])^(a[174] & b[246])^(a[173] & b[247])^(a[172] & b[248])^(a[171] & b[249])^(a[170] & b[250])^(a[169] & b[251])^(a[168] & b[252])^(a[167] & b[253])^(a[166] & b[254])^(a[165] & b[255])^(a[164] & b[256])^(a[163] & b[257])^(a[162] & b[258])^(a[161] & b[259])^(a[160] & b[260])^(a[159] & b[261])^(a[158] & b[262])^(a[157] & b[263])^(a[156] & b[264])^(a[155] & b[265])^(a[154] & b[266])^(a[153] & b[267])^(a[152] & b[268])^(a[151] & b[269])^(a[150] & b[270])^(a[149] & b[271])^(a[148] & b[272])^(a[147] & b[273])^(a[146] & b[274])^(a[145] & b[275])^(a[144] & b[276])^(a[143] & b[277])^(a[142] & b[278])^(a[141] & b[279])^(a[140] & b[280])^(a[139] & b[281])^(a[138] & b[282])^(a[137] & b[283])^(a[136] & b[284])^(a[135] & b[285])^(a[134] & b[286])^(a[133] & b[287])^(a[132] & b[288])^(a[131] & b[289])^(a[130] & b[290])^(a[129] & b[291])^(a[128] & b[292])^(a[127] & b[293])^(a[126] & b[294])^(a[125] & b[295])^(a[124] & b[296])^(a[123] & b[297])^(a[122] & b[298])^(a[121] & b[299])^(a[120] & b[300])^(a[119] & b[301])^(a[118] & b[302])^(a[117] & b[303])^(a[116] & b[304])^(a[115] & b[305])^(a[114] & b[306])^(a[113] & b[307])^(a[112] & b[308])^(a[111] & b[309])^(a[110] & b[310])^(a[109] & b[311])^(a[108] & b[312])^(a[107] & b[313])^(a[106] & b[314])^(a[105] & b[315])^(a[104] & b[316])^(a[103] & b[317])^(a[102] & b[318])^(a[101] & b[319])^(a[100] & b[320])^(a[99] & b[321])^(a[98] & b[322])^(a[97] & b[323])^(a[96] & b[324])^(a[95] & b[325])^(a[94] & b[326])^(a[93] & b[327])^(a[92] & b[328])^(a[91] & b[329])^(a[90] & b[330])^(a[89] & b[331])^(a[88] & b[332])^(a[87] & b[333])^(a[86] & b[334])^(a[85] & b[335])^(a[84] & b[336])^(a[83] & b[337])^(a[82] & b[338])^(a[81] & b[339])^(a[80] & b[340])^(a[79] & b[341])^(a[78] & b[342])^(a[77] & b[343])^(a[76] & b[344])^(a[75] & b[345])^(a[74] & b[346])^(a[73] & b[347])^(a[72] & b[348])^(a[71] & b[349])^(a[70] & b[350])^(a[69] & b[351])^(a[68] & b[352])^(a[67] & b[353])^(a[66] & b[354])^(a[65] & b[355])^(a[64] & b[356])^(a[63] & b[357])^(a[62] & b[358])^(a[61] & b[359])^(a[60] & b[360])^(a[59] & b[361])^(a[58] & b[362])^(a[57] & b[363])^(a[56] & b[364])^(a[55] & b[365])^(a[54] & b[366])^(a[53] & b[367])^(a[52] & b[368])^(a[51] & b[369])^(a[50] & b[370])^(a[49] & b[371])^(a[48] & b[372])^(a[47] & b[373])^(a[46] & b[374])^(a[45] & b[375])^(a[44] & b[376])^(a[43] & b[377])^(a[42] & b[378])^(a[41] & b[379])^(a[40] & b[380])^(a[39] & b[381])^(a[38] & b[382])^(a[37] & b[383])^(a[36] & b[384])^(a[35] & b[385])^(a[34] & b[386])^(a[33] & b[387])^(a[32] & b[388])^(a[31] & b[389])^(a[30] & b[390])^(a[29] & b[391])^(a[28] & b[392])^(a[27] & b[393])^(a[26] & b[394])^(a[25] & b[395])^(a[24] & b[396])^(a[23] & b[397])^(a[22] & b[398])^(a[21] & b[399])^(a[20] & b[400])^(a[19] & b[401])^(a[18] & b[402])^(a[17] & b[403])^(a[16] & b[404])^(a[15] & b[405])^(a[14] & b[406])^(a[13] & b[407])^(a[12] & b[408]);
assign y[421] = (a[408] & b[13])^(a[407] & b[14])^(a[406] & b[15])^(a[405] & b[16])^(a[404] & b[17])^(a[403] & b[18])^(a[402] & b[19])^(a[401] & b[20])^(a[400] & b[21])^(a[399] & b[22])^(a[398] & b[23])^(a[397] & b[24])^(a[396] & b[25])^(a[395] & b[26])^(a[394] & b[27])^(a[393] & b[28])^(a[392] & b[29])^(a[391] & b[30])^(a[390] & b[31])^(a[389] & b[32])^(a[388] & b[33])^(a[387] & b[34])^(a[386] & b[35])^(a[385] & b[36])^(a[384] & b[37])^(a[383] & b[38])^(a[382] & b[39])^(a[381] & b[40])^(a[380] & b[41])^(a[379] & b[42])^(a[378] & b[43])^(a[377] & b[44])^(a[376] & b[45])^(a[375] & b[46])^(a[374] & b[47])^(a[373] & b[48])^(a[372] & b[49])^(a[371] & b[50])^(a[370] & b[51])^(a[369] & b[52])^(a[368] & b[53])^(a[367] & b[54])^(a[366] & b[55])^(a[365] & b[56])^(a[364] & b[57])^(a[363] & b[58])^(a[362] & b[59])^(a[361] & b[60])^(a[360] & b[61])^(a[359] & b[62])^(a[358] & b[63])^(a[357] & b[64])^(a[356] & b[65])^(a[355] & b[66])^(a[354] & b[67])^(a[353] & b[68])^(a[352] & b[69])^(a[351] & b[70])^(a[350] & b[71])^(a[349] & b[72])^(a[348] & b[73])^(a[347] & b[74])^(a[346] & b[75])^(a[345] & b[76])^(a[344] & b[77])^(a[343] & b[78])^(a[342] & b[79])^(a[341] & b[80])^(a[340] & b[81])^(a[339] & b[82])^(a[338] & b[83])^(a[337] & b[84])^(a[336] & b[85])^(a[335] & b[86])^(a[334] & b[87])^(a[333] & b[88])^(a[332] & b[89])^(a[331] & b[90])^(a[330] & b[91])^(a[329] & b[92])^(a[328] & b[93])^(a[327] & b[94])^(a[326] & b[95])^(a[325] & b[96])^(a[324] & b[97])^(a[323] & b[98])^(a[322] & b[99])^(a[321] & b[100])^(a[320] & b[101])^(a[319] & b[102])^(a[318] & b[103])^(a[317] & b[104])^(a[316] & b[105])^(a[315] & b[106])^(a[314] & b[107])^(a[313] & b[108])^(a[312] & b[109])^(a[311] & b[110])^(a[310] & b[111])^(a[309] & b[112])^(a[308] & b[113])^(a[307] & b[114])^(a[306] & b[115])^(a[305] & b[116])^(a[304] & b[117])^(a[303] & b[118])^(a[302] & b[119])^(a[301] & b[120])^(a[300] & b[121])^(a[299] & b[122])^(a[298] & b[123])^(a[297] & b[124])^(a[296] & b[125])^(a[295] & b[126])^(a[294] & b[127])^(a[293] & b[128])^(a[292] & b[129])^(a[291] & b[130])^(a[290] & b[131])^(a[289] & b[132])^(a[288] & b[133])^(a[287] & b[134])^(a[286] & b[135])^(a[285] & b[136])^(a[284] & b[137])^(a[283] & b[138])^(a[282] & b[139])^(a[281] & b[140])^(a[280] & b[141])^(a[279] & b[142])^(a[278] & b[143])^(a[277] & b[144])^(a[276] & b[145])^(a[275] & b[146])^(a[274] & b[147])^(a[273] & b[148])^(a[272] & b[149])^(a[271] & b[150])^(a[270] & b[151])^(a[269] & b[152])^(a[268] & b[153])^(a[267] & b[154])^(a[266] & b[155])^(a[265] & b[156])^(a[264] & b[157])^(a[263] & b[158])^(a[262] & b[159])^(a[261] & b[160])^(a[260] & b[161])^(a[259] & b[162])^(a[258] & b[163])^(a[257] & b[164])^(a[256] & b[165])^(a[255] & b[166])^(a[254] & b[167])^(a[253] & b[168])^(a[252] & b[169])^(a[251] & b[170])^(a[250] & b[171])^(a[249] & b[172])^(a[248] & b[173])^(a[247] & b[174])^(a[246] & b[175])^(a[245] & b[176])^(a[244] & b[177])^(a[243] & b[178])^(a[242] & b[179])^(a[241] & b[180])^(a[240] & b[181])^(a[239] & b[182])^(a[238] & b[183])^(a[237] & b[184])^(a[236] & b[185])^(a[235] & b[186])^(a[234] & b[187])^(a[233] & b[188])^(a[232] & b[189])^(a[231] & b[190])^(a[230] & b[191])^(a[229] & b[192])^(a[228] & b[193])^(a[227] & b[194])^(a[226] & b[195])^(a[225] & b[196])^(a[224] & b[197])^(a[223] & b[198])^(a[222] & b[199])^(a[221] & b[200])^(a[220] & b[201])^(a[219] & b[202])^(a[218] & b[203])^(a[217] & b[204])^(a[216] & b[205])^(a[215] & b[206])^(a[214] & b[207])^(a[213] & b[208])^(a[212] & b[209])^(a[211] & b[210])^(a[210] & b[211])^(a[209] & b[212])^(a[208] & b[213])^(a[207] & b[214])^(a[206] & b[215])^(a[205] & b[216])^(a[204] & b[217])^(a[203] & b[218])^(a[202] & b[219])^(a[201] & b[220])^(a[200] & b[221])^(a[199] & b[222])^(a[198] & b[223])^(a[197] & b[224])^(a[196] & b[225])^(a[195] & b[226])^(a[194] & b[227])^(a[193] & b[228])^(a[192] & b[229])^(a[191] & b[230])^(a[190] & b[231])^(a[189] & b[232])^(a[188] & b[233])^(a[187] & b[234])^(a[186] & b[235])^(a[185] & b[236])^(a[184] & b[237])^(a[183] & b[238])^(a[182] & b[239])^(a[181] & b[240])^(a[180] & b[241])^(a[179] & b[242])^(a[178] & b[243])^(a[177] & b[244])^(a[176] & b[245])^(a[175] & b[246])^(a[174] & b[247])^(a[173] & b[248])^(a[172] & b[249])^(a[171] & b[250])^(a[170] & b[251])^(a[169] & b[252])^(a[168] & b[253])^(a[167] & b[254])^(a[166] & b[255])^(a[165] & b[256])^(a[164] & b[257])^(a[163] & b[258])^(a[162] & b[259])^(a[161] & b[260])^(a[160] & b[261])^(a[159] & b[262])^(a[158] & b[263])^(a[157] & b[264])^(a[156] & b[265])^(a[155] & b[266])^(a[154] & b[267])^(a[153] & b[268])^(a[152] & b[269])^(a[151] & b[270])^(a[150] & b[271])^(a[149] & b[272])^(a[148] & b[273])^(a[147] & b[274])^(a[146] & b[275])^(a[145] & b[276])^(a[144] & b[277])^(a[143] & b[278])^(a[142] & b[279])^(a[141] & b[280])^(a[140] & b[281])^(a[139] & b[282])^(a[138] & b[283])^(a[137] & b[284])^(a[136] & b[285])^(a[135] & b[286])^(a[134] & b[287])^(a[133] & b[288])^(a[132] & b[289])^(a[131] & b[290])^(a[130] & b[291])^(a[129] & b[292])^(a[128] & b[293])^(a[127] & b[294])^(a[126] & b[295])^(a[125] & b[296])^(a[124] & b[297])^(a[123] & b[298])^(a[122] & b[299])^(a[121] & b[300])^(a[120] & b[301])^(a[119] & b[302])^(a[118] & b[303])^(a[117] & b[304])^(a[116] & b[305])^(a[115] & b[306])^(a[114] & b[307])^(a[113] & b[308])^(a[112] & b[309])^(a[111] & b[310])^(a[110] & b[311])^(a[109] & b[312])^(a[108] & b[313])^(a[107] & b[314])^(a[106] & b[315])^(a[105] & b[316])^(a[104] & b[317])^(a[103] & b[318])^(a[102] & b[319])^(a[101] & b[320])^(a[100] & b[321])^(a[99] & b[322])^(a[98] & b[323])^(a[97] & b[324])^(a[96] & b[325])^(a[95] & b[326])^(a[94] & b[327])^(a[93] & b[328])^(a[92] & b[329])^(a[91] & b[330])^(a[90] & b[331])^(a[89] & b[332])^(a[88] & b[333])^(a[87] & b[334])^(a[86] & b[335])^(a[85] & b[336])^(a[84] & b[337])^(a[83] & b[338])^(a[82] & b[339])^(a[81] & b[340])^(a[80] & b[341])^(a[79] & b[342])^(a[78] & b[343])^(a[77] & b[344])^(a[76] & b[345])^(a[75] & b[346])^(a[74] & b[347])^(a[73] & b[348])^(a[72] & b[349])^(a[71] & b[350])^(a[70] & b[351])^(a[69] & b[352])^(a[68] & b[353])^(a[67] & b[354])^(a[66] & b[355])^(a[65] & b[356])^(a[64] & b[357])^(a[63] & b[358])^(a[62] & b[359])^(a[61] & b[360])^(a[60] & b[361])^(a[59] & b[362])^(a[58] & b[363])^(a[57] & b[364])^(a[56] & b[365])^(a[55] & b[366])^(a[54] & b[367])^(a[53] & b[368])^(a[52] & b[369])^(a[51] & b[370])^(a[50] & b[371])^(a[49] & b[372])^(a[48] & b[373])^(a[47] & b[374])^(a[46] & b[375])^(a[45] & b[376])^(a[44] & b[377])^(a[43] & b[378])^(a[42] & b[379])^(a[41] & b[380])^(a[40] & b[381])^(a[39] & b[382])^(a[38] & b[383])^(a[37] & b[384])^(a[36] & b[385])^(a[35] & b[386])^(a[34] & b[387])^(a[33] & b[388])^(a[32] & b[389])^(a[31] & b[390])^(a[30] & b[391])^(a[29] & b[392])^(a[28] & b[393])^(a[27] & b[394])^(a[26] & b[395])^(a[25] & b[396])^(a[24] & b[397])^(a[23] & b[398])^(a[22] & b[399])^(a[21] & b[400])^(a[20] & b[401])^(a[19] & b[402])^(a[18] & b[403])^(a[17] & b[404])^(a[16] & b[405])^(a[15] & b[406])^(a[14] & b[407])^(a[13] & b[408]);
assign y[422] = (a[408] & b[14])^(a[407] & b[15])^(a[406] & b[16])^(a[405] & b[17])^(a[404] & b[18])^(a[403] & b[19])^(a[402] & b[20])^(a[401] & b[21])^(a[400] & b[22])^(a[399] & b[23])^(a[398] & b[24])^(a[397] & b[25])^(a[396] & b[26])^(a[395] & b[27])^(a[394] & b[28])^(a[393] & b[29])^(a[392] & b[30])^(a[391] & b[31])^(a[390] & b[32])^(a[389] & b[33])^(a[388] & b[34])^(a[387] & b[35])^(a[386] & b[36])^(a[385] & b[37])^(a[384] & b[38])^(a[383] & b[39])^(a[382] & b[40])^(a[381] & b[41])^(a[380] & b[42])^(a[379] & b[43])^(a[378] & b[44])^(a[377] & b[45])^(a[376] & b[46])^(a[375] & b[47])^(a[374] & b[48])^(a[373] & b[49])^(a[372] & b[50])^(a[371] & b[51])^(a[370] & b[52])^(a[369] & b[53])^(a[368] & b[54])^(a[367] & b[55])^(a[366] & b[56])^(a[365] & b[57])^(a[364] & b[58])^(a[363] & b[59])^(a[362] & b[60])^(a[361] & b[61])^(a[360] & b[62])^(a[359] & b[63])^(a[358] & b[64])^(a[357] & b[65])^(a[356] & b[66])^(a[355] & b[67])^(a[354] & b[68])^(a[353] & b[69])^(a[352] & b[70])^(a[351] & b[71])^(a[350] & b[72])^(a[349] & b[73])^(a[348] & b[74])^(a[347] & b[75])^(a[346] & b[76])^(a[345] & b[77])^(a[344] & b[78])^(a[343] & b[79])^(a[342] & b[80])^(a[341] & b[81])^(a[340] & b[82])^(a[339] & b[83])^(a[338] & b[84])^(a[337] & b[85])^(a[336] & b[86])^(a[335] & b[87])^(a[334] & b[88])^(a[333] & b[89])^(a[332] & b[90])^(a[331] & b[91])^(a[330] & b[92])^(a[329] & b[93])^(a[328] & b[94])^(a[327] & b[95])^(a[326] & b[96])^(a[325] & b[97])^(a[324] & b[98])^(a[323] & b[99])^(a[322] & b[100])^(a[321] & b[101])^(a[320] & b[102])^(a[319] & b[103])^(a[318] & b[104])^(a[317] & b[105])^(a[316] & b[106])^(a[315] & b[107])^(a[314] & b[108])^(a[313] & b[109])^(a[312] & b[110])^(a[311] & b[111])^(a[310] & b[112])^(a[309] & b[113])^(a[308] & b[114])^(a[307] & b[115])^(a[306] & b[116])^(a[305] & b[117])^(a[304] & b[118])^(a[303] & b[119])^(a[302] & b[120])^(a[301] & b[121])^(a[300] & b[122])^(a[299] & b[123])^(a[298] & b[124])^(a[297] & b[125])^(a[296] & b[126])^(a[295] & b[127])^(a[294] & b[128])^(a[293] & b[129])^(a[292] & b[130])^(a[291] & b[131])^(a[290] & b[132])^(a[289] & b[133])^(a[288] & b[134])^(a[287] & b[135])^(a[286] & b[136])^(a[285] & b[137])^(a[284] & b[138])^(a[283] & b[139])^(a[282] & b[140])^(a[281] & b[141])^(a[280] & b[142])^(a[279] & b[143])^(a[278] & b[144])^(a[277] & b[145])^(a[276] & b[146])^(a[275] & b[147])^(a[274] & b[148])^(a[273] & b[149])^(a[272] & b[150])^(a[271] & b[151])^(a[270] & b[152])^(a[269] & b[153])^(a[268] & b[154])^(a[267] & b[155])^(a[266] & b[156])^(a[265] & b[157])^(a[264] & b[158])^(a[263] & b[159])^(a[262] & b[160])^(a[261] & b[161])^(a[260] & b[162])^(a[259] & b[163])^(a[258] & b[164])^(a[257] & b[165])^(a[256] & b[166])^(a[255] & b[167])^(a[254] & b[168])^(a[253] & b[169])^(a[252] & b[170])^(a[251] & b[171])^(a[250] & b[172])^(a[249] & b[173])^(a[248] & b[174])^(a[247] & b[175])^(a[246] & b[176])^(a[245] & b[177])^(a[244] & b[178])^(a[243] & b[179])^(a[242] & b[180])^(a[241] & b[181])^(a[240] & b[182])^(a[239] & b[183])^(a[238] & b[184])^(a[237] & b[185])^(a[236] & b[186])^(a[235] & b[187])^(a[234] & b[188])^(a[233] & b[189])^(a[232] & b[190])^(a[231] & b[191])^(a[230] & b[192])^(a[229] & b[193])^(a[228] & b[194])^(a[227] & b[195])^(a[226] & b[196])^(a[225] & b[197])^(a[224] & b[198])^(a[223] & b[199])^(a[222] & b[200])^(a[221] & b[201])^(a[220] & b[202])^(a[219] & b[203])^(a[218] & b[204])^(a[217] & b[205])^(a[216] & b[206])^(a[215] & b[207])^(a[214] & b[208])^(a[213] & b[209])^(a[212] & b[210])^(a[211] & b[211])^(a[210] & b[212])^(a[209] & b[213])^(a[208] & b[214])^(a[207] & b[215])^(a[206] & b[216])^(a[205] & b[217])^(a[204] & b[218])^(a[203] & b[219])^(a[202] & b[220])^(a[201] & b[221])^(a[200] & b[222])^(a[199] & b[223])^(a[198] & b[224])^(a[197] & b[225])^(a[196] & b[226])^(a[195] & b[227])^(a[194] & b[228])^(a[193] & b[229])^(a[192] & b[230])^(a[191] & b[231])^(a[190] & b[232])^(a[189] & b[233])^(a[188] & b[234])^(a[187] & b[235])^(a[186] & b[236])^(a[185] & b[237])^(a[184] & b[238])^(a[183] & b[239])^(a[182] & b[240])^(a[181] & b[241])^(a[180] & b[242])^(a[179] & b[243])^(a[178] & b[244])^(a[177] & b[245])^(a[176] & b[246])^(a[175] & b[247])^(a[174] & b[248])^(a[173] & b[249])^(a[172] & b[250])^(a[171] & b[251])^(a[170] & b[252])^(a[169] & b[253])^(a[168] & b[254])^(a[167] & b[255])^(a[166] & b[256])^(a[165] & b[257])^(a[164] & b[258])^(a[163] & b[259])^(a[162] & b[260])^(a[161] & b[261])^(a[160] & b[262])^(a[159] & b[263])^(a[158] & b[264])^(a[157] & b[265])^(a[156] & b[266])^(a[155] & b[267])^(a[154] & b[268])^(a[153] & b[269])^(a[152] & b[270])^(a[151] & b[271])^(a[150] & b[272])^(a[149] & b[273])^(a[148] & b[274])^(a[147] & b[275])^(a[146] & b[276])^(a[145] & b[277])^(a[144] & b[278])^(a[143] & b[279])^(a[142] & b[280])^(a[141] & b[281])^(a[140] & b[282])^(a[139] & b[283])^(a[138] & b[284])^(a[137] & b[285])^(a[136] & b[286])^(a[135] & b[287])^(a[134] & b[288])^(a[133] & b[289])^(a[132] & b[290])^(a[131] & b[291])^(a[130] & b[292])^(a[129] & b[293])^(a[128] & b[294])^(a[127] & b[295])^(a[126] & b[296])^(a[125] & b[297])^(a[124] & b[298])^(a[123] & b[299])^(a[122] & b[300])^(a[121] & b[301])^(a[120] & b[302])^(a[119] & b[303])^(a[118] & b[304])^(a[117] & b[305])^(a[116] & b[306])^(a[115] & b[307])^(a[114] & b[308])^(a[113] & b[309])^(a[112] & b[310])^(a[111] & b[311])^(a[110] & b[312])^(a[109] & b[313])^(a[108] & b[314])^(a[107] & b[315])^(a[106] & b[316])^(a[105] & b[317])^(a[104] & b[318])^(a[103] & b[319])^(a[102] & b[320])^(a[101] & b[321])^(a[100] & b[322])^(a[99] & b[323])^(a[98] & b[324])^(a[97] & b[325])^(a[96] & b[326])^(a[95] & b[327])^(a[94] & b[328])^(a[93] & b[329])^(a[92] & b[330])^(a[91] & b[331])^(a[90] & b[332])^(a[89] & b[333])^(a[88] & b[334])^(a[87] & b[335])^(a[86] & b[336])^(a[85] & b[337])^(a[84] & b[338])^(a[83] & b[339])^(a[82] & b[340])^(a[81] & b[341])^(a[80] & b[342])^(a[79] & b[343])^(a[78] & b[344])^(a[77] & b[345])^(a[76] & b[346])^(a[75] & b[347])^(a[74] & b[348])^(a[73] & b[349])^(a[72] & b[350])^(a[71] & b[351])^(a[70] & b[352])^(a[69] & b[353])^(a[68] & b[354])^(a[67] & b[355])^(a[66] & b[356])^(a[65] & b[357])^(a[64] & b[358])^(a[63] & b[359])^(a[62] & b[360])^(a[61] & b[361])^(a[60] & b[362])^(a[59] & b[363])^(a[58] & b[364])^(a[57] & b[365])^(a[56] & b[366])^(a[55] & b[367])^(a[54] & b[368])^(a[53] & b[369])^(a[52] & b[370])^(a[51] & b[371])^(a[50] & b[372])^(a[49] & b[373])^(a[48] & b[374])^(a[47] & b[375])^(a[46] & b[376])^(a[45] & b[377])^(a[44] & b[378])^(a[43] & b[379])^(a[42] & b[380])^(a[41] & b[381])^(a[40] & b[382])^(a[39] & b[383])^(a[38] & b[384])^(a[37] & b[385])^(a[36] & b[386])^(a[35] & b[387])^(a[34] & b[388])^(a[33] & b[389])^(a[32] & b[390])^(a[31] & b[391])^(a[30] & b[392])^(a[29] & b[393])^(a[28] & b[394])^(a[27] & b[395])^(a[26] & b[396])^(a[25] & b[397])^(a[24] & b[398])^(a[23] & b[399])^(a[22] & b[400])^(a[21] & b[401])^(a[20] & b[402])^(a[19] & b[403])^(a[18] & b[404])^(a[17] & b[405])^(a[16] & b[406])^(a[15] & b[407])^(a[14] & b[408]);
assign y[423] = (a[408] & b[15])^(a[407] & b[16])^(a[406] & b[17])^(a[405] & b[18])^(a[404] & b[19])^(a[403] & b[20])^(a[402] & b[21])^(a[401] & b[22])^(a[400] & b[23])^(a[399] & b[24])^(a[398] & b[25])^(a[397] & b[26])^(a[396] & b[27])^(a[395] & b[28])^(a[394] & b[29])^(a[393] & b[30])^(a[392] & b[31])^(a[391] & b[32])^(a[390] & b[33])^(a[389] & b[34])^(a[388] & b[35])^(a[387] & b[36])^(a[386] & b[37])^(a[385] & b[38])^(a[384] & b[39])^(a[383] & b[40])^(a[382] & b[41])^(a[381] & b[42])^(a[380] & b[43])^(a[379] & b[44])^(a[378] & b[45])^(a[377] & b[46])^(a[376] & b[47])^(a[375] & b[48])^(a[374] & b[49])^(a[373] & b[50])^(a[372] & b[51])^(a[371] & b[52])^(a[370] & b[53])^(a[369] & b[54])^(a[368] & b[55])^(a[367] & b[56])^(a[366] & b[57])^(a[365] & b[58])^(a[364] & b[59])^(a[363] & b[60])^(a[362] & b[61])^(a[361] & b[62])^(a[360] & b[63])^(a[359] & b[64])^(a[358] & b[65])^(a[357] & b[66])^(a[356] & b[67])^(a[355] & b[68])^(a[354] & b[69])^(a[353] & b[70])^(a[352] & b[71])^(a[351] & b[72])^(a[350] & b[73])^(a[349] & b[74])^(a[348] & b[75])^(a[347] & b[76])^(a[346] & b[77])^(a[345] & b[78])^(a[344] & b[79])^(a[343] & b[80])^(a[342] & b[81])^(a[341] & b[82])^(a[340] & b[83])^(a[339] & b[84])^(a[338] & b[85])^(a[337] & b[86])^(a[336] & b[87])^(a[335] & b[88])^(a[334] & b[89])^(a[333] & b[90])^(a[332] & b[91])^(a[331] & b[92])^(a[330] & b[93])^(a[329] & b[94])^(a[328] & b[95])^(a[327] & b[96])^(a[326] & b[97])^(a[325] & b[98])^(a[324] & b[99])^(a[323] & b[100])^(a[322] & b[101])^(a[321] & b[102])^(a[320] & b[103])^(a[319] & b[104])^(a[318] & b[105])^(a[317] & b[106])^(a[316] & b[107])^(a[315] & b[108])^(a[314] & b[109])^(a[313] & b[110])^(a[312] & b[111])^(a[311] & b[112])^(a[310] & b[113])^(a[309] & b[114])^(a[308] & b[115])^(a[307] & b[116])^(a[306] & b[117])^(a[305] & b[118])^(a[304] & b[119])^(a[303] & b[120])^(a[302] & b[121])^(a[301] & b[122])^(a[300] & b[123])^(a[299] & b[124])^(a[298] & b[125])^(a[297] & b[126])^(a[296] & b[127])^(a[295] & b[128])^(a[294] & b[129])^(a[293] & b[130])^(a[292] & b[131])^(a[291] & b[132])^(a[290] & b[133])^(a[289] & b[134])^(a[288] & b[135])^(a[287] & b[136])^(a[286] & b[137])^(a[285] & b[138])^(a[284] & b[139])^(a[283] & b[140])^(a[282] & b[141])^(a[281] & b[142])^(a[280] & b[143])^(a[279] & b[144])^(a[278] & b[145])^(a[277] & b[146])^(a[276] & b[147])^(a[275] & b[148])^(a[274] & b[149])^(a[273] & b[150])^(a[272] & b[151])^(a[271] & b[152])^(a[270] & b[153])^(a[269] & b[154])^(a[268] & b[155])^(a[267] & b[156])^(a[266] & b[157])^(a[265] & b[158])^(a[264] & b[159])^(a[263] & b[160])^(a[262] & b[161])^(a[261] & b[162])^(a[260] & b[163])^(a[259] & b[164])^(a[258] & b[165])^(a[257] & b[166])^(a[256] & b[167])^(a[255] & b[168])^(a[254] & b[169])^(a[253] & b[170])^(a[252] & b[171])^(a[251] & b[172])^(a[250] & b[173])^(a[249] & b[174])^(a[248] & b[175])^(a[247] & b[176])^(a[246] & b[177])^(a[245] & b[178])^(a[244] & b[179])^(a[243] & b[180])^(a[242] & b[181])^(a[241] & b[182])^(a[240] & b[183])^(a[239] & b[184])^(a[238] & b[185])^(a[237] & b[186])^(a[236] & b[187])^(a[235] & b[188])^(a[234] & b[189])^(a[233] & b[190])^(a[232] & b[191])^(a[231] & b[192])^(a[230] & b[193])^(a[229] & b[194])^(a[228] & b[195])^(a[227] & b[196])^(a[226] & b[197])^(a[225] & b[198])^(a[224] & b[199])^(a[223] & b[200])^(a[222] & b[201])^(a[221] & b[202])^(a[220] & b[203])^(a[219] & b[204])^(a[218] & b[205])^(a[217] & b[206])^(a[216] & b[207])^(a[215] & b[208])^(a[214] & b[209])^(a[213] & b[210])^(a[212] & b[211])^(a[211] & b[212])^(a[210] & b[213])^(a[209] & b[214])^(a[208] & b[215])^(a[207] & b[216])^(a[206] & b[217])^(a[205] & b[218])^(a[204] & b[219])^(a[203] & b[220])^(a[202] & b[221])^(a[201] & b[222])^(a[200] & b[223])^(a[199] & b[224])^(a[198] & b[225])^(a[197] & b[226])^(a[196] & b[227])^(a[195] & b[228])^(a[194] & b[229])^(a[193] & b[230])^(a[192] & b[231])^(a[191] & b[232])^(a[190] & b[233])^(a[189] & b[234])^(a[188] & b[235])^(a[187] & b[236])^(a[186] & b[237])^(a[185] & b[238])^(a[184] & b[239])^(a[183] & b[240])^(a[182] & b[241])^(a[181] & b[242])^(a[180] & b[243])^(a[179] & b[244])^(a[178] & b[245])^(a[177] & b[246])^(a[176] & b[247])^(a[175] & b[248])^(a[174] & b[249])^(a[173] & b[250])^(a[172] & b[251])^(a[171] & b[252])^(a[170] & b[253])^(a[169] & b[254])^(a[168] & b[255])^(a[167] & b[256])^(a[166] & b[257])^(a[165] & b[258])^(a[164] & b[259])^(a[163] & b[260])^(a[162] & b[261])^(a[161] & b[262])^(a[160] & b[263])^(a[159] & b[264])^(a[158] & b[265])^(a[157] & b[266])^(a[156] & b[267])^(a[155] & b[268])^(a[154] & b[269])^(a[153] & b[270])^(a[152] & b[271])^(a[151] & b[272])^(a[150] & b[273])^(a[149] & b[274])^(a[148] & b[275])^(a[147] & b[276])^(a[146] & b[277])^(a[145] & b[278])^(a[144] & b[279])^(a[143] & b[280])^(a[142] & b[281])^(a[141] & b[282])^(a[140] & b[283])^(a[139] & b[284])^(a[138] & b[285])^(a[137] & b[286])^(a[136] & b[287])^(a[135] & b[288])^(a[134] & b[289])^(a[133] & b[290])^(a[132] & b[291])^(a[131] & b[292])^(a[130] & b[293])^(a[129] & b[294])^(a[128] & b[295])^(a[127] & b[296])^(a[126] & b[297])^(a[125] & b[298])^(a[124] & b[299])^(a[123] & b[300])^(a[122] & b[301])^(a[121] & b[302])^(a[120] & b[303])^(a[119] & b[304])^(a[118] & b[305])^(a[117] & b[306])^(a[116] & b[307])^(a[115] & b[308])^(a[114] & b[309])^(a[113] & b[310])^(a[112] & b[311])^(a[111] & b[312])^(a[110] & b[313])^(a[109] & b[314])^(a[108] & b[315])^(a[107] & b[316])^(a[106] & b[317])^(a[105] & b[318])^(a[104] & b[319])^(a[103] & b[320])^(a[102] & b[321])^(a[101] & b[322])^(a[100] & b[323])^(a[99] & b[324])^(a[98] & b[325])^(a[97] & b[326])^(a[96] & b[327])^(a[95] & b[328])^(a[94] & b[329])^(a[93] & b[330])^(a[92] & b[331])^(a[91] & b[332])^(a[90] & b[333])^(a[89] & b[334])^(a[88] & b[335])^(a[87] & b[336])^(a[86] & b[337])^(a[85] & b[338])^(a[84] & b[339])^(a[83] & b[340])^(a[82] & b[341])^(a[81] & b[342])^(a[80] & b[343])^(a[79] & b[344])^(a[78] & b[345])^(a[77] & b[346])^(a[76] & b[347])^(a[75] & b[348])^(a[74] & b[349])^(a[73] & b[350])^(a[72] & b[351])^(a[71] & b[352])^(a[70] & b[353])^(a[69] & b[354])^(a[68] & b[355])^(a[67] & b[356])^(a[66] & b[357])^(a[65] & b[358])^(a[64] & b[359])^(a[63] & b[360])^(a[62] & b[361])^(a[61] & b[362])^(a[60] & b[363])^(a[59] & b[364])^(a[58] & b[365])^(a[57] & b[366])^(a[56] & b[367])^(a[55] & b[368])^(a[54] & b[369])^(a[53] & b[370])^(a[52] & b[371])^(a[51] & b[372])^(a[50] & b[373])^(a[49] & b[374])^(a[48] & b[375])^(a[47] & b[376])^(a[46] & b[377])^(a[45] & b[378])^(a[44] & b[379])^(a[43] & b[380])^(a[42] & b[381])^(a[41] & b[382])^(a[40] & b[383])^(a[39] & b[384])^(a[38] & b[385])^(a[37] & b[386])^(a[36] & b[387])^(a[35] & b[388])^(a[34] & b[389])^(a[33] & b[390])^(a[32] & b[391])^(a[31] & b[392])^(a[30] & b[393])^(a[29] & b[394])^(a[28] & b[395])^(a[27] & b[396])^(a[26] & b[397])^(a[25] & b[398])^(a[24] & b[399])^(a[23] & b[400])^(a[22] & b[401])^(a[21] & b[402])^(a[20] & b[403])^(a[19] & b[404])^(a[18] & b[405])^(a[17] & b[406])^(a[16] & b[407])^(a[15] & b[408]);
assign y[424] = (a[408] & b[16])^(a[407] & b[17])^(a[406] & b[18])^(a[405] & b[19])^(a[404] & b[20])^(a[403] & b[21])^(a[402] & b[22])^(a[401] & b[23])^(a[400] & b[24])^(a[399] & b[25])^(a[398] & b[26])^(a[397] & b[27])^(a[396] & b[28])^(a[395] & b[29])^(a[394] & b[30])^(a[393] & b[31])^(a[392] & b[32])^(a[391] & b[33])^(a[390] & b[34])^(a[389] & b[35])^(a[388] & b[36])^(a[387] & b[37])^(a[386] & b[38])^(a[385] & b[39])^(a[384] & b[40])^(a[383] & b[41])^(a[382] & b[42])^(a[381] & b[43])^(a[380] & b[44])^(a[379] & b[45])^(a[378] & b[46])^(a[377] & b[47])^(a[376] & b[48])^(a[375] & b[49])^(a[374] & b[50])^(a[373] & b[51])^(a[372] & b[52])^(a[371] & b[53])^(a[370] & b[54])^(a[369] & b[55])^(a[368] & b[56])^(a[367] & b[57])^(a[366] & b[58])^(a[365] & b[59])^(a[364] & b[60])^(a[363] & b[61])^(a[362] & b[62])^(a[361] & b[63])^(a[360] & b[64])^(a[359] & b[65])^(a[358] & b[66])^(a[357] & b[67])^(a[356] & b[68])^(a[355] & b[69])^(a[354] & b[70])^(a[353] & b[71])^(a[352] & b[72])^(a[351] & b[73])^(a[350] & b[74])^(a[349] & b[75])^(a[348] & b[76])^(a[347] & b[77])^(a[346] & b[78])^(a[345] & b[79])^(a[344] & b[80])^(a[343] & b[81])^(a[342] & b[82])^(a[341] & b[83])^(a[340] & b[84])^(a[339] & b[85])^(a[338] & b[86])^(a[337] & b[87])^(a[336] & b[88])^(a[335] & b[89])^(a[334] & b[90])^(a[333] & b[91])^(a[332] & b[92])^(a[331] & b[93])^(a[330] & b[94])^(a[329] & b[95])^(a[328] & b[96])^(a[327] & b[97])^(a[326] & b[98])^(a[325] & b[99])^(a[324] & b[100])^(a[323] & b[101])^(a[322] & b[102])^(a[321] & b[103])^(a[320] & b[104])^(a[319] & b[105])^(a[318] & b[106])^(a[317] & b[107])^(a[316] & b[108])^(a[315] & b[109])^(a[314] & b[110])^(a[313] & b[111])^(a[312] & b[112])^(a[311] & b[113])^(a[310] & b[114])^(a[309] & b[115])^(a[308] & b[116])^(a[307] & b[117])^(a[306] & b[118])^(a[305] & b[119])^(a[304] & b[120])^(a[303] & b[121])^(a[302] & b[122])^(a[301] & b[123])^(a[300] & b[124])^(a[299] & b[125])^(a[298] & b[126])^(a[297] & b[127])^(a[296] & b[128])^(a[295] & b[129])^(a[294] & b[130])^(a[293] & b[131])^(a[292] & b[132])^(a[291] & b[133])^(a[290] & b[134])^(a[289] & b[135])^(a[288] & b[136])^(a[287] & b[137])^(a[286] & b[138])^(a[285] & b[139])^(a[284] & b[140])^(a[283] & b[141])^(a[282] & b[142])^(a[281] & b[143])^(a[280] & b[144])^(a[279] & b[145])^(a[278] & b[146])^(a[277] & b[147])^(a[276] & b[148])^(a[275] & b[149])^(a[274] & b[150])^(a[273] & b[151])^(a[272] & b[152])^(a[271] & b[153])^(a[270] & b[154])^(a[269] & b[155])^(a[268] & b[156])^(a[267] & b[157])^(a[266] & b[158])^(a[265] & b[159])^(a[264] & b[160])^(a[263] & b[161])^(a[262] & b[162])^(a[261] & b[163])^(a[260] & b[164])^(a[259] & b[165])^(a[258] & b[166])^(a[257] & b[167])^(a[256] & b[168])^(a[255] & b[169])^(a[254] & b[170])^(a[253] & b[171])^(a[252] & b[172])^(a[251] & b[173])^(a[250] & b[174])^(a[249] & b[175])^(a[248] & b[176])^(a[247] & b[177])^(a[246] & b[178])^(a[245] & b[179])^(a[244] & b[180])^(a[243] & b[181])^(a[242] & b[182])^(a[241] & b[183])^(a[240] & b[184])^(a[239] & b[185])^(a[238] & b[186])^(a[237] & b[187])^(a[236] & b[188])^(a[235] & b[189])^(a[234] & b[190])^(a[233] & b[191])^(a[232] & b[192])^(a[231] & b[193])^(a[230] & b[194])^(a[229] & b[195])^(a[228] & b[196])^(a[227] & b[197])^(a[226] & b[198])^(a[225] & b[199])^(a[224] & b[200])^(a[223] & b[201])^(a[222] & b[202])^(a[221] & b[203])^(a[220] & b[204])^(a[219] & b[205])^(a[218] & b[206])^(a[217] & b[207])^(a[216] & b[208])^(a[215] & b[209])^(a[214] & b[210])^(a[213] & b[211])^(a[212] & b[212])^(a[211] & b[213])^(a[210] & b[214])^(a[209] & b[215])^(a[208] & b[216])^(a[207] & b[217])^(a[206] & b[218])^(a[205] & b[219])^(a[204] & b[220])^(a[203] & b[221])^(a[202] & b[222])^(a[201] & b[223])^(a[200] & b[224])^(a[199] & b[225])^(a[198] & b[226])^(a[197] & b[227])^(a[196] & b[228])^(a[195] & b[229])^(a[194] & b[230])^(a[193] & b[231])^(a[192] & b[232])^(a[191] & b[233])^(a[190] & b[234])^(a[189] & b[235])^(a[188] & b[236])^(a[187] & b[237])^(a[186] & b[238])^(a[185] & b[239])^(a[184] & b[240])^(a[183] & b[241])^(a[182] & b[242])^(a[181] & b[243])^(a[180] & b[244])^(a[179] & b[245])^(a[178] & b[246])^(a[177] & b[247])^(a[176] & b[248])^(a[175] & b[249])^(a[174] & b[250])^(a[173] & b[251])^(a[172] & b[252])^(a[171] & b[253])^(a[170] & b[254])^(a[169] & b[255])^(a[168] & b[256])^(a[167] & b[257])^(a[166] & b[258])^(a[165] & b[259])^(a[164] & b[260])^(a[163] & b[261])^(a[162] & b[262])^(a[161] & b[263])^(a[160] & b[264])^(a[159] & b[265])^(a[158] & b[266])^(a[157] & b[267])^(a[156] & b[268])^(a[155] & b[269])^(a[154] & b[270])^(a[153] & b[271])^(a[152] & b[272])^(a[151] & b[273])^(a[150] & b[274])^(a[149] & b[275])^(a[148] & b[276])^(a[147] & b[277])^(a[146] & b[278])^(a[145] & b[279])^(a[144] & b[280])^(a[143] & b[281])^(a[142] & b[282])^(a[141] & b[283])^(a[140] & b[284])^(a[139] & b[285])^(a[138] & b[286])^(a[137] & b[287])^(a[136] & b[288])^(a[135] & b[289])^(a[134] & b[290])^(a[133] & b[291])^(a[132] & b[292])^(a[131] & b[293])^(a[130] & b[294])^(a[129] & b[295])^(a[128] & b[296])^(a[127] & b[297])^(a[126] & b[298])^(a[125] & b[299])^(a[124] & b[300])^(a[123] & b[301])^(a[122] & b[302])^(a[121] & b[303])^(a[120] & b[304])^(a[119] & b[305])^(a[118] & b[306])^(a[117] & b[307])^(a[116] & b[308])^(a[115] & b[309])^(a[114] & b[310])^(a[113] & b[311])^(a[112] & b[312])^(a[111] & b[313])^(a[110] & b[314])^(a[109] & b[315])^(a[108] & b[316])^(a[107] & b[317])^(a[106] & b[318])^(a[105] & b[319])^(a[104] & b[320])^(a[103] & b[321])^(a[102] & b[322])^(a[101] & b[323])^(a[100] & b[324])^(a[99] & b[325])^(a[98] & b[326])^(a[97] & b[327])^(a[96] & b[328])^(a[95] & b[329])^(a[94] & b[330])^(a[93] & b[331])^(a[92] & b[332])^(a[91] & b[333])^(a[90] & b[334])^(a[89] & b[335])^(a[88] & b[336])^(a[87] & b[337])^(a[86] & b[338])^(a[85] & b[339])^(a[84] & b[340])^(a[83] & b[341])^(a[82] & b[342])^(a[81] & b[343])^(a[80] & b[344])^(a[79] & b[345])^(a[78] & b[346])^(a[77] & b[347])^(a[76] & b[348])^(a[75] & b[349])^(a[74] & b[350])^(a[73] & b[351])^(a[72] & b[352])^(a[71] & b[353])^(a[70] & b[354])^(a[69] & b[355])^(a[68] & b[356])^(a[67] & b[357])^(a[66] & b[358])^(a[65] & b[359])^(a[64] & b[360])^(a[63] & b[361])^(a[62] & b[362])^(a[61] & b[363])^(a[60] & b[364])^(a[59] & b[365])^(a[58] & b[366])^(a[57] & b[367])^(a[56] & b[368])^(a[55] & b[369])^(a[54] & b[370])^(a[53] & b[371])^(a[52] & b[372])^(a[51] & b[373])^(a[50] & b[374])^(a[49] & b[375])^(a[48] & b[376])^(a[47] & b[377])^(a[46] & b[378])^(a[45] & b[379])^(a[44] & b[380])^(a[43] & b[381])^(a[42] & b[382])^(a[41] & b[383])^(a[40] & b[384])^(a[39] & b[385])^(a[38] & b[386])^(a[37] & b[387])^(a[36] & b[388])^(a[35] & b[389])^(a[34] & b[390])^(a[33] & b[391])^(a[32] & b[392])^(a[31] & b[393])^(a[30] & b[394])^(a[29] & b[395])^(a[28] & b[396])^(a[27] & b[397])^(a[26] & b[398])^(a[25] & b[399])^(a[24] & b[400])^(a[23] & b[401])^(a[22] & b[402])^(a[21] & b[403])^(a[20] & b[404])^(a[19] & b[405])^(a[18] & b[406])^(a[17] & b[407])^(a[16] & b[408]);
assign y[425] = (a[408] & b[17])^(a[407] & b[18])^(a[406] & b[19])^(a[405] & b[20])^(a[404] & b[21])^(a[403] & b[22])^(a[402] & b[23])^(a[401] & b[24])^(a[400] & b[25])^(a[399] & b[26])^(a[398] & b[27])^(a[397] & b[28])^(a[396] & b[29])^(a[395] & b[30])^(a[394] & b[31])^(a[393] & b[32])^(a[392] & b[33])^(a[391] & b[34])^(a[390] & b[35])^(a[389] & b[36])^(a[388] & b[37])^(a[387] & b[38])^(a[386] & b[39])^(a[385] & b[40])^(a[384] & b[41])^(a[383] & b[42])^(a[382] & b[43])^(a[381] & b[44])^(a[380] & b[45])^(a[379] & b[46])^(a[378] & b[47])^(a[377] & b[48])^(a[376] & b[49])^(a[375] & b[50])^(a[374] & b[51])^(a[373] & b[52])^(a[372] & b[53])^(a[371] & b[54])^(a[370] & b[55])^(a[369] & b[56])^(a[368] & b[57])^(a[367] & b[58])^(a[366] & b[59])^(a[365] & b[60])^(a[364] & b[61])^(a[363] & b[62])^(a[362] & b[63])^(a[361] & b[64])^(a[360] & b[65])^(a[359] & b[66])^(a[358] & b[67])^(a[357] & b[68])^(a[356] & b[69])^(a[355] & b[70])^(a[354] & b[71])^(a[353] & b[72])^(a[352] & b[73])^(a[351] & b[74])^(a[350] & b[75])^(a[349] & b[76])^(a[348] & b[77])^(a[347] & b[78])^(a[346] & b[79])^(a[345] & b[80])^(a[344] & b[81])^(a[343] & b[82])^(a[342] & b[83])^(a[341] & b[84])^(a[340] & b[85])^(a[339] & b[86])^(a[338] & b[87])^(a[337] & b[88])^(a[336] & b[89])^(a[335] & b[90])^(a[334] & b[91])^(a[333] & b[92])^(a[332] & b[93])^(a[331] & b[94])^(a[330] & b[95])^(a[329] & b[96])^(a[328] & b[97])^(a[327] & b[98])^(a[326] & b[99])^(a[325] & b[100])^(a[324] & b[101])^(a[323] & b[102])^(a[322] & b[103])^(a[321] & b[104])^(a[320] & b[105])^(a[319] & b[106])^(a[318] & b[107])^(a[317] & b[108])^(a[316] & b[109])^(a[315] & b[110])^(a[314] & b[111])^(a[313] & b[112])^(a[312] & b[113])^(a[311] & b[114])^(a[310] & b[115])^(a[309] & b[116])^(a[308] & b[117])^(a[307] & b[118])^(a[306] & b[119])^(a[305] & b[120])^(a[304] & b[121])^(a[303] & b[122])^(a[302] & b[123])^(a[301] & b[124])^(a[300] & b[125])^(a[299] & b[126])^(a[298] & b[127])^(a[297] & b[128])^(a[296] & b[129])^(a[295] & b[130])^(a[294] & b[131])^(a[293] & b[132])^(a[292] & b[133])^(a[291] & b[134])^(a[290] & b[135])^(a[289] & b[136])^(a[288] & b[137])^(a[287] & b[138])^(a[286] & b[139])^(a[285] & b[140])^(a[284] & b[141])^(a[283] & b[142])^(a[282] & b[143])^(a[281] & b[144])^(a[280] & b[145])^(a[279] & b[146])^(a[278] & b[147])^(a[277] & b[148])^(a[276] & b[149])^(a[275] & b[150])^(a[274] & b[151])^(a[273] & b[152])^(a[272] & b[153])^(a[271] & b[154])^(a[270] & b[155])^(a[269] & b[156])^(a[268] & b[157])^(a[267] & b[158])^(a[266] & b[159])^(a[265] & b[160])^(a[264] & b[161])^(a[263] & b[162])^(a[262] & b[163])^(a[261] & b[164])^(a[260] & b[165])^(a[259] & b[166])^(a[258] & b[167])^(a[257] & b[168])^(a[256] & b[169])^(a[255] & b[170])^(a[254] & b[171])^(a[253] & b[172])^(a[252] & b[173])^(a[251] & b[174])^(a[250] & b[175])^(a[249] & b[176])^(a[248] & b[177])^(a[247] & b[178])^(a[246] & b[179])^(a[245] & b[180])^(a[244] & b[181])^(a[243] & b[182])^(a[242] & b[183])^(a[241] & b[184])^(a[240] & b[185])^(a[239] & b[186])^(a[238] & b[187])^(a[237] & b[188])^(a[236] & b[189])^(a[235] & b[190])^(a[234] & b[191])^(a[233] & b[192])^(a[232] & b[193])^(a[231] & b[194])^(a[230] & b[195])^(a[229] & b[196])^(a[228] & b[197])^(a[227] & b[198])^(a[226] & b[199])^(a[225] & b[200])^(a[224] & b[201])^(a[223] & b[202])^(a[222] & b[203])^(a[221] & b[204])^(a[220] & b[205])^(a[219] & b[206])^(a[218] & b[207])^(a[217] & b[208])^(a[216] & b[209])^(a[215] & b[210])^(a[214] & b[211])^(a[213] & b[212])^(a[212] & b[213])^(a[211] & b[214])^(a[210] & b[215])^(a[209] & b[216])^(a[208] & b[217])^(a[207] & b[218])^(a[206] & b[219])^(a[205] & b[220])^(a[204] & b[221])^(a[203] & b[222])^(a[202] & b[223])^(a[201] & b[224])^(a[200] & b[225])^(a[199] & b[226])^(a[198] & b[227])^(a[197] & b[228])^(a[196] & b[229])^(a[195] & b[230])^(a[194] & b[231])^(a[193] & b[232])^(a[192] & b[233])^(a[191] & b[234])^(a[190] & b[235])^(a[189] & b[236])^(a[188] & b[237])^(a[187] & b[238])^(a[186] & b[239])^(a[185] & b[240])^(a[184] & b[241])^(a[183] & b[242])^(a[182] & b[243])^(a[181] & b[244])^(a[180] & b[245])^(a[179] & b[246])^(a[178] & b[247])^(a[177] & b[248])^(a[176] & b[249])^(a[175] & b[250])^(a[174] & b[251])^(a[173] & b[252])^(a[172] & b[253])^(a[171] & b[254])^(a[170] & b[255])^(a[169] & b[256])^(a[168] & b[257])^(a[167] & b[258])^(a[166] & b[259])^(a[165] & b[260])^(a[164] & b[261])^(a[163] & b[262])^(a[162] & b[263])^(a[161] & b[264])^(a[160] & b[265])^(a[159] & b[266])^(a[158] & b[267])^(a[157] & b[268])^(a[156] & b[269])^(a[155] & b[270])^(a[154] & b[271])^(a[153] & b[272])^(a[152] & b[273])^(a[151] & b[274])^(a[150] & b[275])^(a[149] & b[276])^(a[148] & b[277])^(a[147] & b[278])^(a[146] & b[279])^(a[145] & b[280])^(a[144] & b[281])^(a[143] & b[282])^(a[142] & b[283])^(a[141] & b[284])^(a[140] & b[285])^(a[139] & b[286])^(a[138] & b[287])^(a[137] & b[288])^(a[136] & b[289])^(a[135] & b[290])^(a[134] & b[291])^(a[133] & b[292])^(a[132] & b[293])^(a[131] & b[294])^(a[130] & b[295])^(a[129] & b[296])^(a[128] & b[297])^(a[127] & b[298])^(a[126] & b[299])^(a[125] & b[300])^(a[124] & b[301])^(a[123] & b[302])^(a[122] & b[303])^(a[121] & b[304])^(a[120] & b[305])^(a[119] & b[306])^(a[118] & b[307])^(a[117] & b[308])^(a[116] & b[309])^(a[115] & b[310])^(a[114] & b[311])^(a[113] & b[312])^(a[112] & b[313])^(a[111] & b[314])^(a[110] & b[315])^(a[109] & b[316])^(a[108] & b[317])^(a[107] & b[318])^(a[106] & b[319])^(a[105] & b[320])^(a[104] & b[321])^(a[103] & b[322])^(a[102] & b[323])^(a[101] & b[324])^(a[100] & b[325])^(a[99] & b[326])^(a[98] & b[327])^(a[97] & b[328])^(a[96] & b[329])^(a[95] & b[330])^(a[94] & b[331])^(a[93] & b[332])^(a[92] & b[333])^(a[91] & b[334])^(a[90] & b[335])^(a[89] & b[336])^(a[88] & b[337])^(a[87] & b[338])^(a[86] & b[339])^(a[85] & b[340])^(a[84] & b[341])^(a[83] & b[342])^(a[82] & b[343])^(a[81] & b[344])^(a[80] & b[345])^(a[79] & b[346])^(a[78] & b[347])^(a[77] & b[348])^(a[76] & b[349])^(a[75] & b[350])^(a[74] & b[351])^(a[73] & b[352])^(a[72] & b[353])^(a[71] & b[354])^(a[70] & b[355])^(a[69] & b[356])^(a[68] & b[357])^(a[67] & b[358])^(a[66] & b[359])^(a[65] & b[360])^(a[64] & b[361])^(a[63] & b[362])^(a[62] & b[363])^(a[61] & b[364])^(a[60] & b[365])^(a[59] & b[366])^(a[58] & b[367])^(a[57] & b[368])^(a[56] & b[369])^(a[55] & b[370])^(a[54] & b[371])^(a[53] & b[372])^(a[52] & b[373])^(a[51] & b[374])^(a[50] & b[375])^(a[49] & b[376])^(a[48] & b[377])^(a[47] & b[378])^(a[46] & b[379])^(a[45] & b[380])^(a[44] & b[381])^(a[43] & b[382])^(a[42] & b[383])^(a[41] & b[384])^(a[40] & b[385])^(a[39] & b[386])^(a[38] & b[387])^(a[37] & b[388])^(a[36] & b[389])^(a[35] & b[390])^(a[34] & b[391])^(a[33] & b[392])^(a[32] & b[393])^(a[31] & b[394])^(a[30] & b[395])^(a[29] & b[396])^(a[28] & b[397])^(a[27] & b[398])^(a[26] & b[399])^(a[25] & b[400])^(a[24] & b[401])^(a[23] & b[402])^(a[22] & b[403])^(a[21] & b[404])^(a[20] & b[405])^(a[19] & b[406])^(a[18] & b[407])^(a[17] & b[408]);
assign y[426] = (a[408] & b[18])^(a[407] & b[19])^(a[406] & b[20])^(a[405] & b[21])^(a[404] & b[22])^(a[403] & b[23])^(a[402] & b[24])^(a[401] & b[25])^(a[400] & b[26])^(a[399] & b[27])^(a[398] & b[28])^(a[397] & b[29])^(a[396] & b[30])^(a[395] & b[31])^(a[394] & b[32])^(a[393] & b[33])^(a[392] & b[34])^(a[391] & b[35])^(a[390] & b[36])^(a[389] & b[37])^(a[388] & b[38])^(a[387] & b[39])^(a[386] & b[40])^(a[385] & b[41])^(a[384] & b[42])^(a[383] & b[43])^(a[382] & b[44])^(a[381] & b[45])^(a[380] & b[46])^(a[379] & b[47])^(a[378] & b[48])^(a[377] & b[49])^(a[376] & b[50])^(a[375] & b[51])^(a[374] & b[52])^(a[373] & b[53])^(a[372] & b[54])^(a[371] & b[55])^(a[370] & b[56])^(a[369] & b[57])^(a[368] & b[58])^(a[367] & b[59])^(a[366] & b[60])^(a[365] & b[61])^(a[364] & b[62])^(a[363] & b[63])^(a[362] & b[64])^(a[361] & b[65])^(a[360] & b[66])^(a[359] & b[67])^(a[358] & b[68])^(a[357] & b[69])^(a[356] & b[70])^(a[355] & b[71])^(a[354] & b[72])^(a[353] & b[73])^(a[352] & b[74])^(a[351] & b[75])^(a[350] & b[76])^(a[349] & b[77])^(a[348] & b[78])^(a[347] & b[79])^(a[346] & b[80])^(a[345] & b[81])^(a[344] & b[82])^(a[343] & b[83])^(a[342] & b[84])^(a[341] & b[85])^(a[340] & b[86])^(a[339] & b[87])^(a[338] & b[88])^(a[337] & b[89])^(a[336] & b[90])^(a[335] & b[91])^(a[334] & b[92])^(a[333] & b[93])^(a[332] & b[94])^(a[331] & b[95])^(a[330] & b[96])^(a[329] & b[97])^(a[328] & b[98])^(a[327] & b[99])^(a[326] & b[100])^(a[325] & b[101])^(a[324] & b[102])^(a[323] & b[103])^(a[322] & b[104])^(a[321] & b[105])^(a[320] & b[106])^(a[319] & b[107])^(a[318] & b[108])^(a[317] & b[109])^(a[316] & b[110])^(a[315] & b[111])^(a[314] & b[112])^(a[313] & b[113])^(a[312] & b[114])^(a[311] & b[115])^(a[310] & b[116])^(a[309] & b[117])^(a[308] & b[118])^(a[307] & b[119])^(a[306] & b[120])^(a[305] & b[121])^(a[304] & b[122])^(a[303] & b[123])^(a[302] & b[124])^(a[301] & b[125])^(a[300] & b[126])^(a[299] & b[127])^(a[298] & b[128])^(a[297] & b[129])^(a[296] & b[130])^(a[295] & b[131])^(a[294] & b[132])^(a[293] & b[133])^(a[292] & b[134])^(a[291] & b[135])^(a[290] & b[136])^(a[289] & b[137])^(a[288] & b[138])^(a[287] & b[139])^(a[286] & b[140])^(a[285] & b[141])^(a[284] & b[142])^(a[283] & b[143])^(a[282] & b[144])^(a[281] & b[145])^(a[280] & b[146])^(a[279] & b[147])^(a[278] & b[148])^(a[277] & b[149])^(a[276] & b[150])^(a[275] & b[151])^(a[274] & b[152])^(a[273] & b[153])^(a[272] & b[154])^(a[271] & b[155])^(a[270] & b[156])^(a[269] & b[157])^(a[268] & b[158])^(a[267] & b[159])^(a[266] & b[160])^(a[265] & b[161])^(a[264] & b[162])^(a[263] & b[163])^(a[262] & b[164])^(a[261] & b[165])^(a[260] & b[166])^(a[259] & b[167])^(a[258] & b[168])^(a[257] & b[169])^(a[256] & b[170])^(a[255] & b[171])^(a[254] & b[172])^(a[253] & b[173])^(a[252] & b[174])^(a[251] & b[175])^(a[250] & b[176])^(a[249] & b[177])^(a[248] & b[178])^(a[247] & b[179])^(a[246] & b[180])^(a[245] & b[181])^(a[244] & b[182])^(a[243] & b[183])^(a[242] & b[184])^(a[241] & b[185])^(a[240] & b[186])^(a[239] & b[187])^(a[238] & b[188])^(a[237] & b[189])^(a[236] & b[190])^(a[235] & b[191])^(a[234] & b[192])^(a[233] & b[193])^(a[232] & b[194])^(a[231] & b[195])^(a[230] & b[196])^(a[229] & b[197])^(a[228] & b[198])^(a[227] & b[199])^(a[226] & b[200])^(a[225] & b[201])^(a[224] & b[202])^(a[223] & b[203])^(a[222] & b[204])^(a[221] & b[205])^(a[220] & b[206])^(a[219] & b[207])^(a[218] & b[208])^(a[217] & b[209])^(a[216] & b[210])^(a[215] & b[211])^(a[214] & b[212])^(a[213] & b[213])^(a[212] & b[214])^(a[211] & b[215])^(a[210] & b[216])^(a[209] & b[217])^(a[208] & b[218])^(a[207] & b[219])^(a[206] & b[220])^(a[205] & b[221])^(a[204] & b[222])^(a[203] & b[223])^(a[202] & b[224])^(a[201] & b[225])^(a[200] & b[226])^(a[199] & b[227])^(a[198] & b[228])^(a[197] & b[229])^(a[196] & b[230])^(a[195] & b[231])^(a[194] & b[232])^(a[193] & b[233])^(a[192] & b[234])^(a[191] & b[235])^(a[190] & b[236])^(a[189] & b[237])^(a[188] & b[238])^(a[187] & b[239])^(a[186] & b[240])^(a[185] & b[241])^(a[184] & b[242])^(a[183] & b[243])^(a[182] & b[244])^(a[181] & b[245])^(a[180] & b[246])^(a[179] & b[247])^(a[178] & b[248])^(a[177] & b[249])^(a[176] & b[250])^(a[175] & b[251])^(a[174] & b[252])^(a[173] & b[253])^(a[172] & b[254])^(a[171] & b[255])^(a[170] & b[256])^(a[169] & b[257])^(a[168] & b[258])^(a[167] & b[259])^(a[166] & b[260])^(a[165] & b[261])^(a[164] & b[262])^(a[163] & b[263])^(a[162] & b[264])^(a[161] & b[265])^(a[160] & b[266])^(a[159] & b[267])^(a[158] & b[268])^(a[157] & b[269])^(a[156] & b[270])^(a[155] & b[271])^(a[154] & b[272])^(a[153] & b[273])^(a[152] & b[274])^(a[151] & b[275])^(a[150] & b[276])^(a[149] & b[277])^(a[148] & b[278])^(a[147] & b[279])^(a[146] & b[280])^(a[145] & b[281])^(a[144] & b[282])^(a[143] & b[283])^(a[142] & b[284])^(a[141] & b[285])^(a[140] & b[286])^(a[139] & b[287])^(a[138] & b[288])^(a[137] & b[289])^(a[136] & b[290])^(a[135] & b[291])^(a[134] & b[292])^(a[133] & b[293])^(a[132] & b[294])^(a[131] & b[295])^(a[130] & b[296])^(a[129] & b[297])^(a[128] & b[298])^(a[127] & b[299])^(a[126] & b[300])^(a[125] & b[301])^(a[124] & b[302])^(a[123] & b[303])^(a[122] & b[304])^(a[121] & b[305])^(a[120] & b[306])^(a[119] & b[307])^(a[118] & b[308])^(a[117] & b[309])^(a[116] & b[310])^(a[115] & b[311])^(a[114] & b[312])^(a[113] & b[313])^(a[112] & b[314])^(a[111] & b[315])^(a[110] & b[316])^(a[109] & b[317])^(a[108] & b[318])^(a[107] & b[319])^(a[106] & b[320])^(a[105] & b[321])^(a[104] & b[322])^(a[103] & b[323])^(a[102] & b[324])^(a[101] & b[325])^(a[100] & b[326])^(a[99] & b[327])^(a[98] & b[328])^(a[97] & b[329])^(a[96] & b[330])^(a[95] & b[331])^(a[94] & b[332])^(a[93] & b[333])^(a[92] & b[334])^(a[91] & b[335])^(a[90] & b[336])^(a[89] & b[337])^(a[88] & b[338])^(a[87] & b[339])^(a[86] & b[340])^(a[85] & b[341])^(a[84] & b[342])^(a[83] & b[343])^(a[82] & b[344])^(a[81] & b[345])^(a[80] & b[346])^(a[79] & b[347])^(a[78] & b[348])^(a[77] & b[349])^(a[76] & b[350])^(a[75] & b[351])^(a[74] & b[352])^(a[73] & b[353])^(a[72] & b[354])^(a[71] & b[355])^(a[70] & b[356])^(a[69] & b[357])^(a[68] & b[358])^(a[67] & b[359])^(a[66] & b[360])^(a[65] & b[361])^(a[64] & b[362])^(a[63] & b[363])^(a[62] & b[364])^(a[61] & b[365])^(a[60] & b[366])^(a[59] & b[367])^(a[58] & b[368])^(a[57] & b[369])^(a[56] & b[370])^(a[55] & b[371])^(a[54] & b[372])^(a[53] & b[373])^(a[52] & b[374])^(a[51] & b[375])^(a[50] & b[376])^(a[49] & b[377])^(a[48] & b[378])^(a[47] & b[379])^(a[46] & b[380])^(a[45] & b[381])^(a[44] & b[382])^(a[43] & b[383])^(a[42] & b[384])^(a[41] & b[385])^(a[40] & b[386])^(a[39] & b[387])^(a[38] & b[388])^(a[37] & b[389])^(a[36] & b[390])^(a[35] & b[391])^(a[34] & b[392])^(a[33] & b[393])^(a[32] & b[394])^(a[31] & b[395])^(a[30] & b[396])^(a[29] & b[397])^(a[28] & b[398])^(a[27] & b[399])^(a[26] & b[400])^(a[25] & b[401])^(a[24] & b[402])^(a[23] & b[403])^(a[22] & b[404])^(a[21] & b[405])^(a[20] & b[406])^(a[19] & b[407])^(a[18] & b[408]);
assign y[427] = (a[408] & b[19])^(a[407] & b[20])^(a[406] & b[21])^(a[405] & b[22])^(a[404] & b[23])^(a[403] & b[24])^(a[402] & b[25])^(a[401] & b[26])^(a[400] & b[27])^(a[399] & b[28])^(a[398] & b[29])^(a[397] & b[30])^(a[396] & b[31])^(a[395] & b[32])^(a[394] & b[33])^(a[393] & b[34])^(a[392] & b[35])^(a[391] & b[36])^(a[390] & b[37])^(a[389] & b[38])^(a[388] & b[39])^(a[387] & b[40])^(a[386] & b[41])^(a[385] & b[42])^(a[384] & b[43])^(a[383] & b[44])^(a[382] & b[45])^(a[381] & b[46])^(a[380] & b[47])^(a[379] & b[48])^(a[378] & b[49])^(a[377] & b[50])^(a[376] & b[51])^(a[375] & b[52])^(a[374] & b[53])^(a[373] & b[54])^(a[372] & b[55])^(a[371] & b[56])^(a[370] & b[57])^(a[369] & b[58])^(a[368] & b[59])^(a[367] & b[60])^(a[366] & b[61])^(a[365] & b[62])^(a[364] & b[63])^(a[363] & b[64])^(a[362] & b[65])^(a[361] & b[66])^(a[360] & b[67])^(a[359] & b[68])^(a[358] & b[69])^(a[357] & b[70])^(a[356] & b[71])^(a[355] & b[72])^(a[354] & b[73])^(a[353] & b[74])^(a[352] & b[75])^(a[351] & b[76])^(a[350] & b[77])^(a[349] & b[78])^(a[348] & b[79])^(a[347] & b[80])^(a[346] & b[81])^(a[345] & b[82])^(a[344] & b[83])^(a[343] & b[84])^(a[342] & b[85])^(a[341] & b[86])^(a[340] & b[87])^(a[339] & b[88])^(a[338] & b[89])^(a[337] & b[90])^(a[336] & b[91])^(a[335] & b[92])^(a[334] & b[93])^(a[333] & b[94])^(a[332] & b[95])^(a[331] & b[96])^(a[330] & b[97])^(a[329] & b[98])^(a[328] & b[99])^(a[327] & b[100])^(a[326] & b[101])^(a[325] & b[102])^(a[324] & b[103])^(a[323] & b[104])^(a[322] & b[105])^(a[321] & b[106])^(a[320] & b[107])^(a[319] & b[108])^(a[318] & b[109])^(a[317] & b[110])^(a[316] & b[111])^(a[315] & b[112])^(a[314] & b[113])^(a[313] & b[114])^(a[312] & b[115])^(a[311] & b[116])^(a[310] & b[117])^(a[309] & b[118])^(a[308] & b[119])^(a[307] & b[120])^(a[306] & b[121])^(a[305] & b[122])^(a[304] & b[123])^(a[303] & b[124])^(a[302] & b[125])^(a[301] & b[126])^(a[300] & b[127])^(a[299] & b[128])^(a[298] & b[129])^(a[297] & b[130])^(a[296] & b[131])^(a[295] & b[132])^(a[294] & b[133])^(a[293] & b[134])^(a[292] & b[135])^(a[291] & b[136])^(a[290] & b[137])^(a[289] & b[138])^(a[288] & b[139])^(a[287] & b[140])^(a[286] & b[141])^(a[285] & b[142])^(a[284] & b[143])^(a[283] & b[144])^(a[282] & b[145])^(a[281] & b[146])^(a[280] & b[147])^(a[279] & b[148])^(a[278] & b[149])^(a[277] & b[150])^(a[276] & b[151])^(a[275] & b[152])^(a[274] & b[153])^(a[273] & b[154])^(a[272] & b[155])^(a[271] & b[156])^(a[270] & b[157])^(a[269] & b[158])^(a[268] & b[159])^(a[267] & b[160])^(a[266] & b[161])^(a[265] & b[162])^(a[264] & b[163])^(a[263] & b[164])^(a[262] & b[165])^(a[261] & b[166])^(a[260] & b[167])^(a[259] & b[168])^(a[258] & b[169])^(a[257] & b[170])^(a[256] & b[171])^(a[255] & b[172])^(a[254] & b[173])^(a[253] & b[174])^(a[252] & b[175])^(a[251] & b[176])^(a[250] & b[177])^(a[249] & b[178])^(a[248] & b[179])^(a[247] & b[180])^(a[246] & b[181])^(a[245] & b[182])^(a[244] & b[183])^(a[243] & b[184])^(a[242] & b[185])^(a[241] & b[186])^(a[240] & b[187])^(a[239] & b[188])^(a[238] & b[189])^(a[237] & b[190])^(a[236] & b[191])^(a[235] & b[192])^(a[234] & b[193])^(a[233] & b[194])^(a[232] & b[195])^(a[231] & b[196])^(a[230] & b[197])^(a[229] & b[198])^(a[228] & b[199])^(a[227] & b[200])^(a[226] & b[201])^(a[225] & b[202])^(a[224] & b[203])^(a[223] & b[204])^(a[222] & b[205])^(a[221] & b[206])^(a[220] & b[207])^(a[219] & b[208])^(a[218] & b[209])^(a[217] & b[210])^(a[216] & b[211])^(a[215] & b[212])^(a[214] & b[213])^(a[213] & b[214])^(a[212] & b[215])^(a[211] & b[216])^(a[210] & b[217])^(a[209] & b[218])^(a[208] & b[219])^(a[207] & b[220])^(a[206] & b[221])^(a[205] & b[222])^(a[204] & b[223])^(a[203] & b[224])^(a[202] & b[225])^(a[201] & b[226])^(a[200] & b[227])^(a[199] & b[228])^(a[198] & b[229])^(a[197] & b[230])^(a[196] & b[231])^(a[195] & b[232])^(a[194] & b[233])^(a[193] & b[234])^(a[192] & b[235])^(a[191] & b[236])^(a[190] & b[237])^(a[189] & b[238])^(a[188] & b[239])^(a[187] & b[240])^(a[186] & b[241])^(a[185] & b[242])^(a[184] & b[243])^(a[183] & b[244])^(a[182] & b[245])^(a[181] & b[246])^(a[180] & b[247])^(a[179] & b[248])^(a[178] & b[249])^(a[177] & b[250])^(a[176] & b[251])^(a[175] & b[252])^(a[174] & b[253])^(a[173] & b[254])^(a[172] & b[255])^(a[171] & b[256])^(a[170] & b[257])^(a[169] & b[258])^(a[168] & b[259])^(a[167] & b[260])^(a[166] & b[261])^(a[165] & b[262])^(a[164] & b[263])^(a[163] & b[264])^(a[162] & b[265])^(a[161] & b[266])^(a[160] & b[267])^(a[159] & b[268])^(a[158] & b[269])^(a[157] & b[270])^(a[156] & b[271])^(a[155] & b[272])^(a[154] & b[273])^(a[153] & b[274])^(a[152] & b[275])^(a[151] & b[276])^(a[150] & b[277])^(a[149] & b[278])^(a[148] & b[279])^(a[147] & b[280])^(a[146] & b[281])^(a[145] & b[282])^(a[144] & b[283])^(a[143] & b[284])^(a[142] & b[285])^(a[141] & b[286])^(a[140] & b[287])^(a[139] & b[288])^(a[138] & b[289])^(a[137] & b[290])^(a[136] & b[291])^(a[135] & b[292])^(a[134] & b[293])^(a[133] & b[294])^(a[132] & b[295])^(a[131] & b[296])^(a[130] & b[297])^(a[129] & b[298])^(a[128] & b[299])^(a[127] & b[300])^(a[126] & b[301])^(a[125] & b[302])^(a[124] & b[303])^(a[123] & b[304])^(a[122] & b[305])^(a[121] & b[306])^(a[120] & b[307])^(a[119] & b[308])^(a[118] & b[309])^(a[117] & b[310])^(a[116] & b[311])^(a[115] & b[312])^(a[114] & b[313])^(a[113] & b[314])^(a[112] & b[315])^(a[111] & b[316])^(a[110] & b[317])^(a[109] & b[318])^(a[108] & b[319])^(a[107] & b[320])^(a[106] & b[321])^(a[105] & b[322])^(a[104] & b[323])^(a[103] & b[324])^(a[102] & b[325])^(a[101] & b[326])^(a[100] & b[327])^(a[99] & b[328])^(a[98] & b[329])^(a[97] & b[330])^(a[96] & b[331])^(a[95] & b[332])^(a[94] & b[333])^(a[93] & b[334])^(a[92] & b[335])^(a[91] & b[336])^(a[90] & b[337])^(a[89] & b[338])^(a[88] & b[339])^(a[87] & b[340])^(a[86] & b[341])^(a[85] & b[342])^(a[84] & b[343])^(a[83] & b[344])^(a[82] & b[345])^(a[81] & b[346])^(a[80] & b[347])^(a[79] & b[348])^(a[78] & b[349])^(a[77] & b[350])^(a[76] & b[351])^(a[75] & b[352])^(a[74] & b[353])^(a[73] & b[354])^(a[72] & b[355])^(a[71] & b[356])^(a[70] & b[357])^(a[69] & b[358])^(a[68] & b[359])^(a[67] & b[360])^(a[66] & b[361])^(a[65] & b[362])^(a[64] & b[363])^(a[63] & b[364])^(a[62] & b[365])^(a[61] & b[366])^(a[60] & b[367])^(a[59] & b[368])^(a[58] & b[369])^(a[57] & b[370])^(a[56] & b[371])^(a[55] & b[372])^(a[54] & b[373])^(a[53] & b[374])^(a[52] & b[375])^(a[51] & b[376])^(a[50] & b[377])^(a[49] & b[378])^(a[48] & b[379])^(a[47] & b[380])^(a[46] & b[381])^(a[45] & b[382])^(a[44] & b[383])^(a[43] & b[384])^(a[42] & b[385])^(a[41] & b[386])^(a[40] & b[387])^(a[39] & b[388])^(a[38] & b[389])^(a[37] & b[390])^(a[36] & b[391])^(a[35] & b[392])^(a[34] & b[393])^(a[33] & b[394])^(a[32] & b[395])^(a[31] & b[396])^(a[30] & b[397])^(a[29] & b[398])^(a[28] & b[399])^(a[27] & b[400])^(a[26] & b[401])^(a[25] & b[402])^(a[24] & b[403])^(a[23] & b[404])^(a[22] & b[405])^(a[21] & b[406])^(a[20] & b[407])^(a[19] & b[408]);
assign y[428] = (a[408] & b[20])^(a[407] & b[21])^(a[406] & b[22])^(a[405] & b[23])^(a[404] & b[24])^(a[403] & b[25])^(a[402] & b[26])^(a[401] & b[27])^(a[400] & b[28])^(a[399] & b[29])^(a[398] & b[30])^(a[397] & b[31])^(a[396] & b[32])^(a[395] & b[33])^(a[394] & b[34])^(a[393] & b[35])^(a[392] & b[36])^(a[391] & b[37])^(a[390] & b[38])^(a[389] & b[39])^(a[388] & b[40])^(a[387] & b[41])^(a[386] & b[42])^(a[385] & b[43])^(a[384] & b[44])^(a[383] & b[45])^(a[382] & b[46])^(a[381] & b[47])^(a[380] & b[48])^(a[379] & b[49])^(a[378] & b[50])^(a[377] & b[51])^(a[376] & b[52])^(a[375] & b[53])^(a[374] & b[54])^(a[373] & b[55])^(a[372] & b[56])^(a[371] & b[57])^(a[370] & b[58])^(a[369] & b[59])^(a[368] & b[60])^(a[367] & b[61])^(a[366] & b[62])^(a[365] & b[63])^(a[364] & b[64])^(a[363] & b[65])^(a[362] & b[66])^(a[361] & b[67])^(a[360] & b[68])^(a[359] & b[69])^(a[358] & b[70])^(a[357] & b[71])^(a[356] & b[72])^(a[355] & b[73])^(a[354] & b[74])^(a[353] & b[75])^(a[352] & b[76])^(a[351] & b[77])^(a[350] & b[78])^(a[349] & b[79])^(a[348] & b[80])^(a[347] & b[81])^(a[346] & b[82])^(a[345] & b[83])^(a[344] & b[84])^(a[343] & b[85])^(a[342] & b[86])^(a[341] & b[87])^(a[340] & b[88])^(a[339] & b[89])^(a[338] & b[90])^(a[337] & b[91])^(a[336] & b[92])^(a[335] & b[93])^(a[334] & b[94])^(a[333] & b[95])^(a[332] & b[96])^(a[331] & b[97])^(a[330] & b[98])^(a[329] & b[99])^(a[328] & b[100])^(a[327] & b[101])^(a[326] & b[102])^(a[325] & b[103])^(a[324] & b[104])^(a[323] & b[105])^(a[322] & b[106])^(a[321] & b[107])^(a[320] & b[108])^(a[319] & b[109])^(a[318] & b[110])^(a[317] & b[111])^(a[316] & b[112])^(a[315] & b[113])^(a[314] & b[114])^(a[313] & b[115])^(a[312] & b[116])^(a[311] & b[117])^(a[310] & b[118])^(a[309] & b[119])^(a[308] & b[120])^(a[307] & b[121])^(a[306] & b[122])^(a[305] & b[123])^(a[304] & b[124])^(a[303] & b[125])^(a[302] & b[126])^(a[301] & b[127])^(a[300] & b[128])^(a[299] & b[129])^(a[298] & b[130])^(a[297] & b[131])^(a[296] & b[132])^(a[295] & b[133])^(a[294] & b[134])^(a[293] & b[135])^(a[292] & b[136])^(a[291] & b[137])^(a[290] & b[138])^(a[289] & b[139])^(a[288] & b[140])^(a[287] & b[141])^(a[286] & b[142])^(a[285] & b[143])^(a[284] & b[144])^(a[283] & b[145])^(a[282] & b[146])^(a[281] & b[147])^(a[280] & b[148])^(a[279] & b[149])^(a[278] & b[150])^(a[277] & b[151])^(a[276] & b[152])^(a[275] & b[153])^(a[274] & b[154])^(a[273] & b[155])^(a[272] & b[156])^(a[271] & b[157])^(a[270] & b[158])^(a[269] & b[159])^(a[268] & b[160])^(a[267] & b[161])^(a[266] & b[162])^(a[265] & b[163])^(a[264] & b[164])^(a[263] & b[165])^(a[262] & b[166])^(a[261] & b[167])^(a[260] & b[168])^(a[259] & b[169])^(a[258] & b[170])^(a[257] & b[171])^(a[256] & b[172])^(a[255] & b[173])^(a[254] & b[174])^(a[253] & b[175])^(a[252] & b[176])^(a[251] & b[177])^(a[250] & b[178])^(a[249] & b[179])^(a[248] & b[180])^(a[247] & b[181])^(a[246] & b[182])^(a[245] & b[183])^(a[244] & b[184])^(a[243] & b[185])^(a[242] & b[186])^(a[241] & b[187])^(a[240] & b[188])^(a[239] & b[189])^(a[238] & b[190])^(a[237] & b[191])^(a[236] & b[192])^(a[235] & b[193])^(a[234] & b[194])^(a[233] & b[195])^(a[232] & b[196])^(a[231] & b[197])^(a[230] & b[198])^(a[229] & b[199])^(a[228] & b[200])^(a[227] & b[201])^(a[226] & b[202])^(a[225] & b[203])^(a[224] & b[204])^(a[223] & b[205])^(a[222] & b[206])^(a[221] & b[207])^(a[220] & b[208])^(a[219] & b[209])^(a[218] & b[210])^(a[217] & b[211])^(a[216] & b[212])^(a[215] & b[213])^(a[214] & b[214])^(a[213] & b[215])^(a[212] & b[216])^(a[211] & b[217])^(a[210] & b[218])^(a[209] & b[219])^(a[208] & b[220])^(a[207] & b[221])^(a[206] & b[222])^(a[205] & b[223])^(a[204] & b[224])^(a[203] & b[225])^(a[202] & b[226])^(a[201] & b[227])^(a[200] & b[228])^(a[199] & b[229])^(a[198] & b[230])^(a[197] & b[231])^(a[196] & b[232])^(a[195] & b[233])^(a[194] & b[234])^(a[193] & b[235])^(a[192] & b[236])^(a[191] & b[237])^(a[190] & b[238])^(a[189] & b[239])^(a[188] & b[240])^(a[187] & b[241])^(a[186] & b[242])^(a[185] & b[243])^(a[184] & b[244])^(a[183] & b[245])^(a[182] & b[246])^(a[181] & b[247])^(a[180] & b[248])^(a[179] & b[249])^(a[178] & b[250])^(a[177] & b[251])^(a[176] & b[252])^(a[175] & b[253])^(a[174] & b[254])^(a[173] & b[255])^(a[172] & b[256])^(a[171] & b[257])^(a[170] & b[258])^(a[169] & b[259])^(a[168] & b[260])^(a[167] & b[261])^(a[166] & b[262])^(a[165] & b[263])^(a[164] & b[264])^(a[163] & b[265])^(a[162] & b[266])^(a[161] & b[267])^(a[160] & b[268])^(a[159] & b[269])^(a[158] & b[270])^(a[157] & b[271])^(a[156] & b[272])^(a[155] & b[273])^(a[154] & b[274])^(a[153] & b[275])^(a[152] & b[276])^(a[151] & b[277])^(a[150] & b[278])^(a[149] & b[279])^(a[148] & b[280])^(a[147] & b[281])^(a[146] & b[282])^(a[145] & b[283])^(a[144] & b[284])^(a[143] & b[285])^(a[142] & b[286])^(a[141] & b[287])^(a[140] & b[288])^(a[139] & b[289])^(a[138] & b[290])^(a[137] & b[291])^(a[136] & b[292])^(a[135] & b[293])^(a[134] & b[294])^(a[133] & b[295])^(a[132] & b[296])^(a[131] & b[297])^(a[130] & b[298])^(a[129] & b[299])^(a[128] & b[300])^(a[127] & b[301])^(a[126] & b[302])^(a[125] & b[303])^(a[124] & b[304])^(a[123] & b[305])^(a[122] & b[306])^(a[121] & b[307])^(a[120] & b[308])^(a[119] & b[309])^(a[118] & b[310])^(a[117] & b[311])^(a[116] & b[312])^(a[115] & b[313])^(a[114] & b[314])^(a[113] & b[315])^(a[112] & b[316])^(a[111] & b[317])^(a[110] & b[318])^(a[109] & b[319])^(a[108] & b[320])^(a[107] & b[321])^(a[106] & b[322])^(a[105] & b[323])^(a[104] & b[324])^(a[103] & b[325])^(a[102] & b[326])^(a[101] & b[327])^(a[100] & b[328])^(a[99] & b[329])^(a[98] & b[330])^(a[97] & b[331])^(a[96] & b[332])^(a[95] & b[333])^(a[94] & b[334])^(a[93] & b[335])^(a[92] & b[336])^(a[91] & b[337])^(a[90] & b[338])^(a[89] & b[339])^(a[88] & b[340])^(a[87] & b[341])^(a[86] & b[342])^(a[85] & b[343])^(a[84] & b[344])^(a[83] & b[345])^(a[82] & b[346])^(a[81] & b[347])^(a[80] & b[348])^(a[79] & b[349])^(a[78] & b[350])^(a[77] & b[351])^(a[76] & b[352])^(a[75] & b[353])^(a[74] & b[354])^(a[73] & b[355])^(a[72] & b[356])^(a[71] & b[357])^(a[70] & b[358])^(a[69] & b[359])^(a[68] & b[360])^(a[67] & b[361])^(a[66] & b[362])^(a[65] & b[363])^(a[64] & b[364])^(a[63] & b[365])^(a[62] & b[366])^(a[61] & b[367])^(a[60] & b[368])^(a[59] & b[369])^(a[58] & b[370])^(a[57] & b[371])^(a[56] & b[372])^(a[55] & b[373])^(a[54] & b[374])^(a[53] & b[375])^(a[52] & b[376])^(a[51] & b[377])^(a[50] & b[378])^(a[49] & b[379])^(a[48] & b[380])^(a[47] & b[381])^(a[46] & b[382])^(a[45] & b[383])^(a[44] & b[384])^(a[43] & b[385])^(a[42] & b[386])^(a[41] & b[387])^(a[40] & b[388])^(a[39] & b[389])^(a[38] & b[390])^(a[37] & b[391])^(a[36] & b[392])^(a[35] & b[393])^(a[34] & b[394])^(a[33] & b[395])^(a[32] & b[396])^(a[31] & b[397])^(a[30] & b[398])^(a[29] & b[399])^(a[28] & b[400])^(a[27] & b[401])^(a[26] & b[402])^(a[25] & b[403])^(a[24] & b[404])^(a[23] & b[405])^(a[22] & b[406])^(a[21] & b[407])^(a[20] & b[408]);
assign y[429] = (a[408] & b[21])^(a[407] & b[22])^(a[406] & b[23])^(a[405] & b[24])^(a[404] & b[25])^(a[403] & b[26])^(a[402] & b[27])^(a[401] & b[28])^(a[400] & b[29])^(a[399] & b[30])^(a[398] & b[31])^(a[397] & b[32])^(a[396] & b[33])^(a[395] & b[34])^(a[394] & b[35])^(a[393] & b[36])^(a[392] & b[37])^(a[391] & b[38])^(a[390] & b[39])^(a[389] & b[40])^(a[388] & b[41])^(a[387] & b[42])^(a[386] & b[43])^(a[385] & b[44])^(a[384] & b[45])^(a[383] & b[46])^(a[382] & b[47])^(a[381] & b[48])^(a[380] & b[49])^(a[379] & b[50])^(a[378] & b[51])^(a[377] & b[52])^(a[376] & b[53])^(a[375] & b[54])^(a[374] & b[55])^(a[373] & b[56])^(a[372] & b[57])^(a[371] & b[58])^(a[370] & b[59])^(a[369] & b[60])^(a[368] & b[61])^(a[367] & b[62])^(a[366] & b[63])^(a[365] & b[64])^(a[364] & b[65])^(a[363] & b[66])^(a[362] & b[67])^(a[361] & b[68])^(a[360] & b[69])^(a[359] & b[70])^(a[358] & b[71])^(a[357] & b[72])^(a[356] & b[73])^(a[355] & b[74])^(a[354] & b[75])^(a[353] & b[76])^(a[352] & b[77])^(a[351] & b[78])^(a[350] & b[79])^(a[349] & b[80])^(a[348] & b[81])^(a[347] & b[82])^(a[346] & b[83])^(a[345] & b[84])^(a[344] & b[85])^(a[343] & b[86])^(a[342] & b[87])^(a[341] & b[88])^(a[340] & b[89])^(a[339] & b[90])^(a[338] & b[91])^(a[337] & b[92])^(a[336] & b[93])^(a[335] & b[94])^(a[334] & b[95])^(a[333] & b[96])^(a[332] & b[97])^(a[331] & b[98])^(a[330] & b[99])^(a[329] & b[100])^(a[328] & b[101])^(a[327] & b[102])^(a[326] & b[103])^(a[325] & b[104])^(a[324] & b[105])^(a[323] & b[106])^(a[322] & b[107])^(a[321] & b[108])^(a[320] & b[109])^(a[319] & b[110])^(a[318] & b[111])^(a[317] & b[112])^(a[316] & b[113])^(a[315] & b[114])^(a[314] & b[115])^(a[313] & b[116])^(a[312] & b[117])^(a[311] & b[118])^(a[310] & b[119])^(a[309] & b[120])^(a[308] & b[121])^(a[307] & b[122])^(a[306] & b[123])^(a[305] & b[124])^(a[304] & b[125])^(a[303] & b[126])^(a[302] & b[127])^(a[301] & b[128])^(a[300] & b[129])^(a[299] & b[130])^(a[298] & b[131])^(a[297] & b[132])^(a[296] & b[133])^(a[295] & b[134])^(a[294] & b[135])^(a[293] & b[136])^(a[292] & b[137])^(a[291] & b[138])^(a[290] & b[139])^(a[289] & b[140])^(a[288] & b[141])^(a[287] & b[142])^(a[286] & b[143])^(a[285] & b[144])^(a[284] & b[145])^(a[283] & b[146])^(a[282] & b[147])^(a[281] & b[148])^(a[280] & b[149])^(a[279] & b[150])^(a[278] & b[151])^(a[277] & b[152])^(a[276] & b[153])^(a[275] & b[154])^(a[274] & b[155])^(a[273] & b[156])^(a[272] & b[157])^(a[271] & b[158])^(a[270] & b[159])^(a[269] & b[160])^(a[268] & b[161])^(a[267] & b[162])^(a[266] & b[163])^(a[265] & b[164])^(a[264] & b[165])^(a[263] & b[166])^(a[262] & b[167])^(a[261] & b[168])^(a[260] & b[169])^(a[259] & b[170])^(a[258] & b[171])^(a[257] & b[172])^(a[256] & b[173])^(a[255] & b[174])^(a[254] & b[175])^(a[253] & b[176])^(a[252] & b[177])^(a[251] & b[178])^(a[250] & b[179])^(a[249] & b[180])^(a[248] & b[181])^(a[247] & b[182])^(a[246] & b[183])^(a[245] & b[184])^(a[244] & b[185])^(a[243] & b[186])^(a[242] & b[187])^(a[241] & b[188])^(a[240] & b[189])^(a[239] & b[190])^(a[238] & b[191])^(a[237] & b[192])^(a[236] & b[193])^(a[235] & b[194])^(a[234] & b[195])^(a[233] & b[196])^(a[232] & b[197])^(a[231] & b[198])^(a[230] & b[199])^(a[229] & b[200])^(a[228] & b[201])^(a[227] & b[202])^(a[226] & b[203])^(a[225] & b[204])^(a[224] & b[205])^(a[223] & b[206])^(a[222] & b[207])^(a[221] & b[208])^(a[220] & b[209])^(a[219] & b[210])^(a[218] & b[211])^(a[217] & b[212])^(a[216] & b[213])^(a[215] & b[214])^(a[214] & b[215])^(a[213] & b[216])^(a[212] & b[217])^(a[211] & b[218])^(a[210] & b[219])^(a[209] & b[220])^(a[208] & b[221])^(a[207] & b[222])^(a[206] & b[223])^(a[205] & b[224])^(a[204] & b[225])^(a[203] & b[226])^(a[202] & b[227])^(a[201] & b[228])^(a[200] & b[229])^(a[199] & b[230])^(a[198] & b[231])^(a[197] & b[232])^(a[196] & b[233])^(a[195] & b[234])^(a[194] & b[235])^(a[193] & b[236])^(a[192] & b[237])^(a[191] & b[238])^(a[190] & b[239])^(a[189] & b[240])^(a[188] & b[241])^(a[187] & b[242])^(a[186] & b[243])^(a[185] & b[244])^(a[184] & b[245])^(a[183] & b[246])^(a[182] & b[247])^(a[181] & b[248])^(a[180] & b[249])^(a[179] & b[250])^(a[178] & b[251])^(a[177] & b[252])^(a[176] & b[253])^(a[175] & b[254])^(a[174] & b[255])^(a[173] & b[256])^(a[172] & b[257])^(a[171] & b[258])^(a[170] & b[259])^(a[169] & b[260])^(a[168] & b[261])^(a[167] & b[262])^(a[166] & b[263])^(a[165] & b[264])^(a[164] & b[265])^(a[163] & b[266])^(a[162] & b[267])^(a[161] & b[268])^(a[160] & b[269])^(a[159] & b[270])^(a[158] & b[271])^(a[157] & b[272])^(a[156] & b[273])^(a[155] & b[274])^(a[154] & b[275])^(a[153] & b[276])^(a[152] & b[277])^(a[151] & b[278])^(a[150] & b[279])^(a[149] & b[280])^(a[148] & b[281])^(a[147] & b[282])^(a[146] & b[283])^(a[145] & b[284])^(a[144] & b[285])^(a[143] & b[286])^(a[142] & b[287])^(a[141] & b[288])^(a[140] & b[289])^(a[139] & b[290])^(a[138] & b[291])^(a[137] & b[292])^(a[136] & b[293])^(a[135] & b[294])^(a[134] & b[295])^(a[133] & b[296])^(a[132] & b[297])^(a[131] & b[298])^(a[130] & b[299])^(a[129] & b[300])^(a[128] & b[301])^(a[127] & b[302])^(a[126] & b[303])^(a[125] & b[304])^(a[124] & b[305])^(a[123] & b[306])^(a[122] & b[307])^(a[121] & b[308])^(a[120] & b[309])^(a[119] & b[310])^(a[118] & b[311])^(a[117] & b[312])^(a[116] & b[313])^(a[115] & b[314])^(a[114] & b[315])^(a[113] & b[316])^(a[112] & b[317])^(a[111] & b[318])^(a[110] & b[319])^(a[109] & b[320])^(a[108] & b[321])^(a[107] & b[322])^(a[106] & b[323])^(a[105] & b[324])^(a[104] & b[325])^(a[103] & b[326])^(a[102] & b[327])^(a[101] & b[328])^(a[100] & b[329])^(a[99] & b[330])^(a[98] & b[331])^(a[97] & b[332])^(a[96] & b[333])^(a[95] & b[334])^(a[94] & b[335])^(a[93] & b[336])^(a[92] & b[337])^(a[91] & b[338])^(a[90] & b[339])^(a[89] & b[340])^(a[88] & b[341])^(a[87] & b[342])^(a[86] & b[343])^(a[85] & b[344])^(a[84] & b[345])^(a[83] & b[346])^(a[82] & b[347])^(a[81] & b[348])^(a[80] & b[349])^(a[79] & b[350])^(a[78] & b[351])^(a[77] & b[352])^(a[76] & b[353])^(a[75] & b[354])^(a[74] & b[355])^(a[73] & b[356])^(a[72] & b[357])^(a[71] & b[358])^(a[70] & b[359])^(a[69] & b[360])^(a[68] & b[361])^(a[67] & b[362])^(a[66] & b[363])^(a[65] & b[364])^(a[64] & b[365])^(a[63] & b[366])^(a[62] & b[367])^(a[61] & b[368])^(a[60] & b[369])^(a[59] & b[370])^(a[58] & b[371])^(a[57] & b[372])^(a[56] & b[373])^(a[55] & b[374])^(a[54] & b[375])^(a[53] & b[376])^(a[52] & b[377])^(a[51] & b[378])^(a[50] & b[379])^(a[49] & b[380])^(a[48] & b[381])^(a[47] & b[382])^(a[46] & b[383])^(a[45] & b[384])^(a[44] & b[385])^(a[43] & b[386])^(a[42] & b[387])^(a[41] & b[388])^(a[40] & b[389])^(a[39] & b[390])^(a[38] & b[391])^(a[37] & b[392])^(a[36] & b[393])^(a[35] & b[394])^(a[34] & b[395])^(a[33] & b[396])^(a[32] & b[397])^(a[31] & b[398])^(a[30] & b[399])^(a[29] & b[400])^(a[28] & b[401])^(a[27] & b[402])^(a[26] & b[403])^(a[25] & b[404])^(a[24] & b[405])^(a[23] & b[406])^(a[22] & b[407])^(a[21] & b[408]);
assign y[430] = (a[408] & b[22])^(a[407] & b[23])^(a[406] & b[24])^(a[405] & b[25])^(a[404] & b[26])^(a[403] & b[27])^(a[402] & b[28])^(a[401] & b[29])^(a[400] & b[30])^(a[399] & b[31])^(a[398] & b[32])^(a[397] & b[33])^(a[396] & b[34])^(a[395] & b[35])^(a[394] & b[36])^(a[393] & b[37])^(a[392] & b[38])^(a[391] & b[39])^(a[390] & b[40])^(a[389] & b[41])^(a[388] & b[42])^(a[387] & b[43])^(a[386] & b[44])^(a[385] & b[45])^(a[384] & b[46])^(a[383] & b[47])^(a[382] & b[48])^(a[381] & b[49])^(a[380] & b[50])^(a[379] & b[51])^(a[378] & b[52])^(a[377] & b[53])^(a[376] & b[54])^(a[375] & b[55])^(a[374] & b[56])^(a[373] & b[57])^(a[372] & b[58])^(a[371] & b[59])^(a[370] & b[60])^(a[369] & b[61])^(a[368] & b[62])^(a[367] & b[63])^(a[366] & b[64])^(a[365] & b[65])^(a[364] & b[66])^(a[363] & b[67])^(a[362] & b[68])^(a[361] & b[69])^(a[360] & b[70])^(a[359] & b[71])^(a[358] & b[72])^(a[357] & b[73])^(a[356] & b[74])^(a[355] & b[75])^(a[354] & b[76])^(a[353] & b[77])^(a[352] & b[78])^(a[351] & b[79])^(a[350] & b[80])^(a[349] & b[81])^(a[348] & b[82])^(a[347] & b[83])^(a[346] & b[84])^(a[345] & b[85])^(a[344] & b[86])^(a[343] & b[87])^(a[342] & b[88])^(a[341] & b[89])^(a[340] & b[90])^(a[339] & b[91])^(a[338] & b[92])^(a[337] & b[93])^(a[336] & b[94])^(a[335] & b[95])^(a[334] & b[96])^(a[333] & b[97])^(a[332] & b[98])^(a[331] & b[99])^(a[330] & b[100])^(a[329] & b[101])^(a[328] & b[102])^(a[327] & b[103])^(a[326] & b[104])^(a[325] & b[105])^(a[324] & b[106])^(a[323] & b[107])^(a[322] & b[108])^(a[321] & b[109])^(a[320] & b[110])^(a[319] & b[111])^(a[318] & b[112])^(a[317] & b[113])^(a[316] & b[114])^(a[315] & b[115])^(a[314] & b[116])^(a[313] & b[117])^(a[312] & b[118])^(a[311] & b[119])^(a[310] & b[120])^(a[309] & b[121])^(a[308] & b[122])^(a[307] & b[123])^(a[306] & b[124])^(a[305] & b[125])^(a[304] & b[126])^(a[303] & b[127])^(a[302] & b[128])^(a[301] & b[129])^(a[300] & b[130])^(a[299] & b[131])^(a[298] & b[132])^(a[297] & b[133])^(a[296] & b[134])^(a[295] & b[135])^(a[294] & b[136])^(a[293] & b[137])^(a[292] & b[138])^(a[291] & b[139])^(a[290] & b[140])^(a[289] & b[141])^(a[288] & b[142])^(a[287] & b[143])^(a[286] & b[144])^(a[285] & b[145])^(a[284] & b[146])^(a[283] & b[147])^(a[282] & b[148])^(a[281] & b[149])^(a[280] & b[150])^(a[279] & b[151])^(a[278] & b[152])^(a[277] & b[153])^(a[276] & b[154])^(a[275] & b[155])^(a[274] & b[156])^(a[273] & b[157])^(a[272] & b[158])^(a[271] & b[159])^(a[270] & b[160])^(a[269] & b[161])^(a[268] & b[162])^(a[267] & b[163])^(a[266] & b[164])^(a[265] & b[165])^(a[264] & b[166])^(a[263] & b[167])^(a[262] & b[168])^(a[261] & b[169])^(a[260] & b[170])^(a[259] & b[171])^(a[258] & b[172])^(a[257] & b[173])^(a[256] & b[174])^(a[255] & b[175])^(a[254] & b[176])^(a[253] & b[177])^(a[252] & b[178])^(a[251] & b[179])^(a[250] & b[180])^(a[249] & b[181])^(a[248] & b[182])^(a[247] & b[183])^(a[246] & b[184])^(a[245] & b[185])^(a[244] & b[186])^(a[243] & b[187])^(a[242] & b[188])^(a[241] & b[189])^(a[240] & b[190])^(a[239] & b[191])^(a[238] & b[192])^(a[237] & b[193])^(a[236] & b[194])^(a[235] & b[195])^(a[234] & b[196])^(a[233] & b[197])^(a[232] & b[198])^(a[231] & b[199])^(a[230] & b[200])^(a[229] & b[201])^(a[228] & b[202])^(a[227] & b[203])^(a[226] & b[204])^(a[225] & b[205])^(a[224] & b[206])^(a[223] & b[207])^(a[222] & b[208])^(a[221] & b[209])^(a[220] & b[210])^(a[219] & b[211])^(a[218] & b[212])^(a[217] & b[213])^(a[216] & b[214])^(a[215] & b[215])^(a[214] & b[216])^(a[213] & b[217])^(a[212] & b[218])^(a[211] & b[219])^(a[210] & b[220])^(a[209] & b[221])^(a[208] & b[222])^(a[207] & b[223])^(a[206] & b[224])^(a[205] & b[225])^(a[204] & b[226])^(a[203] & b[227])^(a[202] & b[228])^(a[201] & b[229])^(a[200] & b[230])^(a[199] & b[231])^(a[198] & b[232])^(a[197] & b[233])^(a[196] & b[234])^(a[195] & b[235])^(a[194] & b[236])^(a[193] & b[237])^(a[192] & b[238])^(a[191] & b[239])^(a[190] & b[240])^(a[189] & b[241])^(a[188] & b[242])^(a[187] & b[243])^(a[186] & b[244])^(a[185] & b[245])^(a[184] & b[246])^(a[183] & b[247])^(a[182] & b[248])^(a[181] & b[249])^(a[180] & b[250])^(a[179] & b[251])^(a[178] & b[252])^(a[177] & b[253])^(a[176] & b[254])^(a[175] & b[255])^(a[174] & b[256])^(a[173] & b[257])^(a[172] & b[258])^(a[171] & b[259])^(a[170] & b[260])^(a[169] & b[261])^(a[168] & b[262])^(a[167] & b[263])^(a[166] & b[264])^(a[165] & b[265])^(a[164] & b[266])^(a[163] & b[267])^(a[162] & b[268])^(a[161] & b[269])^(a[160] & b[270])^(a[159] & b[271])^(a[158] & b[272])^(a[157] & b[273])^(a[156] & b[274])^(a[155] & b[275])^(a[154] & b[276])^(a[153] & b[277])^(a[152] & b[278])^(a[151] & b[279])^(a[150] & b[280])^(a[149] & b[281])^(a[148] & b[282])^(a[147] & b[283])^(a[146] & b[284])^(a[145] & b[285])^(a[144] & b[286])^(a[143] & b[287])^(a[142] & b[288])^(a[141] & b[289])^(a[140] & b[290])^(a[139] & b[291])^(a[138] & b[292])^(a[137] & b[293])^(a[136] & b[294])^(a[135] & b[295])^(a[134] & b[296])^(a[133] & b[297])^(a[132] & b[298])^(a[131] & b[299])^(a[130] & b[300])^(a[129] & b[301])^(a[128] & b[302])^(a[127] & b[303])^(a[126] & b[304])^(a[125] & b[305])^(a[124] & b[306])^(a[123] & b[307])^(a[122] & b[308])^(a[121] & b[309])^(a[120] & b[310])^(a[119] & b[311])^(a[118] & b[312])^(a[117] & b[313])^(a[116] & b[314])^(a[115] & b[315])^(a[114] & b[316])^(a[113] & b[317])^(a[112] & b[318])^(a[111] & b[319])^(a[110] & b[320])^(a[109] & b[321])^(a[108] & b[322])^(a[107] & b[323])^(a[106] & b[324])^(a[105] & b[325])^(a[104] & b[326])^(a[103] & b[327])^(a[102] & b[328])^(a[101] & b[329])^(a[100] & b[330])^(a[99] & b[331])^(a[98] & b[332])^(a[97] & b[333])^(a[96] & b[334])^(a[95] & b[335])^(a[94] & b[336])^(a[93] & b[337])^(a[92] & b[338])^(a[91] & b[339])^(a[90] & b[340])^(a[89] & b[341])^(a[88] & b[342])^(a[87] & b[343])^(a[86] & b[344])^(a[85] & b[345])^(a[84] & b[346])^(a[83] & b[347])^(a[82] & b[348])^(a[81] & b[349])^(a[80] & b[350])^(a[79] & b[351])^(a[78] & b[352])^(a[77] & b[353])^(a[76] & b[354])^(a[75] & b[355])^(a[74] & b[356])^(a[73] & b[357])^(a[72] & b[358])^(a[71] & b[359])^(a[70] & b[360])^(a[69] & b[361])^(a[68] & b[362])^(a[67] & b[363])^(a[66] & b[364])^(a[65] & b[365])^(a[64] & b[366])^(a[63] & b[367])^(a[62] & b[368])^(a[61] & b[369])^(a[60] & b[370])^(a[59] & b[371])^(a[58] & b[372])^(a[57] & b[373])^(a[56] & b[374])^(a[55] & b[375])^(a[54] & b[376])^(a[53] & b[377])^(a[52] & b[378])^(a[51] & b[379])^(a[50] & b[380])^(a[49] & b[381])^(a[48] & b[382])^(a[47] & b[383])^(a[46] & b[384])^(a[45] & b[385])^(a[44] & b[386])^(a[43] & b[387])^(a[42] & b[388])^(a[41] & b[389])^(a[40] & b[390])^(a[39] & b[391])^(a[38] & b[392])^(a[37] & b[393])^(a[36] & b[394])^(a[35] & b[395])^(a[34] & b[396])^(a[33] & b[397])^(a[32] & b[398])^(a[31] & b[399])^(a[30] & b[400])^(a[29] & b[401])^(a[28] & b[402])^(a[27] & b[403])^(a[26] & b[404])^(a[25] & b[405])^(a[24] & b[406])^(a[23] & b[407])^(a[22] & b[408]);
assign y[431] = (a[408] & b[23])^(a[407] & b[24])^(a[406] & b[25])^(a[405] & b[26])^(a[404] & b[27])^(a[403] & b[28])^(a[402] & b[29])^(a[401] & b[30])^(a[400] & b[31])^(a[399] & b[32])^(a[398] & b[33])^(a[397] & b[34])^(a[396] & b[35])^(a[395] & b[36])^(a[394] & b[37])^(a[393] & b[38])^(a[392] & b[39])^(a[391] & b[40])^(a[390] & b[41])^(a[389] & b[42])^(a[388] & b[43])^(a[387] & b[44])^(a[386] & b[45])^(a[385] & b[46])^(a[384] & b[47])^(a[383] & b[48])^(a[382] & b[49])^(a[381] & b[50])^(a[380] & b[51])^(a[379] & b[52])^(a[378] & b[53])^(a[377] & b[54])^(a[376] & b[55])^(a[375] & b[56])^(a[374] & b[57])^(a[373] & b[58])^(a[372] & b[59])^(a[371] & b[60])^(a[370] & b[61])^(a[369] & b[62])^(a[368] & b[63])^(a[367] & b[64])^(a[366] & b[65])^(a[365] & b[66])^(a[364] & b[67])^(a[363] & b[68])^(a[362] & b[69])^(a[361] & b[70])^(a[360] & b[71])^(a[359] & b[72])^(a[358] & b[73])^(a[357] & b[74])^(a[356] & b[75])^(a[355] & b[76])^(a[354] & b[77])^(a[353] & b[78])^(a[352] & b[79])^(a[351] & b[80])^(a[350] & b[81])^(a[349] & b[82])^(a[348] & b[83])^(a[347] & b[84])^(a[346] & b[85])^(a[345] & b[86])^(a[344] & b[87])^(a[343] & b[88])^(a[342] & b[89])^(a[341] & b[90])^(a[340] & b[91])^(a[339] & b[92])^(a[338] & b[93])^(a[337] & b[94])^(a[336] & b[95])^(a[335] & b[96])^(a[334] & b[97])^(a[333] & b[98])^(a[332] & b[99])^(a[331] & b[100])^(a[330] & b[101])^(a[329] & b[102])^(a[328] & b[103])^(a[327] & b[104])^(a[326] & b[105])^(a[325] & b[106])^(a[324] & b[107])^(a[323] & b[108])^(a[322] & b[109])^(a[321] & b[110])^(a[320] & b[111])^(a[319] & b[112])^(a[318] & b[113])^(a[317] & b[114])^(a[316] & b[115])^(a[315] & b[116])^(a[314] & b[117])^(a[313] & b[118])^(a[312] & b[119])^(a[311] & b[120])^(a[310] & b[121])^(a[309] & b[122])^(a[308] & b[123])^(a[307] & b[124])^(a[306] & b[125])^(a[305] & b[126])^(a[304] & b[127])^(a[303] & b[128])^(a[302] & b[129])^(a[301] & b[130])^(a[300] & b[131])^(a[299] & b[132])^(a[298] & b[133])^(a[297] & b[134])^(a[296] & b[135])^(a[295] & b[136])^(a[294] & b[137])^(a[293] & b[138])^(a[292] & b[139])^(a[291] & b[140])^(a[290] & b[141])^(a[289] & b[142])^(a[288] & b[143])^(a[287] & b[144])^(a[286] & b[145])^(a[285] & b[146])^(a[284] & b[147])^(a[283] & b[148])^(a[282] & b[149])^(a[281] & b[150])^(a[280] & b[151])^(a[279] & b[152])^(a[278] & b[153])^(a[277] & b[154])^(a[276] & b[155])^(a[275] & b[156])^(a[274] & b[157])^(a[273] & b[158])^(a[272] & b[159])^(a[271] & b[160])^(a[270] & b[161])^(a[269] & b[162])^(a[268] & b[163])^(a[267] & b[164])^(a[266] & b[165])^(a[265] & b[166])^(a[264] & b[167])^(a[263] & b[168])^(a[262] & b[169])^(a[261] & b[170])^(a[260] & b[171])^(a[259] & b[172])^(a[258] & b[173])^(a[257] & b[174])^(a[256] & b[175])^(a[255] & b[176])^(a[254] & b[177])^(a[253] & b[178])^(a[252] & b[179])^(a[251] & b[180])^(a[250] & b[181])^(a[249] & b[182])^(a[248] & b[183])^(a[247] & b[184])^(a[246] & b[185])^(a[245] & b[186])^(a[244] & b[187])^(a[243] & b[188])^(a[242] & b[189])^(a[241] & b[190])^(a[240] & b[191])^(a[239] & b[192])^(a[238] & b[193])^(a[237] & b[194])^(a[236] & b[195])^(a[235] & b[196])^(a[234] & b[197])^(a[233] & b[198])^(a[232] & b[199])^(a[231] & b[200])^(a[230] & b[201])^(a[229] & b[202])^(a[228] & b[203])^(a[227] & b[204])^(a[226] & b[205])^(a[225] & b[206])^(a[224] & b[207])^(a[223] & b[208])^(a[222] & b[209])^(a[221] & b[210])^(a[220] & b[211])^(a[219] & b[212])^(a[218] & b[213])^(a[217] & b[214])^(a[216] & b[215])^(a[215] & b[216])^(a[214] & b[217])^(a[213] & b[218])^(a[212] & b[219])^(a[211] & b[220])^(a[210] & b[221])^(a[209] & b[222])^(a[208] & b[223])^(a[207] & b[224])^(a[206] & b[225])^(a[205] & b[226])^(a[204] & b[227])^(a[203] & b[228])^(a[202] & b[229])^(a[201] & b[230])^(a[200] & b[231])^(a[199] & b[232])^(a[198] & b[233])^(a[197] & b[234])^(a[196] & b[235])^(a[195] & b[236])^(a[194] & b[237])^(a[193] & b[238])^(a[192] & b[239])^(a[191] & b[240])^(a[190] & b[241])^(a[189] & b[242])^(a[188] & b[243])^(a[187] & b[244])^(a[186] & b[245])^(a[185] & b[246])^(a[184] & b[247])^(a[183] & b[248])^(a[182] & b[249])^(a[181] & b[250])^(a[180] & b[251])^(a[179] & b[252])^(a[178] & b[253])^(a[177] & b[254])^(a[176] & b[255])^(a[175] & b[256])^(a[174] & b[257])^(a[173] & b[258])^(a[172] & b[259])^(a[171] & b[260])^(a[170] & b[261])^(a[169] & b[262])^(a[168] & b[263])^(a[167] & b[264])^(a[166] & b[265])^(a[165] & b[266])^(a[164] & b[267])^(a[163] & b[268])^(a[162] & b[269])^(a[161] & b[270])^(a[160] & b[271])^(a[159] & b[272])^(a[158] & b[273])^(a[157] & b[274])^(a[156] & b[275])^(a[155] & b[276])^(a[154] & b[277])^(a[153] & b[278])^(a[152] & b[279])^(a[151] & b[280])^(a[150] & b[281])^(a[149] & b[282])^(a[148] & b[283])^(a[147] & b[284])^(a[146] & b[285])^(a[145] & b[286])^(a[144] & b[287])^(a[143] & b[288])^(a[142] & b[289])^(a[141] & b[290])^(a[140] & b[291])^(a[139] & b[292])^(a[138] & b[293])^(a[137] & b[294])^(a[136] & b[295])^(a[135] & b[296])^(a[134] & b[297])^(a[133] & b[298])^(a[132] & b[299])^(a[131] & b[300])^(a[130] & b[301])^(a[129] & b[302])^(a[128] & b[303])^(a[127] & b[304])^(a[126] & b[305])^(a[125] & b[306])^(a[124] & b[307])^(a[123] & b[308])^(a[122] & b[309])^(a[121] & b[310])^(a[120] & b[311])^(a[119] & b[312])^(a[118] & b[313])^(a[117] & b[314])^(a[116] & b[315])^(a[115] & b[316])^(a[114] & b[317])^(a[113] & b[318])^(a[112] & b[319])^(a[111] & b[320])^(a[110] & b[321])^(a[109] & b[322])^(a[108] & b[323])^(a[107] & b[324])^(a[106] & b[325])^(a[105] & b[326])^(a[104] & b[327])^(a[103] & b[328])^(a[102] & b[329])^(a[101] & b[330])^(a[100] & b[331])^(a[99] & b[332])^(a[98] & b[333])^(a[97] & b[334])^(a[96] & b[335])^(a[95] & b[336])^(a[94] & b[337])^(a[93] & b[338])^(a[92] & b[339])^(a[91] & b[340])^(a[90] & b[341])^(a[89] & b[342])^(a[88] & b[343])^(a[87] & b[344])^(a[86] & b[345])^(a[85] & b[346])^(a[84] & b[347])^(a[83] & b[348])^(a[82] & b[349])^(a[81] & b[350])^(a[80] & b[351])^(a[79] & b[352])^(a[78] & b[353])^(a[77] & b[354])^(a[76] & b[355])^(a[75] & b[356])^(a[74] & b[357])^(a[73] & b[358])^(a[72] & b[359])^(a[71] & b[360])^(a[70] & b[361])^(a[69] & b[362])^(a[68] & b[363])^(a[67] & b[364])^(a[66] & b[365])^(a[65] & b[366])^(a[64] & b[367])^(a[63] & b[368])^(a[62] & b[369])^(a[61] & b[370])^(a[60] & b[371])^(a[59] & b[372])^(a[58] & b[373])^(a[57] & b[374])^(a[56] & b[375])^(a[55] & b[376])^(a[54] & b[377])^(a[53] & b[378])^(a[52] & b[379])^(a[51] & b[380])^(a[50] & b[381])^(a[49] & b[382])^(a[48] & b[383])^(a[47] & b[384])^(a[46] & b[385])^(a[45] & b[386])^(a[44] & b[387])^(a[43] & b[388])^(a[42] & b[389])^(a[41] & b[390])^(a[40] & b[391])^(a[39] & b[392])^(a[38] & b[393])^(a[37] & b[394])^(a[36] & b[395])^(a[35] & b[396])^(a[34] & b[397])^(a[33] & b[398])^(a[32] & b[399])^(a[31] & b[400])^(a[30] & b[401])^(a[29] & b[402])^(a[28] & b[403])^(a[27] & b[404])^(a[26] & b[405])^(a[25] & b[406])^(a[24] & b[407])^(a[23] & b[408]);
assign y[432] = (a[408] & b[24])^(a[407] & b[25])^(a[406] & b[26])^(a[405] & b[27])^(a[404] & b[28])^(a[403] & b[29])^(a[402] & b[30])^(a[401] & b[31])^(a[400] & b[32])^(a[399] & b[33])^(a[398] & b[34])^(a[397] & b[35])^(a[396] & b[36])^(a[395] & b[37])^(a[394] & b[38])^(a[393] & b[39])^(a[392] & b[40])^(a[391] & b[41])^(a[390] & b[42])^(a[389] & b[43])^(a[388] & b[44])^(a[387] & b[45])^(a[386] & b[46])^(a[385] & b[47])^(a[384] & b[48])^(a[383] & b[49])^(a[382] & b[50])^(a[381] & b[51])^(a[380] & b[52])^(a[379] & b[53])^(a[378] & b[54])^(a[377] & b[55])^(a[376] & b[56])^(a[375] & b[57])^(a[374] & b[58])^(a[373] & b[59])^(a[372] & b[60])^(a[371] & b[61])^(a[370] & b[62])^(a[369] & b[63])^(a[368] & b[64])^(a[367] & b[65])^(a[366] & b[66])^(a[365] & b[67])^(a[364] & b[68])^(a[363] & b[69])^(a[362] & b[70])^(a[361] & b[71])^(a[360] & b[72])^(a[359] & b[73])^(a[358] & b[74])^(a[357] & b[75])^(a[356] & b[76])^(a[355] & b[77])^(a[354] & b[78])^(a[353] & b[79])^(a[352] & b[80])^(a[351] & b[81])^(a[350] & b[82])^(a[349] & b[83])^(a[348] & b[84])^(a[347] & b[85])^(a[346] & b[86])^(a[345] & b[87])^(a[344] & b[88])^(a[343] & b[89])^(a[342] & b[90])^(a[341] & b[91])^(a[340] & b[92])^(a[339] & b[93])^(a[338] & b[94])^(a[337] & b[95])^(a[336] & b[96])^(a[335] & b[97])^(a[334] & b[98])^(a[333] & b[99])^(a[332] & b[100])^(a[331] & b[101])^(a[330] & b[102])^(a[329] & b[103])^(a[328] & b[104])^(a[327] & b[105])^(a[326] & b[106])^(a[325] & b[107])^(a[324] & b[108])^(a[323] & b[109])^(a[322] & b[110])^(a[321] & b[111])^(a[320] & b[112])^(a[319] & b[113])^(a[318] & b[114])^(a[317] & b[115])^(a[316] & b[116])^(a[315] & b[117])^(a[314] & b[118])^(a[313] & b[119])^(a[312] & b[120])^(a[311] & b[121])^(a[310] & b[122])^(a[309] & b[123])^(a[308] & b[124])^(a[307] & b[125])^(a[306] & b[126])^(a[305] & b[127])^(a[304] & b[128])^(a[303] & b[129])^(a[302] & b[130])^(a[301] & b[131])^(a[300] & b[132])^(a[299] & b[133])^(a[298] & b[134])^(a[297] & b[135])^(a[296] & b[136])^(a[295] & b[137])^(a[294] & b[138])^(a[293] & b[139])^(a[292] & b[140])^(a[291] & b[141])^(a[290] & b[142])^(a[289] & b[143])^(a[288] & b[144])^(a[287] & b[145])^(a[286] & b[146])^(a[285] & b[147])^(a[284] & b[148])^(a[283] & b[149])^(a[282] & b[150])^(a[281] & b[151])^(a[280] & b[152])^(a[279] & b[153])^(a[278] & b[154])^(a[277] & b[155])^(a[276] & b[156])^(a[275] & b[157])^(a[274] & b[158])^(a[273] & b[159])^(a[272] & b[160])^(a[271] & b[161])^(a[270] & b[162])^(a[269] & b[163])^(a[268] & b[164])^(a[267] & b[165])^(a[266] & b[166])^(a[265] & b[167])^(a[264] & b[168])^(a[263] & b[169])^(a[262] & b[170])^(a[261] & b[171])^(a[260] & b[172])^(a[259] & b[173])^(a[258] & b[174])^(a[257] & b[175])^(a[256] & b[176])^(a[255] & b[177])^(a[254] & b[178])^(a[253] & b[179])^(a[252] & b[180])^(a[251] & b[181])^(a[250] & b[182])^(a[249] & b[183])^(a[248] & b[184])^(a[247] & b[185])^(a[246] & b[186])^(a[245] & b[187])^(a[244] & b[188])^(a[243] & b[189])^(a[242] & b[190])^(a[241] & b[191])^(a[240] & b[192])^(a[239] & b[193])^(a[238] & b[194])^(a[237] & b[195])^(a[236] & b[196])^(a[235] & b[197])^(a[234] & b[198])^(a[233] & b[199])^(a[232] & b[200])^(a[231] & b[201])^(a[230] & b[202])^(a[229] & b[203])^(a[228] & b[204])^(a[227] & b[205])^(a[226] & b[206])^(a[225] & b[207])^(a[224] & b[208])^(a[223] & b[209])^(a[222] & b[210])^(a[221] & b[211])^(a[220] & b[212])^(a[219] & b[213])^(a[218] & b[214])^(a[217] & b[215])^(a[216] & b[216])^(a[215] & b[217])^(a[214] & b[218])^(a[213] & b[219])^(a[212] & b[220])^(a[211] & b[221])^(a[210] & b[222])^(a[209] & b[223])^(a[208] & b[224])^(a[207] & b[225])^(a[206] & b[226])^(a[205] & b[227])^(a[204] & b[228])^(a[203] & b[229])^(a[202] & b[230])^(a[201] & b[231])^(a[200] & b[232])^(a[199] & b[233])^(a[198] & b[234])^(a[197] & b[235])^(a[196] & b[236])^(a[195] & b[237])^(a[194] & b[238])^(a[193] & b[239])^(a[192] & b[240])^(a[191] & b[241])^(a[190] & b[242])^(a[189] & b[243])^(a[188] & b[244])^(a[187] & b[245])^(a[186] & b[246])^(a[185] & b[247])^(a[184] & b[248])^(a[183] & b[249])^(a[182] & b[250])^(a[181] & b[251])^(a[180] & b[252])^(a[179] & b[253])^(a[178] & b[254])^(a[177] & b[255])^(a[176] & b[256])^(a[175] & b[257])^(a[174] & b[258])^(a[173] & b[259])^(a[172] & b[260])^(a[171] & b[261])^(a[170] & b[262])^(a[169] & b[263])^(a[168] & b[264])^(a[167] & b[265])^(a[166] & b[266])^(a[165] & b[267])^(a[164] & b[268])^(a[163] & b[269])^(a[162] & b[270])^(a[161] & b[271])^(a[160] & b[272])^(a[159] & b[273])^(a[158] & b[274])^(a[157] & b[275])^(a[156] & b[276])^(a[155] & b[277])^(a[154] & b[278])^(a[153] & b[279])^(a[152] & b[280])^(a[151] & b[281])^(a[150] & b[282])^(a[149] & b[283])^(a[148] & b[284])^(a[147] & b[285])^(a[146] & b[286])^(a[145] & b[287])^(a[144] & b[288])^(a[143] & b[289])^(a[142] & b[290])^(a[141] & b[291])^(a[140] & b[292])^(a[139] & b[293])^(a[138] & b[294])^(a[137] & b[295])^(a[136] & b[296])^(a[135] & b[297])^(a[134] & b[298])^(a[133] & b[299])^(a[132] & b[300])^(a[131] & b[301])^(a[130] & b[302])^(a[129] & b[303])^(a[128] & b[304])^(a[127] & b[305])^(a[126] & b[306])^(a[125] & b[307])^(a[124] & b[308])^(a[123] & b[309])^(a[122] & b[310])^(a[121] & b[311])^(a[120] & b[312])^(a[119] & b[313])^(a[118] & b[314])^(a[117] & b[315])^(a[116] & b[316])^(a[115] & b[317])^(a[114] & b[318])^(a[113] & b[319])^(a[112] & b[320])^(a[111] & b[321])^(a[110] & b[322])^(a[109] & b[323])^(a[108] & b[324])^(a[107] & b[325])^(a[106] & b[326])^(a[105] & b[327])^(a[104] & b[328])^(a[103] & b[329])^(a[102] & b[330])^(a[101] & b[331])^(a[100] & b[332])^(a[99] & b[333])^(a[98] & b[334])^(a[97] & b[335])^(a[96] & b[336])^(a[95] & b[337])^(a[94] & b[338])^(a[93] & b[339])^(a[92] & b[340])^(a[91] & b[341])^(a[90] & b[342])^(a[89] & b[343])^(a[88] & b[344])^(a[87] & b[345])^(a[86] & b[346])^(a[85] & b[347])^(a[84] & b[348])^(a[83] & b[349])^(a[82] & b[350])^(a[81] & b[351])^(a[80] & b[352])^(a[79] & b[353])^(a[78] & b[354])^(a[77] & b[355])^(a[76] & b[356])^(a[75] & b[357])^(a[74] & b[358])^(a[73] & b[359])^(a[72] & b[360])^(a[71] & b[361])^(a[70] & b[362])^(a[69] & b[363])^(a[68] & b[364])^(a[67] & b[365])^(a[66] & b[366])^(a[65] & b[367])^(a[64] & b[368])^(a[63] & b[369])^(a[62] & b[370])^(a[61] & b[371])^(a[60] & b[372])^(a[59] & b[373])^(a[58] & b[374])^(a[57] & b[375])^(a[56] & b[376])^(a[55] & b[377])^(a[54] & b[378])^(a[53] & b[379])^(a[52] & b[380])^(a[51] & b[381])^(a[50] & b[382])^(a[49] & b[383])^(a[48] & b[384])^(a[47] & b[385])^(a[46] & b[386])^(a[45] & b[387])^(a[44] & b[388])^(a[43] & b[389])^(a[42] & b[390])^(a[41] & b[391])^(a[40] & b[392])^(a[39] & b[393])^(a[38] & b[394])^(a[37] & b[395])^(a[36] & b[396])^(a[35] & b[397])^(a[34] & b[398])^(a[33] & b[399])^(a[32] & b[400])^(a[31] & b[401])^(a[30] & b[402])^(a[29] & b[403])^(a[28] & b[404])^(a[27] & b[405])^(a[26] & b[406])^(a[25] & b[407])^(a[24] & b[408]);
assign y[433] = (a[408] & b[25])^(a[407] & b[26])^(a[406] & b[27])^(a[405] & b[28])^(a[404] & b[29])^(a[403] & b[30])^(a[402] & b[31])^(a[401] & b[32])^(a[400] & b[33])^(a[399] & b[34])^(a[398] & b[35])^(a[397] & b[36])^(a[396] & b[37])^(a[395] & b[38])^(a[394] & b[39])^(a[393] & b[40])^(a[392] & b[41])^(a[391] & b[42])^(a[390] & b[43])^(a[389] & b[44])^(a[388] & b[45])^(a[387] & b[46])^(a[386] & b[47])^(a[385] & b[48])^(a[384] & b[49])^(a[383] & b[50])^(a[382] & b[51])^(a[381] & b[52])^(a[380] & b[53])^(a[379] & b[54])^(a[378] & b[55])^(a[377] & b[56])^(a[376] & b[57])^(a[375] & b[58])^(a[374] & b[59])^(a[373] & b[60])^(a[372] & b[61])^(a[371] & b[62])^(a[370] & b[63])^(a[369] & b[64])^(a[368] & b[65])^(a[367] & b[66])^(a[366] & b[67])^(a[365] & b[68])^(a[364] & b[69])^(a[363] & b[70])^(a[362] & b[71])^(a[361] & b[72])^(a[360] & b[73])^(a[359] & b[74])^(a[358] & b[75])^(a[357] & b[76])^(a[356] & b[77])^(a[355] & b[78])^(a[354] & b[79])^(a[353] & b[80])^(a[352] & b[81])^(a[351] & b[82])^(a[350] & b[83])^(a[349] & b[84])^(a[348] & b[85])^(a[347] & b[86])^(a[346] & b[87])^(a[345] & b[88])^(a[344] & b[89])^(a[343] & b[90])^(a[342] & b[91])^(a[341] & b[92])^(a[340] & b[93])^(a[339] & b[94])^(a[338] & b[95])^(a[337] & b[96])^(a[336] & b[97])^(a[335] & b[98])^(a[334] & b[99])^(a[333] & b[100])^(a[332] & b[101])^(a[331] & b[102])^(a[330] & b[103])^(a[329] & b[104])^(a[328] & b[105])^(a[327] & b[106])^(a[326] & b[107])^(a[325] & b[108])^(a[324] & b[109])^(a[323] & b[110])^(a[322] & b[111])^(a[321] & b[112])^(a[320] & b[113])^(a[319] & b[114])^(a[318] & b[115])^(a[317] & b[116])^(a[316] & b[117])^(a[315] & b[118])^(a[314] & b[119])^(a[313] & b[120])^(a[312] & b[121])^(a[311] & b[122])^(a[310] & b[123])^(a[309] & b[124])^(a[308] & b[125])^(a[307] & b[126])^(a[306] & b[127])^(a[305] & b[128])^(a[304] & b[129])^(a[303] & b[130])^(a[302] & b[131])^(a[301] & b[132])^(a[300] & b[133])^(a[299] & b[134])^(a[298] & b[135])^(a[297] & b[136])^(a[296] & b[137])^(a[295] & b[138])^(a[294] & b[139])^(a[293] & b[140])^(a[292] & b[141])^(a[291] & b[142])^(a[290] & b[143])^(a[289] & b[144])^(a[288] & b[145])^(a[287] & b[146])^(a[286] & b[147])^(a[285] & b[148])^(a[284] & b[149])^(a[283] & b[150])^(a[282] & b[151])^(a[281] & b[152])^(a[280] & b[153])^(a[279] & b[154])^(a[278] & b[155])^(a[277] & b[156])^(a[276] & b[157])^(a[275] & b[158])^(a[274] & b[159])^(a[273] & b[160])^(a[272] & b[161])^(a[271] & b[162])^(a[270] & b[163])^(a[269] & b[164])^(a[268] & b[165])^(a[267] & b[166])^(a[266] & b[167])^(a[265] & b[168])^(a[264] & b[169])^(a[263] & b[170])^(a[262] & b[171])^(a[261] & b[172])^(a[260] & b[173])^(a[259] & b[174])^(a[258] & b[175])^(a[257] & b[176])^(a[256] & b[177])^(a[255] & b[178])^(a[254] & b[179])^(a[253] & b[180])^(a[252] & b[181])^(a[251] & b[182])^(a[250] & b[183])^(a[249] & b[184])^(a[248] & b[185])^(a[247] & b[186])^(a[246] & b[187])^(a[245] & b[188])^(a[244] & b[189])^(a[243] & b[190])^(a[242] & b[191])^(a[241] & b[192])^(a[240] & b[193])^(a[239] & b[194])^(a[238] & b[195])^(a[237] & b[196])^(a[236] & b[197])^(a[235] & b[198])^(a[234] & b[199])^(a[233] & b[200])^(a[232] & b[201])^(a[231] & b[202])^(a[230] & b[203])^(a[229] & b[204])^(a[228] & b[205])^(a[227] & b[206])^(a[226] & b[207])^(a[225] & b[208])^(a[224] & b[209])^(a[223] & b[210])^(a[222] & b[211])^(a[221] & b[212])^(a[220] & b[213])^(a[219] & b[214])^(a[218] & b[215])^(a[217] & b[216])^(a[216] & b[217])^(a[215] & b[218])^(a[214] & b[219])^(a[213] & b[220])^(a[212] & b[221])^(a[211] & b[222])^(a[210] & b[223])^(a[209] & b[224])^(a[208] & b[225])^(a[207] & b[226])^(a[206] & b[227])^(a[205] & b[228])^(a[204] & b[229])^(a[203] & b[230])^(a[202] & b[231])^(a[201] & b[232])^(a[200] & b[233])^(a[199] & b[234])^(a[198] & b[235])^(a[197] & b[236])^(a[196] & b[237])^(a[195] & b[238])^(a[194] & b[239])^(a[193] & b[240])^(a[192] & b[241])^(a[191] & b[242])^(a[190] & b[243])^(a[189] & b[244])^(a[188] & b[245])^(a[187] & b[246])^(a[186] & b[247])^(a[185] & b[248])^(a[184] & b[249])^(a[183] & b[250])^(a[182] & b[251])^(a[181] & b[252])^(a[180] & b[253])^(a[179] & b[254])^(a[178] & b[255])^(a[177] & b[256])^(a[176] & b[257])^(a[175] & b[258])^(a[174] & b[259])^(a[173] & b[260])^(a[172] & b[261])^(a[171] & b[262])^(a[170] & b[263])^(a[169] & b[264])^(a[168] & b[265])^(a[167] & b[266])^(a[166] & b[267])^(a[165] & b[268])^(a[164] & b[269])^(a[163] & b[270])^(a[162] & b[271])^(a[161] & b[272])^(a[160] & b[273])^(a[159] & b[274])^(a[158] & b[275])^(a[157] & b[276])^(a[156] & b[277])^(a[155] & b[278])^(a[154] & b[279])^(a[153] & b[280])^(a[152] & b[281])^(a[151] & b[282])^(a[150] & b[283])^(a[149] & b[284])^(a[148] & b[285])^(a[147] & b[286])^(a[146] & b[287])^(a[145] & b[288])^(a[144] & b[289])^(a[143] & b[290])^(a[142] & b[291])^(a[141] & b[292])^(a[140] & b[293])^(a[139] & b[294])^(a[138] & b[295])^(a[137] & b[296])^(a[136] & b[297])^(a[135] & b[298])^(a[134] & b[299])^(a[133] & b[300])^(a[132] & b[301])^(a[131] & b[302])^(a[130] & b[303])^(a[129] & b[304])^(a[128] & b[305])^(a[127] & b[306])^(a[126] & b[307])^(a[125] & b[308])^(a[124] & b[309])^(a[123] & b[310])^(a[122] & b[311])^(a[121] & b[312])^(a[120] & b[313])^(a[119] & b[314])^(a[118] & b[315])^(a[117] & b[316])^(a[116] & b[317])^(a[115] & b[318])^(a[114] & b[319])^(a[113] & b[320])^(a[112] & b[321])^(a[111] & b[322])^(a[110] & b[323])^(a[109] & b[324])^(a[108] & b[325])^(a[107] & b[326])^(a[106] & b[327])^(a[105] & b[328])^(a[104] & b[329])^(a[103] & b[330])^(a[102] & b[331])^(a[101] & b[332])^(a[100] & b[333])^(a[99] & b[334])^(a[98] & b[335])^(a[97] & b[336])^(a[96] & b[337])^(a[95] & b[338])^(a[94] & b[339])^(a[93] & b[340])^(a[92] & b[341])^(a[91] & b[342])^(a[90] & b[343])^(a[89] & b[344])^(a[88] & b[345])^(a[87] & b[346])^(a[86] & b[347])^(a[85] & b[348])^(a[84] & b[349])^(a[83] & b[350])^(a[82] & b[351])^(a[81] & b[352])^(a[80] & b[353])^(a[79] & b[354])^(a[78] & b[355])^(a[77] & b[356])^(a[76] & b[357])^(a[75] & b[358])^(a[74] & b[359])^(a[73] & b[360])^(a[72] & b[361])^(a[71] & b[362])^(a[70] & b[363])^(a[69] & b[364])^(a[68] & b[365])^(a[67] & b[366])^(a[66] & b[367])^(a[65] & b[368])^(a[64] & b[369])^(a[63] & b[370])^(a[62] & b[371])^(a[61] & b[372])^(a[60] & b[373])^(a[59] & b[374])^(a[58] & b[375])^(a[57] & b[376])^(a[56] & b[377])^(a[55] & b[378])^(a[54] & b[379])^(a[53] & b[380])^(a[52] & b[381])^(a[51] & b[382])^(a[50] & b[383])^(a[49] & b[384])^(a[48] & b[385])^(a[47] & b[386])^(a[46] & b[387])^(a[45] & b[388])^(a[44] & b[389])^(a[43] & b[390])^(a[42] & b[391])^(a[41] & b[392])^(a[40] & b[393])^(a[39] & b[394])^(a[38] & b[395])^(a[37] & b[396])^(a[36] & b[397])^(a[35] & b[398])^(a[34] & b[399])^(a[33] & b[400])^(a[32] & b[401])^(a[31] & b[402])^(a[30] & b[403])^(a[29] & b[404])^(a[28] & b[405])^(a[27] & b[406])^(a[26] & b[407])^(a[25] & b[408]);
assign y[434] = (a[408] & b[26])^(a[407] & b[27])^(a[406] & b[28])^(a[405] & b[29])^(a[404] & b[30])^(a[403] & b[31])^(a[402] & b[32])^(a[401] & b[33])^(a[400] & b[34])^(a[399] & b[35])^(a[398] & b[36])^(a[397] & b[37])^(a[396] & b[38])^(a[395] & b[39])^(a[394] & b[40])^(a[393] & b[41])^(a[392] & b[42])^(a[391] & b[43])^(a[390] & b[44])^(a[389] & b[45])^(a[388] & b[46])^(a[387] & b[47])^(a[386] & b[48])^(a[385] & b[49])^(a[384] & b[50])^(a[383] & b[51])^(a[382] & b[52])^(a[381] & b[53])^(a[380] & b[54])^(a[379] & b[55])^(a[378] & b[56])^(a[377] & b[57])^(a[376] & b[58])^(a[375] & b[59])^(a[374] & b[60])^(a[373] & b[61])^(a[372] & b[62])^(a[371] & b[63])^(a[370] & b[64])^(a[369] & b[65])^(a[368] & b[66])^(a[367] & b[67])^(a[366] & b[68])^(a[365] & b[69])^(a[364] & b[70])^(a[363] & b[71])^(a[362] & b[72])^(a[361] & b[73])^(a[360] & b[74])^(a[359] & b[75])^(a[358] & b[76])^(a[357] & b[77])^(a[356] & b[78])^(a[355] & b[79])^(a[354] & b[80])^(a[353] & b[81])^(a[352] & b[82])^(a[351] & b[83])^(a[350] & b[84])^(a[349] & b[85])^(a[348] & b[86])^(a[347] & b[87])^(a[346] & b[88])^(a[345] & b[89])^(a[344] & b[90])^(a[343] & b[91])^(a[342] & b[92])^(a[341] & b[93])^(a[340] & b[94])^(a[339] & b[95])^(a[338] & b[96])^(a[337] & b[97])^(a[336] & b[98])^(a[335] & b[99])^(a[334] & b[100])^(a[333] & b[101])^(a[332] & b[102])^(a[331] & b[103])^(a[330] & b[104])^(a[329] & b[105])^(a[328] & b[106])^(a[327] & b[107])^(a[326] & b[108])^(a[325] & b[109])^(a[324] & b[110])^(a[323] & b[111])^(a[322] & b[112])^(a[321] & b[113])^(a[320] & b[114])^(a[319] & b[115])^(a[318] & b[116])^(a[317] & b[117])^(a[316] & b[118])^(a[315] & b[119])^(a[314] & b[120])^(a[313] & b[121])^(a[312] & b[122])^(a[311] & b[123])^(a[310] & b[124])^(a[309] & b[125])^(a[308] & b[126])^(a[307] & b[127])^(a[306] & b[128])^(a[305] & b[129])^(a[304] & b[130])^(a[303] & b[131])^(a[302] & b[132])^(a[301] & b[133])^(a[300] & b[134])^(a[299] & b[135])^(a[298] & b[136])^(a[297] & b[137])^(a[296] & b[138])^(a[295] & b[139])^(a[294] & b[140])^(a[293] & b[141])^(a[292] & b[142])^(a[291] & b[143])^(a[290] & b[144])^(a[289] & b[145])^(a[288] & b[146])^(a[287] & b[147])^(a[286] & b[148])^(a[285] & b[149])^(a[284] & b[150])^(a[283] & b[151])^(a[282] & b[152])^(a[281] & b[153])^(a[280] & b[154])^(a[279] & b[155])^(a[278] & b[156])^(a[277] & b[157])^(a[276] & b[158])^(a[275] & b[159])^(a[274] & b[160])^(a[273] & b[161])^(a[272] & b[162])^(a[271] & b[163])^(a[270] & b[164])^(a[269] & b[165])^(a[268] & b[166])^(a[267] & b[167])^(a[266] & b[168])^(a[265] & b[169])^(a[264] & b[170])^(a[263] & b[171])^(a[262] & b[172])^(a[261] & b[173])^(a[260] & b[174])^(a[259] & b[175])^(a[258] & b[176])^(a[257] & b[177])^(a[256] & b[178])^(a[255] & b[179])^(a[254] & b[180])^(a[253] & b[181])^(a[252] & b[182])^(a[251] & b[183])^(a[250] & b[184])^(a[249] & b[185])^(a[248] & b[186])^(a[247] & b[187])^(a[246] & b[188])^(a[245] & b[189])^(a[244] & b[190])^(a[243] & b[191])^(a[242] & b[192])^(a[241] & b[193])^(a[240] & b[194])^(a[239] & b[195])^(a[238] & b[196])^(a[237] & b[197])^(a[236] & b[198])^(a[235] & b[199])^(a[234] & b[200])^(a[233] & b[201])^(a[232] & b[202])^(a[231] & b[203])^(a[230] & b[204])^(a[229] & b[205])^(a[228] & b[206])^(a[227] & b[207])^(a[226] & b[208])^(a[225] & b[209])^(a[224] & b[210])^(a[223] & b[211])^(a[222] & b[212])^(a[221] & b[213])^(a[220] & b[214])^(a[219] & b[215])^(a[218] & b[216])^(a[217] & b[217])^(a[216] & b[218])^(a[215] & b[219])^(a[214] & b[220])^(a[213] & b[221])^(a[212] & b[222])^(a[211] & b[223])^(a[210] & b[224])^(a[209] & b[225])^(a[208] & b[226])^(a[207] & b[227])^(a[206] & b[228])^(a[205] & b[229])^(a[204] & b[230])^(a[203] & b[231])^(a[202] & b[232])^(a[201] & b[233])^(a[200] & b[234])^(a[199] & b[235])^(a[198] & b[236])^(a[197] & b[237])^(a[196] & b[238])^(a[195] & b[239])^(a[194] & b[240])^(a[193] & b[241])^(a[192] & b[242])^(a[191] & b[243])^(a[190] & b[244])^(a[189] & b[245])^(a[188] & b[246])^(a[187] & b[247])^(a[186] & b[248])^(a[185] & b[249])^(a[184] & b[250])^(a[183] & b[251])^(a[182] & b[252])^(a[181] & b[253])^(a[180] & b[254])^(a[179] & b[255])^(a[178] & b[256])^(a[177] & b[257])^(a[176] & b[258])^(a[175] & b[259])^(a[174] & b[260])^(a[173] & b[261])^(a[172] & b[262])^(a[171] & b[263])^(a[170] & b[264])^(a[169] & b[265])^(a[168] & b[266])^(a[167] & b[267])^(a[166] & b[268])^(a[165] & b[269])^(a[164] & b[270])^(a[163] & b[271])^(a[162] & b[272])^(a[161] & b[273])^(a[160] & b[274])^(a[159] & b[275])^(a[158] & b[276])^(a[157] & b[277])^(a[156] & b[278])^(a[155] & b[279])^(a[154] & b[280])^(a[153] & b[281])^(a[152] & b[282])^(a[151] & b[283])^(a[150] & b[284])^(a[149] & b[285])^(a[148] & b[286])^(a[147] & b[287])^(a[146] & b[288])^(a[145] & b[289])^(a[144] & b[290])^(a[143] & b[291])^(a[142] & b[292])^(a[141] & b[293])^(a[140] & b[294])^(a[139] & b[295])^(a[138] & b[296])^(a[137] & b[297])^(a[136] & b[298])^(a[135] & b[299])^(a[134] & b[300])^(a[133] & b[301])^(a[132] & b[302])^(a[131] & b[303])^(a[130] & b[304])^(a[129] & b[305])^(a[128] & b[306])^(a[127] & b[307])^(a[126] & b[308])^(a[125] & b[309])^(a[124] & b[310])^(a[123] & b[311])^(a[122] & b[312])^(a[121] & b[313])^(a[120] & b[314])^(a[119] & b[315])^(a[118] & b[316])^(a[117] & b[317])^(a[116] & b[318])^(a[115] & b[319])^(a[114] & b[320])^(a[113] & b[321])^(a[112] & b[322])^(a[111] & b[323])^(a[110] & b[324])^(a[109] & b[325])^(a[108] & b[326])^(a[107] & b[327])^(a[106] & b[328])^(a[105] & b[329])^(a[104] & b[330])^(a[103] & b[331])^(a[102] & b[332])^(a[101] & b[333])^(a[100] & b[334])^(a[99] & b[335])^(a[98] & b[336])^(a[97] & b[337])^(a[96] & b[338])^(a[95] & b[339])^(a[94] & b[340])^(a[93] & b[341])^(a[92] & b[342])^(a[91] & b[343])^(a[90] & b[344])^(a[89] & b[345])^(a[88] & b[346])^(a[87] & b[347])^(a[86] & b[348])^(a[85] & b[349])^(a[84] & b[350])^(a[83] & b[351])^(a[82] & b[352])^(a[81] & b[353])^(a[80] & b[354])^(a[79] & b[355])^(a[78] & b[356])^(a[77] & b[357])^(a[76] & b[358])^(a[75] & b[359])^(a[74] & b[360])^(a[73] & b[361])^(a[72] & b[362])^(a[71] & b[363])^(a[70] & b[364])^(a[69] & b[365])^(a[68] & b[366])^(a[67] & b[367])^(a[66] & b[368])^(a[65] & b[369])^(a[64] & b[370])^(a[63] & b[371])^(a[62] & b[372])^(a[61] & b[373])^(a[60] & b[374])^(a[59] & b[375])^(a[58] & b[376])^(a[57] & b[377])^(a[56] & b[378])^(a[55] & b[379])^(a[54] & b[380])^(a[53] & b[381])^(a[52] & b[382])^(a[51] & b[383])^(a[50] & b[384])^(a[49] & b[385])^(a[48] & b[386])^(a[47] & b[387])^(a[46] & b[388])^(a[45] & b[389])^(a[44] & b[390])^(a[43] & b[391])^(a[42] & b[392])^(a[41] & b[393])^(a[40] & b[394])^(a[39] & b[395])^(a[38] & b[396])^(a[37] & b[397])^(a[36] & b[398])^(a[35] & b[399])^(a[34] & b[400])^(a[33] & b[401])^(a[32] & b[402])^(a[31] & b[403])^(a[30] & b[404])^(a[29] & b[405])^(a[28] & b[406])^(a[27] & b[407])^(a[26] & b[408]);
assign y[435] = (a[408] & b[27])^(a[407] & b[28])^(a[406] & b[29])^(a[405] & b[30])^(a[404] & b[31])^(a[403] & b[32])^(a[402] & b[33])^(a[401] & b[34])^(a[400] & b[35])^(a[399] & b[36])^(a[398] & b[37])^(a[397] & b[38])^(a[396] & b[39])^(a[395] & b[40])^(a[394] & b[41])^(a[393] & b[42])^(a[392] & b[43])^(a[391] & b[44])^(a[390] & b[45])^(a[389] & b[46])^(a[388] & b[47])^(a[387] & b[48])^(a[386] & b[49])^(a[385] & b[50])^(a[384] & b[51])^(a[383] & b[52])^(a[382] & b[53])^(a[381] & b[54])^(a[380] & b[55])^(a[379] & b[56])^(a[378] & b[57])^(a[377] & b[58])^(a[376] & b[59])^(a[375] & b[60])^(a[374] & b[61])^(a[373] & b[62])^(a[372] & b[63])^(a[371] & b[64])^(a[370] & b[65])^(a[369] & b[66])^(a[368] & b[67])^(a[367] & b[68])^(a[366] & b[69])^(a[365] & b[70])^(a[364] & b[71])^(a[363] & b[72])^(a[362] & b[73])^(a[361] & b[74])^(a[360] & b[75])^(a[359] & b[76])^(a[358] & b[77])^(a[357] & b[78])^(a[356] & b[79])^(a[355] & b[80])^(a[354] & b[81])^(a[353] & b[82])^(a[352] & b[83])^(a[351] & b[84])^(a[350] & b[85])^(a[349] & b[86])^(a[348] & b[87])^(a[347] & b[88])^(a[346] & b[89])^(a[345] & b[90])^(a[344] & b[91])^(a[343] & b[92])^(a[342] & b[93])^(a[341] & b[94])^(a[340] & b[95])^(a[339] & b[96])^(a[338] & b[97])^(a[337] & b[98])^(a[336] & b[99])^(a[335] & b[100])^(a[334] & b[101])^(a[333] & b[102])^(a[332] & b[103])^(a[331] & b[104])^(a[330] & b[105])^(a[329] & b[106])^(a[328] & b[107])^(a[327] & b[108])^(a[326] & b[109])^(a[325] & b[110])^(a[324] & b[111])^(a[323] & b[112])^(a[322] & b[113])^(a[321] & b[114])^(a[320] & b[115])^(a[319] & b[116])^(a[318] & b[117])^(a[317] & b[118])^(a[316] & b[119])^(a[315] & b[120])^(a[314] & b[121])^(a[313] & b[122])^(a[312] & b[123])^(a[311] & b[124])^(a[310] & b[125])^(a[309] & b[126])^(a[308] & b[127])^(a[307] & b[128])^(a[306] & b[129])^(a[305] & b[130])^(a[304] & b[131])^(a[303] & b[132])^(a[302] & b[133])^(a[301] & b[134])^(a[300] & b[135])^(a[299] & b[136])^(a[298] & b[137])^(a[297] & b[138])^(a[296] & b[139])^(a[295] & b[140])^(a[294] & b[141])^(a[293] & b[142])^(a[292] & b[143])^(a[291] & b[144])^(a[290] & b[145])^(a[289] & b[146])^(a[288] & b[147])^(a[287] & b[148])^(a[286] & b[149])^(a[285] & b[150])^(a[284] & b[151])^(a[283] & b[152])^(a[282] & b[153])^(a[281] & b[154])^(a[280] & b[155])^(a[279] & b[156])^(a[278] & b[157])^(a[277] & b[158])^(a[276] & b[159])^(a[275] & b[160])^(a[274] & b[161])^(a[273] & b[162])^(a[272] & b[163])^(a[271] & b[164])^(a[270] & b[165])^(a[269] & b[166])^(a[268] & b[167])^(a[267] & b[168])^(a[266] & b[169])^(a[265] & b[170])^(a[264] & b[171])^(a[263] & b[172])^(a[262] & b[173])^(a[261] & b[174])^(a[260] & b[175])^(a[259] & b[176])^(a[258] & b[177])^(a[257] & b[178])^(a[256] & b[179])^(a[255] & b[180])^(a[254] & b[181])^(a[253] & b[182])^(a[252] & b[183])^(a[251] & b[184])^(a[250] & b[185])^(a[249] & b[186])^(a[248] & b[187])^(a[247] & b[188])^(a[246] & b[189])^(a[245] & b[190])^(a[244] & b[191])^(a[243] & b[192])^(a[242] & b[193])^(a[241] & b[194])^(a[240] & b[195])^(a[239] & b[196])^(a[238] & b[197])^(a[237] & b[198])^(a[236] & b[199])^(a[235] & b[200])^(a[234] & b[201])^(a[233] & b[202])^(a[232] & b[203])^(a[231] & b[204])^(a[230] & b[205])^(a[229] & b[206])^(a[228] & b[207])^(a[227] & b[208])^(a[226] & b[209])^(a[225] & b[210])^(a[224] & b[211])^(a[223] & b[212])^(a[222] & b[213])^(a[221] & b[214])^(a[220] & b[215])^(a[219] & b[216])^(a[218] & b[217])^(a[217] & b[218])^(a[216] & b[219])^(a[215] & b[220])^(a[214] & b[221])^(a[213] & b[222])^(a[212] & b[223])^(a[211] & b[224])^(a[210] & b[225])^(a[209] & b[226])^(a[208] & b[227])^(a[207] & b[228])^(a[206] & b[229])^(a[205] & b[230])^(a[204] & b[231])^(a[203] & b[232])^(a[202] & b[233])^(a[201] & b[234])^(a[200] & b[235])^(a[199] & b[236])^(a[198] & b[237])^(a[197] & b[238])^(a[196] & b[239])^(a[195] & b[240])^(a[194] & b[241])^(a[193] & b[242])^(a[192] & b[243])^(a[191] & b[244])^(a[190] & b[245])^(a[189] & b[246])^(a[188] & b[247])^(a[187] & b[248])^(a[186] & b[249])^(a[185] & b[250])^(a[184] & b[251])^(a[183] & b[252])^(a[182] & b[253])^(a[181] & b[254])^(a[180] & b[255])^(a[179] & b[256])^(a[178] & b[257])^(a[177] & b[258])^(a[176] & b[259])^(a[175] & b[260])^(a[174] & b[261])^(a[173] & b[262])^(a[172] & b[263])^(a[171] & b[264])^(a[170] & b[265])^(a[169] & b[266])^(a[168] & b[267])^(a[167] & b[268])^(a[166] & b[269])^(a[165] & b[270])^(a[164] & b[271])^(a[163] & b[272])^(a[162] & b[273])^(a[161] & b[274])^(a[160] & b[275])^(a[159] & b[276])^(a[158] & b[277])^(a[157] & b[278])^(a[156] & b[279])^(a[155] & b[280])^(a[154] & b[281])^(a[153] & b[282])^(a[152] & b[283])^(a[151] & b[284])^(a[150] & b[285])^(a[149] & b[286])^(a[148] & b[287])^(a[147] & b[288])^(a[146] & b[289])^(a[145] & b[290])^(a[144] & b[291])^(a[143] & b[292])^(a[142] & b[293])^(a[141] & b[294])^(a[140] & b[295])^(a[139] & b[296])^(a[138] & b[297])^(a[137] & b[298])^(a[136] & b[299])^(a[135] & b[300])^(a[134] & b[301])^(a[133] & b[302])^(a[132] & b[303])^(a[131] & b[304])^(a[130] & b[305])^(a[129] & b[306])^(a[128] & b[307])^(a[127] & b[308])^(a[126] & b[309])^(a[125] & b[310])^(a[124] & b[311])^(a[123] & b[312])^(a[122] & b[313])^(a[121] & b[314])^(a[120] & b[315])^(a[119] & b[316])^(a[118] & b[317])^(a[117] & b[318])^(a[116] & b[319])^(a[115] & b[320])^(a[114] & b[321])^(a[113] & b[322])^(a[112] & b[323])^(a[111] & b[324])^(a[110] & b[325])^(a[109] & b[326])^(a[108] & b[327])^(a[107] & b[328])^(a[106] & b[329])^(a[105] & b[330])^(a[104] & b[331])^(a[103] & b[332])^(a[102] & b[333])^(a[101] & b[334])^(a[100] & b[335])^(a[99] & b[336])^(a[98] & b[337])^(a[97] & b[338])^(a[96] & b[339])^(a[95] & b[340])^(a[94] & b[341])^(a[93] & b[342])^(a[92] & b[343])^(a[91] & b[344])^(a[90] & b[345])^(a[89] & b[346])^(a[88] & b[347])^(a[87] & b[348])^(a[86] & b[349])^(a[85] & b[350])^(a[84] & b[351])^(a[83] & b[352])^(a[82] & b[353])^(a[81] & b[354])^(a[80] & b[355])^(a[79] & b[356])^(a[78] & b[357])^(a[77] & b[358])^(a[76] & b[359])^(a[75] & b[360])^(a[74] & b[361])^(a[73] & b[362])^(a[72] & b[363])^(a[71] & b[364])^(a[70] & b[365])^(a[69] & b[366])^(a[68] & b[367])^(a[67] & b[368])^(a[66] & b[369])^(a[65] & b[370])^(a[64] & b[371])^(a[63] & b[372])^(a[62] & b[373])^(a[61] & b[374])^(a[60] & b[375])^(a[59] & b[376])^(a[58] & b[377])^(a[57] & b[378])^(a[56] & b[379])^(a[55] & b[380])^(a[54] & b[381])^(a[53] & b[382])^(a[52] & b[383])^(a[51] & b[384])^(a[50] & b[385])^(a[49] & b[386])^(a[48] & b[387])^(a[47] & b[388])^(a[46] & b[389])^(a[45] & b[390])^(a[44] & b[391])^(a[43] & b[392])^(a[42] & b[393])^(a[41] & b[394])^(a[40] & b[395])^(a[39] & b[396])^(a[38] & b[397])^(a[37] & b[398])^(a[36] & b[399])^(a[35] & b[400])^(a[34] & b[401])^(a[33] & b[402])^(a[32] & b[403])^(a[31] & b[404])^(a[30] & b[405])^(a[29] & b[406])^(a[28] & b[407])^(a[27] & b[408]);
assign y[436] = (a[408] & b[28])^(a[407] & b[29])^(a[406] & b[30])^(a[405] & b[31])^(a[404] & b[32])^(a[403] & b[33])^(a[402] & b[34])^(a[401] & b[35])^(a[400] & b[36])^(a[399] & b[37])^(a[398] & b[38])^(a[397] & b[39])^(a[396] & b[40])^(a[395] & b[41])^(a[394] & b[42])^(a[393] & b[43])^(a[392] & b[44])^(a[391] & b[45])^(a[390] & b[46])^(a[389] & b[47])^(a[388] & b[48])^(a[387] & b[49])^(a[386] & b[50])^(a[385] & b[51])^(a[384] & b[52])^(a[383] & b[53])^(a[382] & b[54])^(a[381] & b[55])^(a[380] & b[56])^(a[379] & b[57])^(a[378] & b[58])^(a[377] & b[59])^(a[376] & b[60])^(a[375] & b[61])^(a[374] & b[62])^(a[373] & b[63])^(a[372] & b[64])^(a[371] & b[65])^(a[370] & b[66])^(a[369] & b[67])^(a[368] & b[68])^(a[367] & b[69])^(a[366] & b[70])^(a[365] & b[71])^(a[364] & b[72])^(a[363] & b[73])^(a[362] & b[74])^(a[361] & b[75])^(a[360] & b[76])^(a[359] & b[77])^(a[358] & b[78])^(a[357] & b[79])^(a[356] & b[80])^(a[355] & b[81])^(a[354] & b[82])^(a[353] & b[83])^(a[352] & b[84])^(a[351] & b[85])^(a[350] & b[86])^(a[349] & b[87])^(a[348] & b[88])^(a[347] & b[89])^(a[346] & b[90])^(a[345] & b[91])^(a[344] & b[92])^(a[343] & b[93])^(a[342] & b[94])^(a[341] & b[95])^(a[340] & b[96])^(a[339] & b[97])^(a[338] & b[98])^(a[337] & b[99])^(a[336] & b[100])^(a[335] & b[101])^(a[334] & b[102])^(a[333] & b[103])^(a[332] & b[104])^(a[331] & b[105])^(a[330] & b[106])^(a[329] & b[107])^(a[328] & b[108])^(a[327] & b[109])^(a[326] & b[110])^(a[325] & b[111])^(a[324] & b[112])^(a[323] & b[113])^(a[322] & b[114])^(a[321] & b[115])^(a[320] & b[116])^(a[319] & b[117])^(a[318] & b[118])^(a[317] & b[119])^(a[316] & b[120])^(a[315] & b[121])^(a[314] & b[122])^(a[313] & b[123])^(a[312] & b[124])^(a[311] & b[125])^(a[310] & b[126])^(a[309] & b[127])^(a[308] & b[128])^(a[307] & b[129])^(a[306] & b[130])^(a[305] & b[131])^(a[304] & b[132])^(a[303] & b[133])^(a[302] & b[134])^(a[301] & b[135])^(a[300] & b[136])^(a[299] & b[137])^(a[298] & b[138])^(a[297] & b[139])^(a[296] & b[140])^(a[295] & b[141])^(a[294] & b[142])^(a[293] & b[143])^(a[292] & b[144])^(a[291] & b[145])^(a[290] & b[146])^(a[289] & b[147])^(a[288] & b[148])^(a[287] & b[149])^(a[286] & b[150])^(a[285] & b[151])^(a[284] & b[152])^(a[283] & b[153])^(a[282] & b[154])^(a[281] & b[155])^(a[280] & b[156])^(a[279] & b[157])^(a[278] & b[158])^(a[277] & b[159])^(a[276] & b[160])^(a[275] & b[161])^(a[274] & b[162])^(a[273] & b[163])^(a[272] & b[164])^(a[271] & b[165])^(a[270] & b[166])^(a[269] & b[167])^(a[268] & b[168])^(a[267] & b[169])^(a[266] & b[170])^(a[265] & b[171])^(a[264] & b[172])^(a[263] & b[173])^(a[262] & b[174])^(a[261] & b[175])^(a[260] & b[176])^(a[259] & b[177])^(a[258] & b[178])^(a[257] & b[179])^(a[256] & b[180])^(a[255] & b[181])^(a[254] & b[182])^(a[253] & b[183])^(a[252] & b[184])^(a[251] & b[185])^(a[250] & b[186])^(a[249] & b[187])^(a[248] & b[188])^(a[247] & b[189])^(a[246] & b[190])^(a[245] & b[191])^(a[244] & b[192])^(a[243] & b[193])^(a[242] & b[194])^(a[241] & b[195])^(a[240] & b[196])^(a[239] & b[197])^(a[238] & b[198])^(a[237] & b[199])^(a[236] & b[200])^(a[235] & b[201])^(a[234] & b[202])^(a[233] & b[203])^(a[232] & b[204])^(a[231] & b[205])^(a[230] & b[206])^(a[229] & b[207])^(a[228] & b[208])^(a[227] & b[209])^(a[226] & b[210])^(a[225] & b[211])^(a[224] & b[212])^(a[223] & b[213])^(a[222] & b[214])^(a[221] & b[215])^(a[220] & b[216])^(a[219] & b[217])^(a[218] & b[218])^(a[217] & b[219])^(a[216] & b[220])^(a[215] & b[221])^(a[214] & b[222])^(a[213] & b[223])^(a[212] & b[224])^(a[211] & b[225])^(a[210] & b[226])^(a[209] & b[227])^(a[208] & b[228])^(a[207] & b[229])^(a[206] & b[230])^(a[205] & b[231])^(a[204] & b[232])^(a[203] & b[233])^(a[202] & b[234])^(a[201] & b[235])^(a[200] & b[236])^(a[199] & b[237])^(a[198] & b[238])^(a[197] & b[239])^(a[196] & b[240])^(a[195] & b[241])^(a[194] & b[242])^(a[193] & b[243])^(a[192] & b[244])^(a[191] & b[245])^(a[190] & b[246])^(a[189] & b[247])^(a[188] & b[248])^(a[187] & b[249])^(a[186] & b[250])^(a[185] & b[251])^(a[184] & b[252])^(a[183] & b[253])^(a[182] & b[254])^(a[181] & b[255])^(a[180] & b[256])^(a[179] & b[257])^(a[178] & b[258])^(a[177] & b[259])^(a[176] & b[260])^(a[175] & b[261])^(a[174] & b[262])^(a[173] & b[263])^(a[172] & b[264])^(a[171] & b[265])^(a[170] & b[266])^(a[169] & b[267])^(a[168] & b[268])^(a[167] & b[269])^(a[166] & b[270])^(a[165] & b[271])^(a[164] & b[272])^(a[163] & b[273])^(a[162] & b[274])^(a[161] & b[275])^(a[160] & b[276])^(a[159] & b[277])^(a[158] & b[278])^(a[157] & b[279])^(a[156] & b[280])^(a[155] & b[281])^(a[154] & b[282])^(a[153] & b[283])^(a[152] & b[284])^(a[151] & b[285])^(a[150] & b[286])^(a[149] & b[287])^(a[148] & b[288])^(a[147] & b[289])^(a[146] & b[290])^(a[145] & b[291])^(a[144] & b[292])^(a[143] & b[293])^(a[142] & b[294])^(a[141] & b[295])^(a[140] & b[296])^(a[139] & b[297])^(a[138] & b[298])^(a[137] & b[299])^(a[136] & b[300])^(a[135] & b[301])^(a[134] & b[302])^(a[133] & b[303])^(a[132] & b[304])^(a[131] & b[305])^(a[130] & b[306])^(a[129] & b[307])^(a[128] & b[308])^(a[127] & b[309])^(a[126] & b[310])^(a[125] & b[311])^(a[124] & b[312])^(a[123] & b[313])^(a[122] & b[314])^(a[121] & b[315])^(a[120] & b[316])^(a[119] & b[317])^(a[118] & b[318])^(a[117] & b[319])^(a[116] & b[320])^(a[115] & b[321])^(a[114] & b[322])^(a[113] & b[323])^(a[112] & b[324])^(a[111] & b[325])^(a[110] & b[326])^(a[109] & b[327])^(a[108] & b[328])^(a[107] & b[329])^(a[106] & b[330])^(a[105] & b[331])^(a[104] & b[332])^(a[103] & b[333])^(a[102] & b[334])^(a[101] & b[335])^(a[100] & b[336])^(a[99] & b[337])^(a[98] & b[338])^(a[97] & b[339])^(a[96] & b[340])^(a[95] & b[341])^(a[94] & b[342])^(a[93] & b[343])^(a[92] & b[344])^(a[91] & b[345])^(a[90] & b[346])^(a[89] & b[347])^(a[88] & b[348])^(a[87] & b[349])^(a[86] & b[350])^(a[85] & b[351])^(a[84] & b[352])^(a[83] & b[353])^(a[82] & b[354])^(a[81] & b[355])^(a[80] & b[356])^(a[79] & b[357])^(a[78] & b[358])^(a[77] & b[359])^(a[76] & b[360])^(a[75] & b[361])^(a[74] & b[362])^(a[73] & b[363])^(a[72] & b[364])^(a[71] & b[365])^(a[70] & b[366])^(a[69] & b[367])^(a[68] & b[368])^(a[67] & b[369])^(a[66] & b[370])^(a[65] & b[371])^(a[64] & b[372])^(a[63] & b[373])^(a[62] & b[374])^(a[61] & b[375])^(a[60] & b[376])^(a[59] & b[377])^(a[58] & b[378])^(a[57] & b[379])^(a[56] & b[380])^(a[55] & b[381])^(a[54] & b[382])^(a[53] & b[383])^(a[52] & b[384])^(a[51] & b[385])^(a[50] & b[386])^(a[49] & b[387])^(a[48] & b[388])^(a[47] & b[389])^(a[46] & b[390])^(a[45] & b[391])^(a[44] & b[392])^(a[43] & b[393])^(a[42] & b[394])^(a[41] & b[395])^(a[40] & b[396])^(a[39] & b[397])^(a[38] & b[398])^(a[37] & b[399])^(a[36] & b[400])^(a[35] & b[401])^(a[34] & b[402])^(a[33] & b[403])^(a[32] & b[404])^(a[31] & b[405])^(a[30] & b[406])^(a[29] & b[407])^(a[28] & b[408]);
assign y[437] = (a[408] & b[29])^(a[407] & b[30])^(a[406] & b[31])^(a[405] & b[32])^(a[404] & b[33])^(a[403] & b[34])^(a[402] & b[35])^(a[401] & b[36])^(a[400] & b[37])^(a[399] & b[38])^(a[398] & b[39])^(a[397] & b[40])^(a[396] & b[41])^(a[395] & b[42])^(a[394] & b[43])^(a[393] & b[44])^(a[392] & b[45])^(a[391] & b[46])^(a[390] & b[47])^(a[389] & b[48])^(a[388] & b[49])^(a[387] & b[50])^(a[386] & b[51])^(a[385] & b[52])^(a[384] & b[53])^(a[383] & b[54])^(a[382] & b[55])^(a[381] & b[56])^(a[380] & b[57])^(a[379] & b[58])^(a[378] & b[59])^(a[377] & b[60])^(a[376] & b[61])^(a[375] & b[62])^(a[374] & b[63])^(a[373] & b[64])^(a[372] & b[65])^(a[371] & b[66])^(a[370] & b[67])^(a[369] & b[68])^(a[368] & b[69])^(a[367] & b[70])^(a[366] & b[71])^(a[365] & b[72])^(a[364] & b[73])^(a[363] & b[74])^(a[362] & b[75])^(a[361] & b[76])^(a[360] & b[77])^(a[359] & b[78])^(a[358] & b[79])^(a[357] & b[80])^(a[356] & b[81])^(a[355] & b[82])^(a[354] & b[83])^(a[353] & b[84])^(a[352] & b[85])^(a[351] & b[86])^(a[350] & b[87])^(a[349] & b[88])^(a[348] & b[89])^(a[347] & b[90])^(a[346] & b[91])^(a[345] & b[92])^(a[344] & b[93])^(a[343] & b[94])^(a[342] & b[95])^(a[341] & b[96])^(a[340] & b[97])^(a[339] & b[98])^(a[338] & b[99])^(a[337] & b[100])^(a[336] & b[101])^(a[335] & b[102])^(a[334] & b[103])^(a[333] & b[104])^(a[332] & b[105])^(a[331] & b[106])^(a[330] & b[107])^(a[329] & b[108])^(a[328] & b[109])^(a[327] & b[110])^(a[326] & b[111])^(a[325] & b[112])^(a[324] & b[113])^(a[323] & b[114])^(a[322] & b[115])^(a[321] & b[116])^(a[320] & b[117])^(a[319] & b[118])^(a[318] & b[119])^(a[317] & b[120])^(a[316] & b[121])^(a[315] & b[122])^(a[314] & b[123])^(a[313] & b[124])^(a[312] & b[125])^(a[311] & b[126])^(a[310] & b[127])^(a[309] & b[128])^(a[308] & b[129])^(a[307] & b[130])^(a[306] & b[131])^(a[305] & b[132])^(a[304] & b[133])^(a[303] & b[134])^(a[302] & b[135])^(a[301] & b[136])^(a[300] & b[137])^(a[299] & b[138])^(a[298] & b[139])^(a[297] & b[140])^(a[296] & b[141])^(a[295] & b[142])^(a[294] & b[143])^(a[293] & b[144])^(a[292] & b[145])^(a[291] & b[146])^(a[290] & b[147])^(a[289] & b[148])^(a[288] & b[149])^(a[287] & b[150])^(a[286] & b[151])^(a[285] & b[152])^(a[284] & b[153])^(a[283] & b[154])^(a[282] & b[155])^(a[281] & b[156])^(a[280] & b[157])^(a[279] & b[158])^(a[278] & b[159])^(a[277] & b[160])^(a[276] & b[161])^(a[275] & b[162])^(a[274] & b[163])^(a[273] & b[164])^(a[272] & b[165])^(a[271] & b[166])^(a[270] & b[167])^(a[269] & b[168])^(a[268] & b[169])^(a[267] & b[170])^(a[266] & b[171])^(a[265] & b[172])^(a[264] & b[173])^(a[263] & b[174])^(a[262] & b[175])^(a[261] & b[176])^(a[260] & b[177])^(a[259] & b[178])^(a[258] & b[179])^(a[257] & b[180])^(a[256] & b[181])^(a[255] & b[182])^(a[254] & b[183])^(a[253] & b[184])^(a[252] & b[185])^(a[251] & b[186])^(a[250] & b[187])^(a[249] & b[188])^(a[248] & b[189])^(a[247] & b[190])^(a[246] & b[191])^(a[245] & b[192])^(a[244] & b[193])^(a[243] & b[194])^(a[242] & b[195])^(a[241] & b[196])^(a[240] & b[197])^(a[239] & b[198])^(a[238] & b[199])^(a[237] & b[200])^(a[236] & b[201])^(a[235] & b[202])^(a[234] & b[203])^(a[233] & b[204])^(a[232] & b[205])^(a[231] & b[206])^(a[230] & b[207])^(a[229] & b[208])^(a[228] & b[209])^(a[227] & b[210])^(a[226] & b[211])^(a[225] & b[212])^(a[224] & b[213])^(a[223] & b[214])^(a[222] & b[215])^(a[221] & b[216])^(a[220] & b[217])^(a[219] & b[218])^(a[218] & b[219])^(a[217] & b[220])^(a[216] & b[221])^(a[215] & b[222])^(a[214] & b[223])^(a[213] & b[224])^(a[212] & b[225])^(a[211] & b[226])^(a[210] & b[227])^(a[209] & b[228])^(a[208] & b[229])^(a[207] & b[230])^(a[206] & b[231])^(a[205] & b[232])^(a[204] & b[233])^(a[203] & b[234])^(a[202] & b[235])^(a[201] & b[236])^(a[200] & b[237])^(a[199] & b[238])^(a[198] & b[239])^(a[197] & b[240])^(a[196] & b[241])^(a[195] & b[242])^(a[194] & b[243])^(a[193] & b[244])^(a[192] & b[245])^(a[191] & b[246])^(a[190] & b[247])^(a[189] & b[248])^(a[188] & b[249])^(a[187] & b[250])^(a[186] & b[251])^(a[185] & b[252])^(a[184] & b[253])^(a[183] & b[254])^(a[182] & b[255])^(a[181] & b[256])^(a[180] & b[257])^(a[179] & b[258])^(a[178] & b[259])^(a[177] & b[260])^(a[176] & b[261])^(a[175] & b[262])^(a[174] & b[263])^(a[173] & b[264])^(a[172] & b[265])^(a[171] & b[266])^(a[170] & b[267])^(a[169] & b[268])^(a[168] & b[269])^(a[167] & b[270])^(a[166] & b[271])^(a[165] & b[272])^(a[164] & b[273])^(a[163] & b[274])^(a[162] & b[275])^(a[161] & b[276])^(a[160] & b[277])^(a[159] & b[278])^(a[158] & b[279])^(a[157] & b[280])^(a[156] & b[281])^(a[155] & b[282])^(a[154] & b[283])^(a[153] & b[284])^(a[152] & b[285])^(a[151] & b[286])^(a[150] & b[287])^(a[149] & b[288])^(a[148] & b[289])^(a[147] & b[290])^(a[146] & b[291])^(a[145] & b[292])^(a[144] & b[293])^(a[143] & b[294])^(a[142] & b[295])^(a[141] & b[296])^(a[140] & b[297])^(a[139] & b[298])^(a[138] & b[299])^(a[137] & b[300])^(a[136] & b[301])^(a[135] & b[302])^(a[134] & b[303])^(a[133] & b[304])^(a[132] & b[305])^(a[131] & b[306])^(a[130] & b[307])^(a[129] & b[308])^(a[128] & b[309])^(a[127] & b[310])^(a[126] & b[311])^(a[125] & b[312])^(a[124] & b[313])^(a[123] & b[314])^(a[122] & b[315])^(a[121] & b[316])^(a[120] & b[317])^(a[119] & b[318])^(a[118] & b[319])^(a[117] & b[320])^(a[116] & b[321])^(a[115] & b[322])^(a[114] & b[323])^(a[113] & b[324])^(a[112] & b[325])^(a[111] & b[326])^(a[110] & b[327])^(a[109] & b[328])^(a[108] & b[329])^(a[107] & b[330])^(a[106] & b[331])^(a[105] & b[332])^(a[104] & b[333])^(a[103] & b[334])^(a[102] & b[335])^(a[101] & b[336])^(a[100] & b[337])^(a[99] & b[338])^(a[98] & b[339])^(a[97] & b[340])^(a[96] & b[341])^(a[95] & b[342])^(a[94] & b[343])^(a[93] & b[344])^(a[92] & b[345])^(a[91] & b[346])^(a[90] & b[347])^(a[89] & b[348])^(a[88] & b[349])^(a[87] & b[350])^(a[86] & b[351])^(a[85] & b[352])^(a[84] & b[353])^(a[83] & b[354])^(a[82] & b[355])^(a[81] & b[356])^(a[80] & b[357])^(a[79] & b[358])^(a[78] & b[359])^(a[77] & b[360])^(a[76] & b[361])^(a[75] & b[362])^(a[74] & b[363])^(a[73] & b[364])^(a[72] & b[365])^(a[71] & b[366])^(a[70] & b[367])^(a[69] & b[368])^(a[68] & b[369])^(a[67] & b[370])^(a[66] & b[371])^(a[65] & b[372])^(a[64] & b[373])^(a[63] & b[374])^(a[62] & b[375])^(a[61] & b[376])^(a[60] & b[377])^(a[59] & b[378])^(a[58] & b[379])^(a[57] & b[380])^(a[56] & b[381])^(a[55] & b[382])^(a[54] & b[383])^(a[53] & b[384])^(a[52] & b[385])^(a[51] & b[386])^(a[50] & b[387])^(a[49] & b[388])^(a[48] & b[389])^(a[47] & b[390])^(a[46] & b[391])^(a[45] & b[392])^(a[44] & b[393])^(a[43] & b[394])^(a[42] & b[395])^(a[41] & b[396])^(a[40] & b[397])^(a[39] & b[398])^(a[38] & b[399])^(a[37] & b[400])^(a[36] & b[401])^(a[35] & b[402])^(a[34] & b[403])^(a[33] & b[404])^(a[32] & b[405])^(a[31] & b[406])^(a[30] & b[407])^(a[29] & b[408]);
assign y[438] = (a[408] & b[30])^(a[407] & b[31])^(a[406] & b[32])^(a[405] & b[33])^(a[404] & b[34])^(a[403] & b[35])^(a[402] & b[36])^(a[401] & b[37])^(a[400] & b[38])^(a[399] & b[39])^(a[398] & b[40])^(a[397] & b[41])^(a[396] & b[42])^(a[395] & b[43])^(a[394] & b[44])^(a[393] & b[45])^(a[392] & b[46])^(a[391] & b[47])^(a[390] & b[48])^(a[389] & b[49])^(a[388] & b[50])^(a[387] & b[51])^(a[386] & b[52])^(a[385] & b[53])^(a[384] & b[54])^(a[383] & b[55])^(a[382] & b[56])^(a[381] & b[57])^(a[380] & b[58])^(a[379] & b[59])^(a[378] & b[60])^(a[377] & b[61])^(a[376] & b[62])^(a[375] & b[63])^(a[374] & b[64])^(a[373] & b[65])^(a[372] & b[66])^(a[371] & b[67])^(a[370] & b[68])^(a[369] & b[69])^(a[368] & b[70])^(a[367] & b[71])^(a[366] & b[72])^(a[365] & b[73])^(a[364] & b[74])^(a[363] & b[75])^(a[362] & b[76])^(a[361] & b[77])^(a[360] & b[78])^(a[359] & b[79])^(a[358] & b[80])^(a[357] & b[81])^(a[356] & b[82])^(a[355] & b[83])^(a[354] & b[84])^(a[353] & b[85])^(a[352] & b[86])^(a[351] & b[87])^(a[350] & b[88])^(a[349] & b[89])^(a[348] & b[90])^(a[347] & b[91])^(a[346] & b[92])^(a[345] & b[93])^(a[344] & b[94])^(a[343] & b[95])^(a[342] & b[96])^(a[341] & b[97])^(a[340] & b[98])^(a[339] & b[99])^(a[338] & b[100])^(a[337] & b[101])^(a[336] & b[102])^(a[335] & b[103])^(a[334] & b[104])^(a[333] & b[105])^(a[332] & b[106])^(a[331] & b[107])^(a[330] & b[108])^(a[329] & b[109])^(a[328] & b[110])^(a[327] & b[111])^(a[326] & b[112])^(a[325] & b[113])^(a[324] & b[114])^(a[323] & b[115])^(a[322] & b[116])^(a[321] & b[117])^(a[320] & b[118])^(a[319] & b[119])^(a[318] & b[120])^(a[317] & b[121])^(a[316] & b[122])^(a[315] & b[123])^(a[314] & b[124])^(a[313] & b[125])^(a[312] & b[126])^(a[311] & b[127])^(a[310] & b[128])^(a[309] & b[129])^(a[308] & b[130])^(a[307] & b[131])^(a[306] & b[132])^(a[305] & b[133])^(a[304] & b[134])^(a[303] & b[135])^(a[302] & b[136])^(a[301] & b[137])^(a[300] & b[138])^(a[299] & b[139])^(a[298] & b[140])^(a[297] & b[141])^(a[296] & b[142])^(a[295] & b[143])^(a[294] & b[144])^(a[293] & b[145])^(a[292] & b[146])^(a[291] & b[147])^(a[290] & b[148])^(a[289] & b[149])^(a[288] & b[150])^(a[287] & b[151])^(a[286] & b[152])^(a[285] & b[153])^(a[284] & b[154])^(a[283] & b[155])^(a[282] & b[156])^(a[281] & b[157])^(a[280] & b[158])^(a[279] & b[159])^(a[278] & b[160])^(a[277] & b[161])^(a[276] & b[162])^(a[275] & b[163])^(a[274] & b[164])^(a[273] & b[165])^(a[272] & b[166])^(a[271] & b[167])^(a[270] & b[168])^(a[269] & b[169])^(a[268] & b[170])^(a[267] & b[171])^(a[266] & b[172])^(a[265] & b[173])^(a[264] & b[174])^(a[263] & b[175])^(a[262] & b[176])^(a[261] & b[177])^(a[260] & b[178])^(a[259] & b[179])^(a[258] & b[180])^(a[257] & b[181])^(a[256] & b[182])^(a[255] & b[183])^(a[254] & b[184])^(a[253] & b[185])^(a[252] & b[186])^(a[251] & b[187])^(a[250] & b[188])^(a[249] & b[189])^(a[248] & b[190])^(a[247] & b[191])^(a[246] & b[192])^(a[245] & b[193])^(a[244] & b[194])^(a[243] & b[195])^(a[242] & b[196])^(a[241] & b[197])^(a[240] & b[198])^(a[239] & b[199])^(a[238] & b[200])^(a[237] & b[201])^(a[236] & b[202])^(a[235] & b[203])^(a[234] & b[204])^(a[233] & b[205])^(a[232] & b[206])^(a[231] & b[207])^(a[230] & b[208])^(a[229] & b[209])^(a[228] & b[210])^(a[227] & b[211])^(a[226] & b[212])^(a[225] & b[213])^(a[224] & b[214])^(a[223] & b[215])^(a[222] & b[216])^(a[221] & b[217])^(a[220] & b[218])^(a[219] & b[219])^(a[218] & b[220])^(a[217] & b[221])^(a[216] & b[222])^(a[215] & b[223])^(a[214] & b[224])^(a[213] & b[225])^(a[212] & b[226])^(a[211] & b[227])^(a[210] & b[228])^(a[209] & b[229])^(a[208] & b[230])^(a[207] & b[231])^(a[206] & b[232])^(a[205] & b[233])^(a[204] & b[234])^(a[203] & b[235])^(a[202] & b[236])^(a[201] & b[237])^(a[200] & b[238])^(a[199] & b[239])^(a[198] & b[240])^(a[197] & b[241])^(a[196] & b[242])^(a[195] & b[243])^(a[194] & b[244])^(a[193] & b[245])^(a[192] & b[246])^(a[191] & b[247])^(a[190] & b[248])^(a[189] & b[249])^(a[188] & b[250])^(a[187] & b[251])^(a[186] & b[252])^(a[185] & b[253])^(a[184] & b[254])^(a[183] & b[255])^(a[182] & b[256])^(a[181] & b[257])^(a[180] & b[258])^(a[179] & b[259])^(a[178] & b[260])^(a[177] & b[261])^(a[176] & b[262])^(a[175] & b[263])^(a[174] & b[264])^(a[173] & b[265])^(a[172] & b[266])^(a[171] & b[267])^(a[170] & b[268])^(a[169] & b[269])^(a[168] & b[270])^(a[167] & b[271])^(a[166] & b[272])^(a[165] & b[273])^(a[164] & b[274])^(a[163] & b[275])^(a[162] & b[276])^(a[161] & b[277])^(a[160] & b[278])^(a[159] & b[279])^(a[158] & b[280])^(a[157] & b[281])^(a[156] & b[282])^(a[155] & b[283])^(a[154] & b[284])^(a[153] & b[285])^(a[152] & b[286])^(a[151] & b[287])^(a[150] & b[288])^(a[149] & b[289])^(a[148] & b[290])^(a[147] & b[291])^(a[146] & b[292])^(a[145] & b[293])^(a[144] & b[294])^(a[143] & b[295])^(a[142] & b[296])^(a[141] & b[297])^(a[140] & b[298])^(a[139] & b[299])^(a[138] & b[300])^(a[137] & b[301])^(a[136] & b[302])^(a[135] & b[303])^(a[134] & b[304])^(a[133] & b[305])^(a[132] & b[306])^(a[131] & b[307])^(a[130] & b[308])^(a[129] & b[309])^(a[128] & b[310])^(a[127] & b[311])^(a[126] & b[312])^(a[125] & b[313])^(a[124] & b[314])^(a[123] & b[315])^(a[122] & b[316])^(a[121] & b[317])^(a[120] & b[318])^(a[119] & b[319])^(a[118] & b[320])^(a[117] & b[321])^(a[116] & b[322])^(a[115] & b[323])^(a[114] & b[324])^(a[113] & b[325])^(a[112] & b[326])^(a[111] & b[327])^(a[110] & b[328])^(a[109] & b[329])^(a[108] & b[330])^(a[107] & b[331])^(a[106] & b[332])^(a[105] & b[333])^(a[104] & b[334])^(a[103] & b[335])^(a[102] & b[336])^(a[101] & b[337])^(a[100] & b[338])^(a[99] & b[339])^(a[98] & b[340])^(a[97] & b[341])^(a[96] & b[342])^(a[95] & b[343])^(a[94] & b[344])^(a[93] & b[345])^(a[92] & b[346])^(a[91] & b[347])^(a[90] & b[348])^(a[89] & b[349])^(a[88] & b[350])^(a[87] & b[351])^(a[86] & b[352])^(a[85] & b[353])^(a[84] & b[354])^(a[83] & b[355])^(a[82] & b[356])^(a[81] & b[357])^(a[80] & b[358])^(a[79] & b[359])^(a[78] & b[360])^(a[77] & b[361])^(a[76] & b[362])^(a[75] & b[363])^(a[74] & b[364])^(a[73] & b[365])^(a[72] & b[366])^(a[71] & b[367])^(a[70] & b[368])^(a[69] & b[369])^(a[68] & b[370])^(a[67] & b[371])^(a[66] & b[372])^(a[65] & b[373])^(a[64] & b[374])^(a[63] & b[375])^(a[62] & b[376])^(a[61] & b[377])^(a[60] & b[378])^(a[59] & b[379])^(a[58] & b[380])^(a[57] & b[381])^(a[56] & b[382])^(a[55] & b[383])^(a[54] & b[384])^(a[53] & b[385])^(a[52] & b[386])^(a[51] & b[387])^(a[50] & b[388])^(a[49] & b[389])^(a[48] & b[390])^(a[47] & b[391])^(a[46] & b[392])^(a[45] & b[393])^(a[44] & b[394])^(a[43] & b[395])^(a[42] & b[396])^(a[41] & b[397])^(a[40] & b[398])^(a[39] & b[399])^(a[38] & b[400])^(a[37] & b[401])^(a[36] & b[402])^(a[35] & b[403])^(a[34] & b[404])^(a[33] & b[405])^(a[32] & b[406])^(a[31] & b[407])^(a[30] & b[408]);
assign y[439] = (a[408] & b[31])^(a[407] & b[32])^(a[406] & b[33])^(a[405] & b[34])^(a[404] & b[35])^(a[403] & b[36])^(a[402] & b[37])^(a[401] & b[38])^(a[400] & b[39])^(a[399] & b[40])^(a[398] & b[41])^(a[397] & b[42])^(a[396] & b[43])^(a[395] & b[44])^(a[394] & b[45])^(a[393] & b[46])^(a[392] & b[47])^(a[391] & b[48])^(a[390] & b[49])^(a[389] & b[50])^(a[388] & b[51])^(a[387] & b[52])^(a[386] & b[53])^(a[385] & b[54])^(a[384] & b[55])^(a[383] & b[56])^(a[382] & b[57])^(a[381] & b[58])^(a[380] & b[59])^(a[379] & b[60])^(a[378] & b[61])^(a[377] & b[62])^(a[376] & b[63])^(a[375] & b[64])^(a[374] & b[65])^(a[373] & b[66])^(a[372] & b[67])^(a[371] & b[68])^(a[370] & b[69])^(a[369] & b[70])^(a[368] & b[71])^(a[367] & b[72])^(a[366] & b[73])^(a[365] & b[74])^(a[364] & b[75])^(a[363] & b[76])^(a[362] & b[77])^(a[361] & b[78])^(a[360] & b[79])^(a[359] & b[80])^(a[358] & b[81])^(a[357] & b[82])^(a[356] & b[83])^(a[355] & b[84])^(a[354] & b[85])^(a[353] & b[86])^(a[352] & b[87])^(a[351] & b[88])^(a[350] & b[89])^(a[349] & b[90])^(a[348] & b[91])^(a[347] & b[92])^(a[346] & b[93])^(a[345] & b[94])^(a[344] & b[95])^(a[343] & b[96])^(a[342] & b[97])^(a[341] & b[98])^(a[340] & b[99])^(a[339] & b[100])^(a[338] & b[101])^(a[337] & b[102])^(a[336] & b[103])^(a[335] & b[104])^(a[334] & b[105])^(a[333] & b[106])^(a[332] & b[107])^(a[331] & b[108])^(a[330] & b[109])^(a[329] & b[110])^(a[328] & b[111])^(a[327] & b[112])^(a[326] & b[113])^(a[325] & b[114])^(a[324] & b[115])^(a[323] & b[116])^(a[322] & b[117])^(a[321] & b[118])^(a[320] & b[119])^(a[319] & b[120])^(a[318] & b[121])^(a[317] & b[122])^(a[316] & b[123])^(a[315] & b[124])^(a[314] & b[125])^(a[313] & b[126])^(a[312] & b[127])^(a[311] & b[128])^(a[310] & b[129])^(a[309] & b[130])^(a[308] & b[131])^(a[307] & b[132])^(a[306] & b[133])^(a[305] & b[134])^(a[304] & b[135])^(a[303] & b[136])^(a[302] & b[137])^(a[301] & b[138])^(a[300] & b[139])^(a[299] & b[140])^(a[298] & b[141])^(a[297] & b[142])^(a[296] & b[143])^(a[295] & b[144])^(a[294] & b[145])^(a[293] & b[146])^(a[292] & b[147])^(a[291] & b[148])^(a[290] & b[149])^(a[289] & b[150])^(a[288] & b[151])^(a[287] & b[152])^(a[286] & b[153])^(a[285] & b[154])^(a[284] & b[155])^(a[283] & b[156])^(a[282] & b[157])^(a[281] & b[158])^(a[280] & b[159])^(a[279] & b[160])^(a[278] & b[161])^(a[277] & b[162])^(a[276] & b[163])^(a[275] & b[164])^(a[274] & b[165])^(a[273] & b[166])^(a[272] & b[167])^(a[271] & b[168])^(a[270] & b[169])^(a[269] & b[170])^(a[268] & b[171])^(a[267] & b[172])^(a[266] & b[173])^(a[265] & b[174])^(a[264] & b[175])^(a[263] & b[176])^(a[262] & b[177])^(a[261] & b[178])^(a[260] & b[179])^(a[259] & b[180])^(a[258] & b[181])^(a[257] & b[182])^(a[256] & b[183])^(a[255] & b[184])^(a[254] & b[185])^(a[253] & b[186])^(a[252] & b[187])^(a[251] & b[188])^(a[250] & b[189])^(a[249] & b[190])^(a[248] & b[191])^(a[247] & b[192])^(a[246] & b[193])^(a[245] & b[194])^(a[244] & b[195])^(a[243] & b[196])^(a[242] & b[197])^(a[241] & b[198])^(a[240] & b[199])^(a[239] & b[200])^(a[238] & b[201])^(a[237] & b[202])^(a[236] & b[203])^(a[235] & b[204])^(a[234] & b[205])^(a[233] & b[206])^(a[232] & b[207])^(a[231] & b[208])^(a[230] & b[209])^(a[229] & b[210])^(a[228] & b[211])^(a[227] & b[212])^(a[226] & b[213])^(a[225] & b[214])^(a[224] & b[215])^(a[223] & b[216])^(a[222] & b[217])^(a[221] & b[218])^(a[220] & b[219])^(a[219] & b[220])^(a[218] & b[221])^(a[217] & b[222])^(a[216] & b[223])^(a[215] & b[224])^(a[214] & b[225])^(a[213] & b[226])^(a[212] & b[227])^(a[211] & b[228])^(a[210] & b[229])^(a[209] & b[230])^(a[208] & b[231])^(a[207] & b[232])^(a[206] & b[233])^(a[205] & b[234])^(a[204] & b[235])^(a[203] & b[236])^(a[202] & b[237])^(a[201] & b[238])^(a[200] & b[239])^(a[199] & b[240])^(a[198] & b[241])^(a[197] & b[242])^(a[196] & b[243])^(a[195] & b[244])^(a[194] & b[245])^(a[193] & b[246])^(a[192] & b[247])^(a[191] & b[248])^(a[190] & b[249])^(a[189] & b[250])^(a[188] & b[251])^(a[187] & b[252])^(a[186] & b[253])^(a[185] & b[254])^(a[184] & b[255])^(a[183] & b[256])^(a[182] & b[257])^(a[181] & b[258])^(a[180] & b[259])^(a[179] & b[260])^(a[178] & b[261])^(a[177] & b[262])^(a[176] & b[263])^(a[175] & b[264])^(a[174] & b[265])^(a[173] & b[266])^(a[172] & b[267])^(a[171] & b[268])^(a[170] & b[269])^(a[169] & b[270])^(a[168] & b[271])^(a[167] & b[272])^(a[166] & b[273])^(a[165] & b[274])^(a[164] & b[275])^(a[163] & b[276])^(a[162] & b[277])^(a[161] & b[278])^(a[160] & b[279])^(a[159] & b[280])^(a[158] & b[281])^(a[157] & b[282])^(a[156] & b[283])^(a[155] & b[284])^(a[154] & b[285])^(a[153] & b[286])^(a[152] & b[287])^(a[151] & b[288])^(a[150] & b[289])^(a[149] & b[290])^(a[148] & b[291])^(a[147] & b[292])^(a[146] & b[293])^(a[145] & b[294])^(a[144] & b[295])^(a[143] & b[296])^(a[142] & b[297])^(a[141] & b[298])^(a[140] & b[299])^(a[139] & b[300])^(a[138] & b[301])^(a[137] & b[302])^(a[136] & b[303])^(a[135] & b[304])^(a[134] & b[305])^(a[133] & b[306])^(a[132] & b[307])^(a[131] & b[308])^(a[130] & b[309])^(a[129] & b[310])^(a[128] & b[311])^(a[127] & b[312])^(a[126] & b[313])^(a[125] & b[314])^(a[124] & b[315])^(a[123] & b[316])^(a[122] & b[317])^(a[121] & b[318])^(a[120] & b[319])^(a[119] & b[320])^(a[118] & b[321])^(a[117] & b[322])^(a[116] & b[323])^(a[115] & b[324])^(a[114] & b[325])^(a[113] & b[326])^(a[112] & b[327])^(a[111] & b[328])^(a[110] & b[329])^(a[109] & b[330])^(a[108] & b[331])^(a[107] & b[332])^(a[106] & b[333])^(a[105] & b[334])^(a[104] & b[335])^(a[103] & b[336])^(a[102] & b[337])^(a[101] & b[338])^(a[100] & b[339])^(a[99] & b[340])^(a[98] & b[341])^(a[97] & b[342])^(a[96] & b[343])^(a[95] & b[344])^(a[94] & b[345])^(a[93] & b[346])^(a[92] & b[347])^(a[91] & b[348])^(a[90] & b[349])^(a[89] & b[350])^(a[88] & b[351])^(a[87] & b[352])^(a[86] & b[353])^(a[85] & b[354])^(a[84] & b[355])^(a[83] & b[356])^(a[82] & b[357])^(a[81] & b[358])^(a[80] & b[359])^(a[79] & b[360])^(a[78] & b[361])^(a[77] & b[362])^(a[76] & b[363])^(a[75] & b[364])^(a[74] & b[365])^(a[73] & b[366])^(a[72] & b[367])^(a[71] & b[368])^(a[70] & b[369])^(a[69] & b[370])^(a[68] & b[371])^(a[67] & b[372])^(a[66] & b[373])^(a[65] & b[374])^(a[64] & b[375])^(a[63] & b[376])^(a[62] & b[377])^(a[61] & b[378])^(a[60] & b[379])^(a[59] & b[380])^(a[58] & b[381])^(a[57] & b[382])^(a[56] & b[383])^(a[55] & b[384])^(a[54] & b[385])^(a[53] & b[386])^(a[52] & b[387])^(a[51] & b[388])^(a[50] & b[389])^(a[49] & b[390])^(a[48] & b[391])^(a[47] & b[392])^(a[46] & b[393])^(a[45] & b[394])^(a[44] & b[395])^(a[43] & b[396])^(a[42] & b[397])^(a[41] & b[398])^(a[40] & b[399])^(a[39] & b[400])^(a[38] & b[401])^(a[37] & b[402])^(a[36] & b[403])^(a[35] & b[404])^(a[34] & b[405])^(a[33] & b[406])^(a[32] & b[407])^(a[31] & b[408]);
assign y[440] = (a[408] & b[32])^(a[407] & b[33])^(a[406] & b[34])^(a[405] & b[35])^(a[404] & b[36])^(a[403] & b[37])^(a[402] & b[38])^(a[401] & b[39])^(a[400] & b[40])^(a[399] & b[41])^(a[398] & b[42])^(a[397] & b[43])^(a[396] & b[44])^(a[395] & b[45])^(a[394] & b[46])^(a[393] & b[47])^(a[392] & b[48])^(a[391] & b[49])^(a[390] & b[50])^(a[389] & b[51])^(a[388] & b[52])^(a[387] & b[53])^(a[386] & b[54])^(a[385] & b[55])^(a[384] & b[56])^(a[383] & b[57])^(a[382] & b[58])^(a[381] & b[59])^(a[380] & b[60])^(a[379] & b[61])^(a[378] & b[62])^(a[377] & b[63])^(a[376] & b[64])^(a[375] & b[65])^(a[374] & b[66])^(a[373] & b[67])^(a[372] & b[68])^(a[371] & b[69])^(a[370] & b[70])^(a[369] & b[71])^(a[368] & b[72])^(a[367] & b[73])^(a[366] & b[74])^(a[365] & b[75])^(a[364] & b[76])^(a[363] & b[77])^(a[362] & b[78])^(a[361] & b[79])^(a[360] & b[80])^(a[359] & b[81])^(a[358] & b[82])^(a[357] & b[83])^(a[356] & b[84])^(a[355] & b[85])^(a[354] & b[86])^(a[353] & b[87])^(a[352] & b[88])^(a[351] & b[89])^(a[350] & b[90])^(a[349] & b[91])^(a[348] & b[92])^(a[347] & b[93])^(a[346] & b[94])^(a[345] & b[95])^(a[344] & b[96])^(a[343] & b[97])^(a[342] & b[98])^(a[341] & b[99])^(a[340] & b[100])^(a[339] & b[101])^(a[338] & b[102])^(a[337] & b[103])^(a[336] & b[104])^(a[335] & b[105])^(a[334] & b[106])^(a[333] & b[107])^(a[332] & b[108])^(a[331] & b[109])^(a[330] & b[110])^(a[329] & b[111])^(a[328] & b[112])^(a[327] & b[113])^(a[326] & b[114])^(a[325] & b[115])^(a[324] & b[116])^(a[323] & b[117])^(a[322] & b[118])^(a[321] & b[119])^(a[320] & b[120])^(a[319] & b[121])^(a[318] & b[122])^(a[317] & b[123])^(a[316] & b[124])^(a[315] & b[125])^(a[314] & b[126])^(a[313] & b[127])^(a[312] & b[128])^(a[311] & b[129])^(a[310] & b[130])^(a[309] & b[131])^(a[308] & b[132])^(a[307] & b[133])^(a[306] & b[134])^(a[305] & b[135])^(a[304] & b[136])^(a[303] & b[137])^(a[302] & b[138])^(a[301] & b[139])^(a[300] & b[140])^(a[299] & b[141])^(a[298] & b[142])^(a[297] & b[143])^(a[296] & b[144])^(a[295] & b[145])^(a[294] & b[146])^(a[293] & b[147])^(a[292] & b[148])^(a[291] & b[149])^(a[290] & b[150])^(a[289] & b[151])^(a[288] & b[152])^(a[287] & b[153])^(a[286] & b[154])^(a[285] & b[155])^(a[284] & b[156])^(a[283] & b[157])^(a[282] & b[158])^(a[281] & b[159])^(a[280] & b[160])^(a[279] & b[161])^(a[278] & b[162])^(a[277] & b[163])^(a[276] & b[164])^(a[275] & b[165])^(a[274] & b[166])^(a[273] & b[167])^(a[272] & b[168])^(a[271] & b[169])^(a[270] & b[170])^(a[269] & b[171])^(a[268] & b[172])^(a[267] & b[173])^(a[266] & b[174])^(a[265] & b[175])^(a[264] & b[176])^(a[263] & b[177])^(a[262] & b[178])^(a[261] & b[179])^(a[260] & b[180])^(a[259] & b[181])^(a[258] & b[182])^(a[257] & b[183])^(a[256] & b[184])^(a[255] & b[185])^(a[254] & b[186])^(a[253] & b[187])^(a[252] & b[188])^(a[251] & b[189])^(a[250] & b[190])^(a[249] & b[191])^(a[248] & b[192])^(a[247] & b[193])^(a[246] & b[194])^(a[245] & b[195])^(a[244] & b[196])^(a[243] & b[197])^(a[242] & b[198])^(a[241] & b[199])^(a[240] & b[200])^(a[239] & b[201])^(a[238] & b[202])^(a[237] & b[203])^(a[236] & b[204])^(a[235] & b[205])^(a[234] & b[206])^(a[233] & b[207])^(a[232] & b[208])^(a[231] & b[209])^(a[230] & b[210])^(a[229] & b[211])^(a[228] & b[212])^(a[227] & b[213])^(a[226] & b[214])^(a[225] & b[215])^(a[224] & b[216])^(a[223] & b[217])^(a[222] & b[218])^(a[221] & b[219])^(a[220] & b[220])^(a[219] & b[221])^(a[218] & b[222])^(a[217] & b[223])^(a[216] & b[224])^(a[215] & b[225])^(a[214] & b[226])^(a[213] & b[227])^(a[212] & b[228])^(a[211] & b[229])^(a[210] & b[230])^(a[209] & b[231])^(a[208] & b[232])^(a[207] & b[233])^(a[206] & b[234])^(a[205] & b[235])^(a[204] & b[236])^(a[203] & b[237])^(a[202] & b[238])^(a[201] & b[239])^(a[200] & b[240])^(a[199] & b[241])^(a[198] & b[242])^(a[197] & b[243])^(a[196] & b[244])^(a[195] & b[245])^(a[194] & b[246])^(a[193] & b[247])^(a[192] & b[248])^(a[191] & b[249])^(a[190] & b[250])^(a[189] & b[251])^(a[188] & b[252])^(a[187] & b[253])^(a[186] & b[254])^(a[185] & b[255])^(a[184] & b[256])^(a[183] & b[257])^(a[182] & b[258])^(a[181] & b[259])^(a[180] & b[260])^(a[179] & b[261])^(a[178] & b[262])^(a[177] & b[263])^(a[176] & b[264])^(a[175] & b[265])^(a[174] & b[266])^(a[173] & b[267])^(a[172] & b[268])^(a[171] & b[269])^(a[170] & b[270])^(a[169] & b[271])^(a[168] & b[272])^(a[167] & b[273])^(a[166] & b[274])^(a[165] & b[275])^(a[164] & b[276])^(a[163] & b[277])^(a[162] & b[278])^(a[161] & b[279])^(a[160] & b[280])^(a[159] & b[281])^(a[158] & b[282])^(a[157] & b[283])^(a[156] & b[284])^(a[155] & b[285])^(a[154] & b[286])^(a[153] & b[287])^(a[152] & b[288])^(a[151] & b[289])^(a[150] & b[290])^(a[149] & b[291])^(a[148] & b[292])^(a[147] & b[293])^(a[146] & b[294])^(a[145] & b[295])^(a[144] & b[296])^(a[143] & b[297])^(a[142] & b[298])^(a[141] & b[299])^(a[140] & b[300])^(a[139] & b[301])^(a[138] & b[302])^(a[137] & b[303])^(a[136] & b[304])^(a[135] & b[305])^(a[134] & b[306])^(a[133] & b[307])^(a[132] & b[308])^(a[131] & b[309])^(a[130] & b[310])^(a[129] & b[311])^(a[128] & b[312])^(a[127] & b[313])^(a[126] & b[314])^(a[125] & b[315])^(a[124] & b[316])^(a[123] & b[317])^(a[122] & b[318])^(a[121] & b[319])^(a[120] & b[320])^(a[119] & b[321])^(a[118] & b[322])^(a[117] & b[323])^(a[116] & b[324])^(a[115] & b[325])^(a[114] & b[326])^(a[113] & b[327])^(a[112] & b[328])^(a[111] & b[329])^(a[110] & b[330])^(a[109] & b[331])^(a[108] & b[332])^(a[107] & b[333])^(a[106] & b[334])^(a[105] & b[335])^(a[104] & b[336])^(a[103] & b[337])^(a[102] & b[338])^(a[101] & b[339])^(a[100] & b[340])^(a[99] & b[341])^(a[98] & b[342])^(a[97] & b[343])^(a[96] & b[344])^(a[95] & b[345])^(a[94] & b[346])^(a[93] & b[347])^(a[92] & b[348])^(a[91] & b[349])^(a[90] & b[350])^(a[89] & b[351])^(a[88] & b[352])^(a[87] & b[353])^(a[86] & b[354])^(a[85] & b[355])^(a[84] & b[356])^(a[83] & b[357])^(a[82] & b[358])^(a[81] & b[359])^(a[80] & b[360])^(a[79] & b[361])^(a[78] & b[362])^(a[77] & b[363])^(a[76] & b[364])^(a[75] & b[365])^(a[74] & b[366])^(a[73] & b[367])^(a[72] & b[368])^(a[71] & b[369])^(a[70] & b[370])^(a[69] & b[371])^(a[68] & b[372])^(a[67] & b[373])^(a[66] & b[374])^(a[65] & b[375])^(a[64] & b[376])^(a[63] & b[377])^(a[62] & b[378])^(a[61] & b[379])^(a[60] & b[380])^(a[59] & b[381])^(a[58] & b[382])^(a[57] & b[383])^(a[56] & b[384])^(a[55] & b[385])^(a[54] & b[386])^(a[53] & b[387])^(a[52] & b[388])^(a[51] & b[389])^(a[50] & b[390])^(a[49] & b[391])^(a[48] & b[392])^(a[47] & b[393])^(a[46] & b[394])^(a[45] & b[395])^(a[44] & b[396])^(a[43] & b[397])^(a[42] & b[398])^(a[41] & b[399])^(a[40] & b[400])^(a[39] & b[401])^(a[38] & b[402])^(a[37] & b[403])^(a[36] & b[404])^(a[35] & b[405])^(a[34] & b[406])^(a[33] & b[407])^(a[32] & b[408]);
assign y[441] = (a[408] & b[33])^(a[407] & b[34])^(a[406] & b[35])^(a[405] & b[36])^(a[404] & b[37])^(a[403] & b[38])^(a[402] & b[39])^(a[401] & b[40])^(a[400] & b[41])^(a[399] & b[42])^(a[398] & b[43])^(a[397] & b[44])^(a[396] & b[45])^(a[395] & b[46])^(a[394] & b[47])^(a[393] & b[48])^(a[392] & b[49])^(a[391] & b[50])^(a[390] & b[51])^(a[389] & b[52])^(a[388] & b[53])^(a[387] & b[54])^(a[386] & b[55])^(a[385] & b[56])^(a[384] & b[57])^(a[383] & b[58])^(a[382] & b[59])^(a[381] & b[60])^(a[380] & b[61])^(a[379] & b[62])^(a[378] & b[63])^(a[377] & b[64])^(a[376] & b[65])^(a[375] & b[66])^(a[374] & b[67])^(a[373] & b[68])^(a[372] & b[69])^(a[371] & b[70])^(a[370] & b[71])^(a[369] & b[72])^(a[368] & b[73])^(a[367] & b[74])^(a[366] & b[75])^(a[365] & b[76])^(a[364] & b[77])^(a[363] & b[78])^(a[362] & b[79])^(a[361] & b[80])^(a[360] & b[81])^(a[359] & b[82])^(a[358] & b[83])^(a[357] & b[84])^(a[356] & b[85])^(a[355] & b[86])^(a[354] & b[87])^(a[353] & b[88])^(a[352] & b[89])^(a[351] & b[90])^(a[350] & b[91])^(a[349] & b[92])^(a[348] & b[93])^(a[347] & b[94])^(a[346] & b[95])^(a[345] & b[96])^(a[344] & b[97])^(a[343] & b[98])^(a[342] & b[99])^(a[341] & b[100])^(a[340] & b[101])^(a[339] & b[102])^(a[338] & b[103])^(a[337] & b[104])^(a[336] & b[105])^(a[335] & b[106])^(a[334] & b[107])^(a[333] & b[108])^(a[332] & b[109])^(a[331] & b[110])^(a[330] & b[111])^(a[329] & b[112])^(a[328] & b[113])^(a[327] & b[114])^(a[326] & b[115])^(a[325] & b[116])^(a[324] & b[117])^(a[323] & b[118])^(a[322] & b[119])^(a[321] & b[120])^(a[320] & b[121])^(a[319] & b[122])^(a[318] & b[123])^(a[317] & b[124])^(a[316] & b[125])^(a[315] & b[126])^(a[314] & b[127])^(a[313] & b[128])^(a[312] & b[129])^(a[311] & b[130])^(a[310] & b[131])^(a[309] & b[132])^(a[308] & b[133])^(a[307] & b[134])^(a[306] & b[135])^(a[305] & b[136])^(a[304] & b[137])^(a[303] & b[138])^(a[302] & b[139])^(a[301] & b[140])^(a[300] & b[141])^(a[299] & b[142])^(a[298] & b[143])^(a[297] & b[144])^(a[296] & b[145])^(a[295] & b[146])^(a[294] & b[147])^(a[293] & b[148])^(a[292] & b[149])^(a[291] & b[150])^(a[290] & b[151])^(a[289] & b[152])^(a[288] & b[153])^(a[287] & b[154])^(a[286] & b[155])^(a[285] & b[156])^(a[284] & b[157])^(a[283] & b[158])^(a[282] & b[159])^(a[281] & b[160])^(a[280] & b[161])^(a[279] & b[162])^(a[278] & b[163])^(a[277] & b[164])^(a[276] & b[165])^(a[275] & b[166])^(a[274] & b[167])^(a[273] & b[168])^(a[272] & b[169])^(a[271] & b[170])^(a[270] & b[171])^(a[269] & b[172])^(a[268] & b[173])^(a[267] & b[174])^(a[266] & b[175])^(a[265] & b[176])^(a[264] & b[177])^(a[263] & b[178])^(a[262] & b[179])^(a[261] & b[180])^(a[260] & b[181])^(a[259] & b[182])^(a[258] & b[183])^(a[257] & b[184])^(a[256] & b[185])^(a[255] & b[186])^(a[254] & b[187])^(a[253] & b[188])^(a[252] & b[189])^(a[251] & b[190])^(a[250] & b[191])^(a[249] & b[192])^(a[248] & b[193])^(a[247] & b[194])^(a[246] & b[195])^(a[245] & b[196])^(a[244] & b[197])^(a[243] & b[198])^(a[242] & b[199])^(a[241] & b[200])^(a[240] & b[201])^(a[239] & b[202])^(a[238] & b[203])^(a[237] & b[204])^(a[236] & b[205])^(a[235] & b[206])^(a[234] & b[207])^(a[233] & b[208])^(a[232] & b[209])^(a[231] & b[210])^(a[230] & b[211])^(a[229] & b[212])^(a[228] & b[213])^(a[227] & b[214])^(a[226] & b[215])^(a[225] & b[216])^(a[224] & b[217])^(a[223] & b[218])^(a[222] & b[219])^(a[221] & b[220])^(a[220] & b[221])^(a[219] & b[222])^(a[218] & b[223])^(a[217] & b[224])^(a[216] & b[225])^(a[215] & b[226])^(a[214] & b[227])^(a[213] & b[228])^(a[212] & b[229])^(a[211] & b[230])^(a[210] & b[231])^(a[209] & b[232])^(a[208] & b[233])^(a[207] & b[234])^(a[206] & b[235])^(a[205] & b[236])^(a[204] & b[237])^(a[203] & b[238])^(a[202] & b[239])^(a[201] & b[240])^(a[200] & b[241])^(a[199] & b[242])^(a[198] & b[243])^(a[197] & b[244])^(a[196] & b[245])^(a[195] & b[246])^(a[194] & b[247])^(a[193] & b[248])^(a[192] & b[249])^(a[191] & b[250])^(a[190] & b[251])^(a[189] & b[252])^(a[188] & b[253])^(a[187] & b[254])^(a[186] & b[255])^(a[185] & b[256])^(a[184] & b[257])^(a[183] & b[258])^(a[182] & b[259])^(a[181] & b[260])^(a[180] & b[261])^(a[179] & b[262])^(a[178] & b[263])^(a[177] & b[264])^(a[176] & b[265])^(a[175] & b[266])^(a[174] & b[267])^(a[173] & b[268])^(a[172] & b[269])^(a[171] & b[270])^(a[170] & b[271])^(a[169] & b[272])^(a[168] & b[273])^(a[167] & b[274])^(a[166] & b[275])^(a[165] & b[276])^(a[164] & b[277])^(a[163] & b[278])^(a[162] & b[279])^(a[161] & b[280])^(a[160] & b[281])^(a[159] & b[282])^(a[158] & b[283])^(a[157] & b[284])^(a[156] & b[285])^(a[155] & b[286])^(a[154] & b[287])^(a[153] & b[288])^(a[152] & b[289])^(a[151] & b[290])^(a[150] & b[291])^(a[149] & b[292])^(a[148] & b[293])^(a[147] & b[294])^(a[146] & b[295])^(a[145] & b[296])^(a[144] & b[297])^(a[143] & b[298])^(a[142] & b[299])^(a[141] & b[300])^(a[140] & b[301])^(a[139] & b[302])^(a[138] & b[303])^(a[137] & b[304])^(a[136] & b[305])^(a[135] & b[306])^(a[134] & b[307])^(a[133] & b[308])^(a[132] & b[309])^(a[131] & b[310])^(a[130] & b[311])^(a[129] & b[312])^(a[128] & b[313])^(a[127] & b[314])^(a[126] & b[315])^(a[125] & b[316])^(a[124] & b[317])^(a[123] & b[318])^(a[122] & b[319])^(a[121] & b[320])^(a[120] & b[321])^(a[119] & b[322])^(a[118] & b[323])^(a[117] & b[324])^(a[116] & b[325])^(a[115] & b[326])^(a[114] & b[327])^(a[113] & b[328])^(a[112] & b[329])^(a[111] & b[330])^(a[110] & b[331])^(a[109] & b[332])^(a[108] & b[333])^(a[107] & b[334])^(a[106] & b[335])^(a[105] & b[336])^(a[104] & b[337])^(a[103] & b[338])^(a[102] & b[339])^(a[101] & b[340])^(a[100] & b[341])^(a[99] & b[342])^(a[98] & b[343])^(a[97] & b[344])^(a[96] & b[345])^(a[95] & b[346])^(a[94] & b[347])^(a[93] & b[348])^(a[92] & b[349])^(a[91] & b[350])^(a[90] & b[351])^(a[89] & b[352])^(a[88] & b[353])^(a[87] & b[354])^(a[86] & b[355])^(a[85] & b[356])^(a[84] & b[357])^(a[83] & b[358])^(a[82] & b[359])^(a[81] & b[360])^(a[80] & b[361])^(a[79] & b[362])^(a[78] & b[363])^(a[77] & b[364])^(a[76] & b[365])^(a[75] & b[366])^(a[74] & b[367])^(a[73] & b[368])^(a[72] & b[369])^(a[71] & b[370])^(a[70] & b[371])^(a[69] & b[372])^(a[68] & b[373])^(a[67] & b[374])^(a[66] & b[375])^(a[65] & b[376])^(a[64] & b[377])^(a[63] & b[378])^(a[62] & b[379])^(a[61] & b[380])^(a[60] & b[381])^(a[59] & b[382])^(a[58] & b[383])^(a[57] & b[384])^(a[56] & b[385])^(a[55] & b[386])^(a[54] & b[387])^(a[53] & b[388])^(a[52] & b[389])^(a[51] & b[390])^(a[50] & b[391])^(a[49] & b[392])^(a[48] & b[393])^(a[47] & b[394])^(a[46] & b[395])^(a[45] & b[396])^(a[44] & b[397])^(a[43] & b[398])^(a[42] & b[399])^(a[41] & b[400])^(a[40] & b[401])^(a[39] & b[402])^(a[38] & b[403])^(a[37] & b[404])^(a[36] & b[405])^(a[35] & b[406])^(a[34] & b[407])^(a[33] & b[408]);
assign y[442] = (a[408] & b[34])^(a[407] & b[35])^(a[406] & b[36])^(a[405] & b[37])^(a[404] & b[38])^(a[403] & b[39])^(a[402] & b[40])^(a[401] & b[41])^(a[400] & b[42])^(a[399] & b[43])^(a[398] & b[44])^(a[397] & b[45])^(a[396] & b[46])^(a[395] & b[47])^(a[394] & b[48])^(a[393] & b[49])^(a[392] & b[50])^(a[391] & b[51])^(a[390] & b[52])^(a[389] & b[53])^(a[388] & b[54])^(a[387] & b[55])^(a[386] & b[56])^(a[385] & b[57])^(a[384] & b[58])^(a[383] & b[59])^(a[382] & b[60])^(a[381] & b[61])^(a[380] & b[62])^(a[379] & b[63])^(a[378] & b[64])^(a[377] & b[65])^(a[376] & b[66])^(a[375] & b[67])^(a[374] & b[68])^(a[373] & b[69])^(a[372] & b[70])^(a[371] & b[71])^(a[370] & b[72])^(a[369] & b[73])^(a[368] & b[74])^(a[367] & b[75])^(a[366] & b[76])^(a[365] & b[77])^(a[364] & b[78])^(a[363] & b[79])^(a[362] & b[80])^(a[361] & b[81])^(a[360] & b[82])^(a[359] & b[83])^(a[358] & b[84])^(a[357] & b[85])^(a[356] & b[86])^(a[355] & b[87])^(a[354] & b[88])^(a[353] & b[89])^(a[352] & b[90])^(a[351] & b[91])^(a[350] & b[92])^(a[349] & b[93])^(a[348] & b[94])^(a[347] & b[95])^(a[346] & b[96])^(a[345] & b[97])^(a[344] & b[98])^(a[343] & b[99])^(a[342] & b[100])^(a[341] & b[101])^(a[340] & b[102])^(a[339] & b[103])^(a[338] & b[104])^(a[337] & b[105])^(a[336] & b[106])^(a[335] & b[107])^(a[334] & b[108])^(a[333] & b[109])^(a[332] & b[110])^(a[331] & b[111])^(a[330] & b[112])^(a[329] & b[113])^(a[328] & b[114])^(a[327] & b[115])^(a[326] & b[116])^(a[325] & b[117])^(a[324] & b[118])^(a[323] & b[119])^(a[322] & b[120])^(a[321] & b[121])^(a[320] & b[122])^(a[319] & b[123])^(a[318] & b[124])^(a[317] & b[125])^(a[316] & b[126])^(a[315] & b[127])^(a[314] & b[128])^(a[313] & b[129])^(a[312] & b[130])^(a[311] & b[131])^(a[310] & b[132])^(a[309] & b[133])^(a[308] & b[134])^(a[307] & b[135])^(a[306] & b[136])^(a[305] & b[137])^(a[304] & b[138])^(a[303] & b[139])^(a[302] & b[140])^(a[301] & b[141])^(a[300] & b[142])^(a[299] & b[143])^(a[298] & b[144])^(a[297] & b[145])^(a[296] & b[146])^(a[295] & b[147])^(a[294] & b[148])^(a[293] & b[149])^(a[292] & b[150])^(a[291] & b[151])^(a[290] & b[152])^(a[289] & b[153])^(a[288] & b[154])^(a[287] & b[155])^(a[286] & b[156])^(a[285] & b[157])^(a[284] & b[158])^(a[283] & b[159])^(a[282] & b[160])^(a[281] & b[161])^(a[280] & b[162])^(a[279] & b[163])^(a[278] & b[164])^(a[277] & b[165])^(a[276] & b[166])^(a[275] & b[167])^(a[274] & b[168])^(a[273] & b[169])^(a[272] & b[170])^(a[271] & b[171])^(a[270] & b[172])^(a[269] & b[173])^(a[268] & b[174])^(a[267] & b[175])^(a[266] & b[176])^(a[265] & b[177])^(a[264] & b[178])^(a[263] & b[179])^(a[262] & b[180])^(a[261] & b[181])^(a[260] & b[182])^(a[259] & b[183])^(a[258] & b[184])^(a[257] & b[185])^(a[256] & b[186])^(a[255] & b[187])^(a[254] & b[188])^(a[253] & b[189])^(a[252] & b[190])^(a[251] & b[191])^(a[250] & b[192])^(a[249] & b[193])^(a[248] & b[194])^(a[247] & b[195])^(a[246] & b[196])^(a[245] & b[197])^(a[244] & b[198])^(a[243] & b[199])^(a[242] & b[200])^(a[241] & b[201])^(a[240] & b[202])^(a[239] & b[203])^(a[238] & b[204])^(a[237] & b[205])^(a[236] & b[206])^(a[235] & b[207])^(a[234] & b[208])^(a[233] & b[209])^(a[232] & b[210])^(a[231] & b[211])^(a[230] & b[212])^(a[229] & b[213])^(a[228] & b[214])^(a[227] & b[215])^(a[226] & b[216])^(a[225] & b[217])^(a[224] & b[218])^(a[223] & b[219])^(a[222] & b[220])^(a[221] & b[221])^(a[220] & b[222])^(a[219] & b[223])^(a[218] & b[224])^(a[217] & b[225])^(a[216] & b[226])^(a[215] & b[227])^(a[214] & b[228])^(a[213] & b[229])^(a[212] & b[230])^(a[211] & b[231])^(a[210] & b[232])^(a[209] & b[233])^(a[208] & b[234])^(a[207] & b[235])^(a[206] & b[236])^(a[205] & b[237])^(a[204] & b[238])^(a[203] & b[239])^(a[202] & b[240])^(a[201] & b[241])^(a[200] & b[242])^(a[199] & b[243])^(a[198] & b[244])^(a[197] & b[245])^(a[196] & b[246])^(a[195] & b[247])^(a[194] & b[248])^(a[193] & b[249])^(a[192] & b[250])^(a[191] & b[251])^(a[190] & b[252])^(a[189] & b[253])^(a[188] & b[254])^(a[187] & b[255])^(a[186] & b[256])^(a[185] & b[257])^(a[184] & b[258])^(a[183] & b[259])^(a[182] & b[260])^(a[181] & b[261])^(a[180] & b[262])^(a[179] & b[263])^(a[178] & b[264])^(a[177] & b[265])^(a[176] & b[266])^(a[175] & b[267])^(a[174] & b[268])^(a[173] & b[269])^(a[172] & b[270])^(a[171] & b[271])^(a[170] & b[272])^(a[169] & b[273])^(a[168] & b[274])^(a[167] & b[275])^(a[166] & b[276])^(a[165] & b[277])^(a[164] & b[278])^(a[163] & b[279])^(a[162] & b[280])^(a[161] & b[281])^(a[160] & b[282])^(a[159] & b[283])^(a[158] & b[284])^(a[157] & b[285])^(a[156] & b[286])^(a[155] & b[287])^(a[154] & b[288])^(a[153] & b[289])^(a[152] & b[290])^(a[151] & b[291])^(a[150] & b[292])^(a[149] & b[293])^(a[148] & b[294])^(a[147] & b[295])^(a[146] & b[296])^(a[145] & b[297])^(a[144] & b[298])^(a[143] & b[299])^(a[142] & b[300])^(a[141] & b[301])^(a[140] & b[302])^(a[139] & b[303])^(a[138] & b[304])^(a[137] & b[305])^(a[136] & b[306])^(a[135] & b[307])^(a[134] & b[308])^(a[133] & b[309])^(a[132] & b[310])^(a[131] & b[311])^(a[130] & b[312])^(a[129] & b[313])^(a[128] & b[314])^(a[127] & b[315])^(a[126] & b[316])^(a[125] & b[317])^(a[124] & b[318])^(a[123] & b[319])^(a[122] & b[320])^(a[121] & b[321])^(a[120] & b[322])^(a[119] & b[323])^(a[118] & b[324])^(a[117] & b[325])^(a[116] & b[326])^(a[115] & b[327])^(a[114] & b[328])^(a[113] & b[329])^(a[112] & b[330])^(a[111] & b[331])^(a[110] & b[332])^(a[109] & b[333])^(a[108] & b[334])^(a[107] & b[335])^(a[106] & b[336])^(a[105] & b[337])^(a[104] & b[338])^(a[103] & b[339])^(a[102] & b[340])^(a[101] & b[341])^(a[100] & b[342])^(a[99] & b[343])^(a[98] & b[344])^(a[97] & b[345])^(a[96] & b[346])^(a[95] & b[347])^(a[94] & b[348])^(a[93] & b[349])^(a[92] & b[350])^(a[91] & b[351])^(a[90] & b[352])^(a[89] & b[353])^(a[88] & b[354])^(a[87] & b[355])^(a[86] & b[356])^(a[85] & b[357])^(a[84] & b[358])^(a[83] & b[359])^(a[82] & b[360])^(a[81] & b[361])^(a[80] & b[362])^(a[79] & b[363])^(a[78] & b[364])^(a[77] & b[365])^(a[76] & b[366])^(a[75] & b[367])^(a[74] & b[368])^(a[73] & b[369])^(a[72] & b[370])^(a[71] & b[371])^(a[70] & b[372])^(a[69] & b[373])^(a[68] & b[374])^(a[67] & b[375])^(a[66] & b[376])^(a[65] & b[377])^(a[64] & b[378])^(a[63] & b[379])^(a[62] & b[380])^(a[61] & b[381])^(a[60] & b[382])^(a[59] & b[383])^(a[58] & b[384])^(a[57] & b[385])^(a[56] & b[386])^(a[55] & b[387])^(a[54] & b[388])^(a[53] & b[389])^(a[52] & b[390])^(a[51] & b[391])^(a[50] & b[392])^(a[49] & b[393])^(a[48] & b[394])^(a[47] & b[395])^(a[46] & b[396])^(a[45] & b[397])^(a[44] & b[398])^(a[43] & b[399])^(a[42] & b[400])^(a[41] & b[401])^(a[40] & b[402])^(a[39] & b[403])^(a[38] & b[404])^(a[37] & b[405])^(a[36] & b[406])^(a[35] & b[407])^(a[34] & b[408]);
assign y[443] = (a[408] & b[35])^(a[407] & b[36])^(a[406] & b[37])^(a[405] & b[38])^(a[404] & b[39])^(a[403] & b[40])^(a[402] & b[41])^(a[401] & b[42])^(a[400] & b[43])^(a[399] & b[44])^(a[398] & b[45])^(a[397] & b[46])^(a[396] & b[47])^(a[395] & b[48])^(a[394] & b[49])^(a[393] & b[50])^(a[392] & b[51])^(a[391] & b[52])^(a[390] & b[53])^(a[389] & b[54])^(a[388] & b[55])^(a[387] & b[56])^(a[386] & b[57])^(a[385] & b[58])^(a[384] & b[59])^(a[383] & b[60])^(a[382] & b[61])^(a[381] & b[62])^(a[380] & b[63])^(a[379] & b[64])^(a[378] & b[65])^(a[377] & b[66])^(a[376] & b[67])^(a[375] & b[68])^(a[374] & b[69])^(a[373] & b[70])^(a[372] & b[71])^(a[371] & b[72])^(a[370] & b[73])^(a[369] & b[74])^(a[368] & b[75])^(a[367] & b[76])^(a[366] & b[77])^(a[365] & b[78])^(a[364] & b[79])^(a[363] & b[80])^(a[362] & b[81])^(a[361] & b[82])^(a[360] & b[83])^(a[359] & b[84])^(a[358] & b[85])^(a[357] & b[86])^(a[356] & b[87])^(a[355] & b[88])^(a[354] & b[89])^(a[353] & b[90])^(a[352] & b[91])^(a[351] & b[92])^(a[350] & b[93])^(a[349] & b[94])^(a[348] & b[95])^(a[347] & b[96])^(a[346] & b[97])^(a[345] & b[98])^(a[344] & b[99])^(a[343] & b[100])^(a[342] & b[101])^(a[341] & b[102])^(a[340] & b[103])^(a[339] & b[104])^(a[338] & b[105])^(a[337] & b[106])^(a[336] & b[107])^(a[335] & b[108])^(a[334] & b[109])^(a[333] & b[110])^(a[332] & b[111])^(a[331] & b[112])^(a[330] & b[113])^(a[329] & b[114])^(a[328] & b[115])^(a[327] & b[116])^(a[326] & b[117])^(a[325] & b[118])^(a[324] & b[119])^(a[323] & b[120])^(a[322] & b[121])^(a[321] & b[122])^(a[320] & b[123])^(a[319] & b[124])^(a[318] & b[125])^(a[317] & b[126])^(a[316] & b[127])^(a[315] & b[128])^(a[314] & b[129])^(a[313] & b[130])^(a[312] & b[131])^(a[311] & b[132])^(a[310] & b[133])^(a[309] & b[134])^(a[308] & b[135])^(a[307] & b[136])^(a[306] & b[137])^(a[305] & b[138])^(a[304] & b[139])^(a[303] & b[140])^(a[302] & b[141])^(a[301] & b[142])^(a[300] & b[143])^(a[299] & b[144])^(a[298] & b[145])^(a[297] & b[146])^(a[296] & b[147])^(a[295] & b[148])^(a[294] & b[149])^(a[293] & b[150])^(a[292] & b[151])^(a[291] & b[152])^(a[290] & b[153])^(a[289] & b[154])^(a[288] & b[155])^(a[287] & b[156])^(a[286] & b[157])^(a[285] & b[158])^(a[284] & b[159])^(a[283] & b[160])^(a[282] & b[161])^(a[281] & b[162])^(a[280] & b[163])^(a[279] & b[164])^(a[278] & b[165])^(a[277] & b[166])^(a[276] & b[167])^(a[275] & b[168])^(a[274] & b[169])^(a[273] & b[170])^(a[272] & b[171])^(a[271] & b[172])^(a[270] & b[173])^(a[269] & b[174])^(a[268] & b[175])^(a[267] & b[176])^(a[266] & b[177])^(a[265] & b[178])^(a[264] & b[179])^(a[263] & b[180])^(a[262] & b[181])^(a[261] & b[182])^(a[260] & b[183])^(a[259] & b[184])^(a[258] & b[185])^(a[257] & b[186])^(a[256] & b[187])^(a[255] & b[188])^(a[254] & b[189])^(a[253] & b[190])^(a[252] & b[191])^(a[251] & b[192])^(a[250] & b[193])^(a[249] & b[194])^(a[248] & b[195])^(a[247] & b[196])^(a[246] & b[197])^(a[245] & b[198])^(a[244] & b[199])^(a[243] & b[200])^(a[242] & b[201])^(a[241] & b[202])^(a[240] & b[203])^(a[239] & b[204])^(a[238] & b[205])^(a[237] & b[206])^(a[236] & b[207])^(a[235] & b[208])^(a[234] & b[209])^(a[233] & b[210])^(a[232] & b[211])^(a[231] & b[212])^(a[230] & b[213])^(a[229] & b[214])^(a[228] & b[215])^(a[227] & b[216])^(a[226] & b[217])^(a[225] & b[218])^(a[224] & b[219])^(a[223] & b[220])^(a[222] & b[221])^(a[221] & b[222])^(a[220] & b[223])^(a[219] & b[224])^(a[218] & b[225])^(a[217] & b[226])^(a[216] & b[227])^(a[215] & b[228])^(a[214] & b[229])^(a[213] & b[230])^(a[212] & b[231])^(a[211] & b[232])^(a[210] & b[233])^(a[209] & b[234])^(a[208] & b[235])^(a[207] & b[236])^(a[206] & b[237])^(a[205] & b[238])^(a[204] & b[239])^(a[203] & b[240])^(a[202] & b[241])^(a[201] & b[242])^(a[200] & b[243])^(a[199] & b[244])^(a[198] & b[245])^(a[197] & b[246])^(a[196] & b[247])^(a[195] & b[248])^(a[194] & b[249])^(a[193] & b[250])^(a[192] & b[251])^(a[191] & b[252])^(a[190] & b[253])^(a[189] & b[254])^(a[188] & b[255])^(a[187] & b[256])^(a[186] & b[257])^(a[185] & b[258])^(a[184] & b[259])^(a[183] & b[260])^(a[182] & b[261])^(a[181] & b[262])^(a[180] & b[263])^(a[179] & b[264])^(a[178] & b[265])^(a[177] & b[266])^(a[176] & b[267])^(a[175] & b[268])^(a[174] & b[269])^(a[173] & b[270])^(a[172] & b[271])^(a[171] & b[272])^(a[170] & b[273])^(a[169] & b[274])^(a[168] & b[275])^(a[167] & b[276])^(a[166] & b[277])^(a[165] & b[278])^(a[164] & b[279])^(a[163] & b[280])^(a[162] & b[281])^(a[161] & b[282])^(a[160] & b[283])^(a[159] & b[284])^(a[158] & b[285])^(a[157] & b[286])^(a[156] & b[287])^(a[155] & b[288])^(a[154] & b[289])^(a[153] & b[290])^(a[152] & b[291])^(a[151] & b[292])^(a[150] & b[293])^(a[149] & b[294])^(a[148] & b[295])^(a[147] & b[296])^(a[146] & b[297])^(a[145] & b[298])^(a[144] & b[299])^(a[143] & b[300])^(a[142] & b[301])^(a[141] & b[302])^(a[140] & b[303])^(a[139] & b[304])^(a[138] & b[305])^(a[137] & b[306])^(a[136] & b[307])^(a[135] & b[308])^(a[134] & b[309])^(a[133] & b[310])^(a[132] & b[311])^(a[131] & b[312])^(a[130] & b[313])^(a[129] & b[314])^(a[128] & b[315])^(a[127] & b[316])^(a[126] & b[317])^(a[125] & b[318])^(a[124] & b[319])^(a[123] & b[320])^(a[122] & b[321])^(a[121] & b[322])^(a[120] & b[323])^(a[119] & b[324])^(a[118] & b[325])^(a[117] & b[326])^(a[116] & b[327])^(a[115] & b[328])^(a[114] & b[329])^(a[113] & b[330])^(a[112] & b[331])^(a[111] & b[332])^(a[110] & b[333])^(a[109] & b[334])^(a[108] & b[335])^(a[107] & b[336])^(a[106] & b[337])^(a[105] & b[338])^(a[104] & b[339])^(a[103] & b[340])^(a[102] & b[341])^(a[101] & b[342])^(a[100] & b[343])^(a[99] & b[344])^(a[98] & b[345])^(a[97] & b[346])^(a[96] & b[347])^(a[95] & b[348])^(a[94] & b[349])^(a[93] & b[350])^(a[92] & b[351])^(a[91] & b[352])^(a[90] & b[353])^(a[89] & b[354])^(a[88] & b[355])^(a[87] & b[356])^(a[86] & b[357])^(a[85] & b[358])^(a[84] & b[359])^(a[83] & b[360])^(a[82] & b[361])^(a[81] & b[362])^(a[80] & b[363])^(a[79] & b[364])^(a[78] & b[365])^(a[77] & b[366])^(a[76] & b[367])^(a[75] & b[368])^(a[74] & b[369])^(a[73] & b[370])^(a[72] & b[371])^(a[71] & b[372])^(a[70] & b[373])^(a[69] & b[374])^(a[68] & b[375])^(a[67] & b[376])^(a[66] & b[377])^(a[65] & b[378])^(a[64] & b[379])^(a[63] & b[380])^(a[62] & b[381])^(a[61] & b[382])^(a[60] & b[383])^(a[59] & b[384])^(a[58] & b[385])^(a[57] & b[386])^(a[56] & b[387])^(a[55] & b[388])^(a[54] & b[389])^(a[53] & b[390])^(a[52] & b[391])^(a[51] & b[392])^(a[50] & b[393])^(a[49] & b[394])^(a[48] & b[395])^(a[47] & b[396])^(a[46] & b[397])^(a[45] & b[398])^(a[44] & b[399])^(a[43] & b[400])^(a[42] & b[401])^(a[41] & b[402])^(a[40] & b[403])^(a[39] & b[404])^(a[38] & b[405])^(a[37] & b[406])^(a[36] & b[407])^(a[35] & b[408]);
assign y[444] = (a[408] & b[36])^(a[407] & b[37])^(a[406] & b[38])^(a[405] & b[39])^(a[404] & b[40])^(a[403] & b[41])^(a[402] & b[42])^(a[401] & b[43])^(a[400] & b[44])^(a[399] & b[45])^(a[398] & b[46])^(a[397] & b[47])^(a[396] & b[48])^(a[395] & b[49])^(a[394] & b[50])^(a[393] & b[51])^(a[392] & b[52])^(a[391] & b[53])^(a[390] & b[54])^(a[389] & b[55])^(a[388] & b[56])^(a[387] & b[57])^(a[386] & b[58])^(a[385] & b[59])^(a[384] & b[60])^(a[383] & b[61])^(a[382] & b[62])^(a[381] & b[63])^(a[380] & b[64])^(a[379] & b[65])^(a[378] & b[66])^(a[377] & b[67])^(a[376] & b[68])^(a[375] & b[69])^(a[374] & b[70])^(a[373] & b[71])^(a[372] & b[72])^(a[371] & b[73])^(a[370] & b[74])^(a[369] & b[75])^(a[368] & b[76])^(a[367] & b[77])^(a[366] & b[78])^(a[365] & b[79])^(a[364] & b[80])^(a[363] & b[81])^(a[362] & b[82])^(a[361] & b[83])^(a[360] & b[84])^(a[359] & b[85])^(a[358] & b[86])^(a[357] & b[87])^(a[356] & b[88])^(a[355] & b[89])^(a[354] & b[90])^(a[353] & b[91])^(a[352] & b[92])^(a[351] & b[93])^(a[350] & b[94])^(a[349] & b[95])^(a[348] & b[96])^(a[347] & b[97])^(a[346] & b[98])^(a[345] & b[99])^(a[344] & b[100])^(a[343] & b[101])^(a[342] & b[102])^(a[341] & b[103])^(a[340] & b[104])^(a[339] & b[105])^(a[338] & b[106])^(a[337] & b[107])^(a[336] & b[108])^(a[335] & b[109])^(a[334] & b[110])^(a[333] & b[111])^(a[332] & b[112])^(a[331] & b[113])^(a[330] & b[114])^(a[329] & b[115])^(a[328] & b[116])^(a[327] & b[117])^(a[326] & b[118])^(a[325] & b[119])^(a[324] & b[120])^(a[323] & b[121])^(a[322] & b[122])^(a[321] & b[123])^(a[320] & b[124])^(a[319] & b[125])^(a[318] & b[126])^(a[317] & b[127])^(a[316] & b[128])^(a[315] & b[129])^(a[314] & b[130])^(a[313] & b[131])^(a[312] & b[132])^(a[311] & b[133])^(a[310] & b[134])^(a[309] & b[135])^(a[308] & b[136])^(a[307] & b[137])^(a[306] & b[138])^(a[305] & b[139])^(a[304] & b[140])^(a[303] & b[141])^(a[302] & b[142])^(a[301] & b[143])^(a[300] & b[144])^(a[299] & b[145])^(a[298] & b[146])^(a[297] & b[147])^(a[296] & b[148])^(a[295] & b[149])^(a[294] & b[150])^(a[293] & b[151])^(a[292] & b[152])^(a[291] & b[153])^(a[290] & b[154])^(a[289] & b[155])^(a[288] & b[156])^(a[287] & b[157])^(a[286] & b[158])^(a[285] & b[159])^(a[284] & b[160])^(a[283] & b[161])^(a[282] & b[162])^(a[281] & b[163])^(a[280] & b[164])^(a[279] & b[165])^(a[278] & b[166])^(a[277] & b[167])^(a[276] & b[168])^(a[275] & b[169])^(a[274] & b[170])^(a[273] & b[171])^(a[272] & b[172])^(a[271] & b[173])^(a[270] & b[174])^(a[269] & b[175])^(a[268] & b[176])^(a[267] & b[177])^(a[266] & b[178])^(a[265] & b[179])^(a[264] & b[180])^(a[263] & b[181])^(a[262] & b[182])^(a[261] & b[183])^(a[260] & b[184])^(a[259] & b[185])^(a[258] & b[186])^(a[257] & b[187])^(a[256] & b[188])^(a[255] & b[189])^(a[254] & b[190])^(a[253] & b[191])^(a[252] & b[192])^(a[251] & b[193])^(a[250] & b[194])^(a[249] & b[195])^(a[248] & b[196])^(a[247] & b[197])^(a[246] & b[198])^(a[245] & b[199])^(a[244] & b[200])^(a[243] & b[201])^(a[242] & b[202])^(a[241] & b[203])^(a[240] & b[204])^(a[239] & b[205])^(a[238] & b[206])^(a[237] & b[207])^(a[236] & b[208])^(a[235] & b[209])^(a[234] & b[210])^(a[233] & b[211])^(a[232] & b[212])^(a[231] & b[213])^(a[230] & b[214])^(a[229] & b[215])^(a[228] & b[216])^(a[227] & b[217])^(a[226] & b[218])^(a[225] & b[219])^(a[224] & b[220])^(a[223] & b[221])^(a[222] & b[222])^(a[221] & b[223])^(a[220] & b[224])^(a[219] & b[225])^(a[218] & b[226])^(a[217] & b[227])^(a[216] & b[228])^(a[215] & b[229])^(a[214] & b[230])^(a[213] & b[231])^(a[212] & b[232])^(a[211] & b[233])^(a[210] & b[234])^(a[209] & b[235])^(a[208] & b[236])^(a[207] & b[237])^(a[206] & b[238])^(a[205] & b[239])^(a[204] & b[240])^(a[203] & b[241])^(a[202] & b[242])^(a[201] & b[243])^(a[200] & b[244])^(a[199] & b[245])^(a[198] & b[246])^(a[197] & b[247])^(a[196] & b[248])^(a[195] & b[249])^(a[194] & b[250])^(a[193] & b[251])^(a[192] & b[252])^(a[191] & b[253])^(a[190] & b[254])^(a[189] & b[255])^(a[188] & b[256])^(a[187] & b[257])^(a[186] & b[258])^(a[185] & b[259])^(a[184] & b[260])^(a[183] & b[261])^(a[182] & b[262])^(a[181] & b[263])^(a[180] & b[264])^(a[179] & b[265])^(a[178] & b[266])^(a[177] & b[267])^(a[176] & b[268])^(a[175] & b[269])^(a[174] & b[270])^(a[173] & b[271])^(a[172] & b[272])^(a[171] & b[273])^(a[170] & b[274])^(a[169] & b[275])^(a[168] & b[276])^(a[167] & b[277])^(a[166] & b[278])^(a[165] & b[279])^(a[164] & b[280])^(a[163] & b[281])^(a[162] & b[282])^(a[161] & b[283])^(a[160] & b[284])^(a[159] & b[285])^(a[158] & b[286])^(a[157] & b[287])^(a[156] & b[288])^(a[155] & b[289])^(a[154] & b[290])^(a[153] & b[291])^(a[152] & b[292])^(a[151] & b[293])^(a[150] & b[294])^(a[149] & b[295])^(a[148] & b[296])^(a[147] & b[297])^(a[146] & b[298])^(a[145] & b[299])^(a[144] & b[300])^(a[143] & b[301])^(a[142] & b[302])^(a[141] & b[303])^(a[140] & b[304])^(a[139] & b[305])^(a[138] & b[306])^(a[137] & b[307])^(a[136] & b[308])^(a[135] & b[309])^(a[134] & b[310])^(a[133] & b[311])^(a[132] & b[312])^(a[131] & b[313])^(a[130] & b[314])^(a[129] & b[315])^(a[128] & b[316])^(a[127] & b[317])^(a[126] & b[318])^(a[125] & b[319])^(a[124] & b[320])^(a[123] & b[321])^(a[122] & b[322])^(a[121] & b[323])^(a[120] & b[324])^(a[119] & b[325])^(a[118] & b[326])^(a[117] & b[327])^(a[116] & b[328])^(a[115] & b[329])^(a[114] & b[330])^(a[113] & b[331])^(a[112] & b[332])^(a[111] & b[333])^(a[110] & b[334])^(a[109] & b[335])^(a[108] & b[336])^(a[107] & b[337])^(a[106] & b[338])^(a[105] & b[339])^(a[104] & b[340])^(a[103] & b[341])^(a[102] & b[342])^(a[101] & b[343])^(a[100] & b[344])^(a[99] & b[345])^(a[98] & b[346])^(a[97] & b[347])^(a[96] & b[348])^(a[95] & b[349])^(a[94] & b[350])^(a[93] & b[351])^(a[92] & b[352])^(a[91] & b[353])^(a[90] & b[354])^(a[89] & b[355])^(a[88] & b[356])^(a[87] & b[357])^(a[86] & b[358])^(a[85] & b[359])^(a[84] & b[360])^(a[83] & b[361])^(a[82] & b[362])^(a[81] & b[363])^(a[80] & b[364])^(a[79] & b[365])^(a[78] & b[366])^(a[77] & b[367])^(a[76] & b[368])^(a[75] & b[369])^(a[74] & b[370])^(a[73] & b[371])^(a[72] & b[372])^(a[71] & b[373])^(a[70] & b[374])^(a[69] & b[375])^(a[68] & b[376])^(a[67] & b[377])^(a[66] & b[378])^(a[65] & b[379])^(a[64] & b[380])^(a[63] & b[381])^(a[62] & b[382])^(a[61] & b[383])^(a[60] & b[384])^(a[59] & b[385])^(a[58] & b[386])^(a[57] & b[387])^(a[56] & b[388])^(a[55] & b[389])^(a[54] & b[390])^(a[53] & b[391])^(a[52] & b[392])^(a[51] & b[393])^(a[50] & b[394])^(a[49] & b[395])^(a[48] & b[396])^(a[47] & b[397])^(a[46] & b[398])^(a[45] & b[399])^(a[44] & b[400])^(a[43] & b[401])^(a[42] & b[402])^(a[41] & b[403])^(a[40] & b[404])^(a[39] & b[405])^(a[38] & b[406])^(a[37] & b[407])^(a[36] & b[408]);
assign y[445] = (a[408] & b[37])^(a[407] & b[38])^(a[406] & b[39])^(a[405] & b[40])^(a[404] & b[41])^(a[403] & b[42])^(a[402] & b[43])^(a[401] & b[44])^(a[400] & b[45])^(a[399] & b[46])^(a[398] & b[47])^(a[397] & b[48])^(a[396] & b[49])^(a[395] & b[50])^(a[394] & b[51])^(a[393] & b[52])^(a[392] & b[53])^(a[391] & b[54])^(a[390] & b[55])^(a[389] & b[56])^(a[388] & b[57])^(a[387] & b[58])^(a[386] & b[59])^(a[385] & b[60])^(a[384] & b[61])^(a[383] & b[62])^(a[382] & b[63])^(a[381] & b[64])^(a[380] & b[65])^(a[379] & b[66])^(a[378] & b[67])^(a[377] & b[68])^(a[376] & b[69])^(a[375] & b[70])^(a[374] & b[71])^(a[373] & b[72])^(a[372] & b[73])^(a[371] & b[74])^(a[370] & b[75])^(a[369] & b[76])^(a[368] & b[77])^(a[367] & b[78])^(a[366] & b[79])^(a[365] & b[80])^(a[364] & b[81])^(a[363] & b[82])^(a[362] & b[83])^(a[361] & b[84])^(a[360] & b[85])^(a[359] & b[86])^(a[358] & b[87])^(a[357] & b[88])^(a[356] & b[89])^(a[355] & b[90])^(a[354] & b[91])^(a[353] & b[92])^(a[352] & b[93])^(a[351] & b[94])^(a[350] & b[95])^(a[349] & b[96])^(a[348] & b[97])^(a[347] & b[98])^(a[346] & b[99])^(a[345] & b[100])^(a[344] & b[101])^(a[343] & b[102])^(a[342] & b[103])^(a[341] & b[104])^(a[340] & b[105])^(a[339] & b[106])^(a[338] & b[107])^(a[337] & b[108])^(a[336] & b[109])^(a[335] & b[110])^(a[334] & b[111])^(a[333] & b[112])^(a[332] & b[113])^(a[331] & b[114])^(a[330] & b[115])^(a[329] & b[116])^(a[328] & b[117])^(a[327] & b[118])^(a[326] & b[119])^(a[325] & b[120])^(a[324] & b[121])^(a[323] & b[122])^(a[322] & b[123])^(a[321] & b[124])^(a[320] & b[125])^(a[319] & b[126])^(a[318] & b[127])^(a[317] & b[128])^(a[316] & b[129])^(a[315] & b[130])^(a[314] & b[131])^(a[313] & b[132])^(a[312] & b[133])^(a[311] & b[134])^(a[310] & b[135])^(a[309] & b[136])^(a[308] & b[137])^(a[307] & b[138])^(a[306] & b[139])^(a[305] & b[140])^(a[304] & b[141])^(a[303] & b[142])^(a[302] & b[143])^(a[301] & b[144])^(a[300] & b[145])^(a[299] & b[146])^(a[298] & b[147])^(a[297] & b[148])^(a[296] & b[149])^(a[295] & b[150])^(a[294] & b[151])^(a[293] & b[152])^(a[292] & b[153])^(a[291] & b[154])^(a[290] & b[155])^(a[289] & b[156])^(a[288] & b[157])^(a[287] & b[158])^(a[286] & b[159])^(a[285] & b[160])^(a[284] & b[161])^(a[283] & b[162])^(a[282] & b[163])^(a[281] & b[164])^(a[280] & b[165])^(a[279] & b[166])^(a[278] & b[167])^(a[277] & b[168])^(a[276] & b[169])^(a[275] & b[170])^(a[274] & b[171])^(a[273] & b[172])^(a[272] & b[173])^(a[271] & b[174])^(a[270] & b[175])^(a[269] & b[176])^(a[268] & b[177])^(a[267] & b[178])^(a[266] & b[179])^(a[265] & b[180])^(a[264] & b[181])^(a[263] & b[182])^(a[262] & b[183])^(a[261] & b[184])^(a[260] & b[185])^(a[259] & b[186])^(a[258] & b[187])^(a[257] & b[188])^(a[256] & b[189])^(a[255] & b[190])^(a[254] & b[191])^(a[253] & b[192])^(a[252] & b[193])^(a[251] & b[194])^(a[250] & b[195])^(a[249] & b[196])^(a[248] & b[197])^(a[247] & b[198])^(a[246] & b[199])^(a[245] & b[200])^(a[244] & b[201])^(a[243] & b[202])^(a[242] & b[203])^(a[241] & b[204])^(a[240] & b[205])^(a[239] & b[206])^(a[238] & b[207])^(a[237] & b[208])^(a[236] & b[209])^(a[235] & b[210])^(a[234] & b[211])^(a[233] & b[212])^(a[232] & b[213])^(a[231] & b[214])^(a[230] & b[215])^(a[229] & b[216])^(a[228] & b[217])^(a[227] & b[218])^(a[226] & b[219])^(a[225] & b[220])^(a[224] & b[221])^(a[223] & b[222])^(a[222] & b[223])^(a[221] & b[224])^(a[220] & b[225])^(a[219] & b[226])^(a[218] & b[227])^(a[217] & b[228])^(a[216] & b[229])^(a[215] & b[230])^(a[214] & b[231])^(a[213] & b[232])^(a[212] & b[233])^(a[211] & b[234])^(a[210] & b[235])^(a[209] & b[236])^(a[208] & b[237])^(a[207] & b[238])^(a[206] & b[239])^(a[205] & b[240])^(a[204] & b[241])^(a[203] & b[242])^(a[202] & b[243])^(a[201] & b[244])^(a[200] & b[245])^(a[199] & b[246])^(a[198] & b[247])^(a[197] & b[248])^(a[196] & b[249])^(a[195] & b[250])^(a[194] & b[251])^(a[193] & b[252])^(a[192] & b[253])^(a[191] & b[254])^(a[190] & b[255])^(a[189] & b[256])^(a[188] & b[257])^(a[187] & b[258])^(a[186] & b[259])^(a[185] & b[260])^(a[184] & b[261])^(a[183] & b[262])^(a[182] & b[263])^(a[181] & b[264])^(a[180] & b[265])^(a[179] & b[266])^(a[178] & b[267])^(a[177] & b[268])^(a[176] & b[269])^(a[175] & b[270])^(a[174] & b[271])^(a[173] & b[272])^(a[172] & b[273])^(a[171] & b[274])^(a[170] & b[275])^(a[169] & b[276])^(a[168] & b[277])^(a[167] & b[278])^(a[166] & b[279])^(a[165] & b[280])^(a[164] & b[281])^(a[163] & b[282])^(a[162] & b[283])^(a[161] & b[284])^(a[160] & b[285])^(a[159] & b[286])^(a[158] & b[287])^(a[157] & b[288])^(a[156] & b[289])^(a[155] & b[290])^(a[154] & b[291])^(a[153] & b[292])^(a[152] & b[293])^(a[151] & b[294])^(a[150] & b[295])^(a[149] & b[296])^(a[148] & b[297])^(a[147] & b[298])^(a[146] & b[299])^(a[145] & b[300])^(a[144] & b[301])^(a[143] & b[302])^(a[142] & b[303])^(a[141] & b[304])^(a[140] & b[305])^(a[139] & b[306])^(a[138] & b[307])^(a[137] & b[308])^(a[136] & b[309])^(a[135] & b[310])^(a[134] & b[311])^(a[133] & b[312])^(a[132] & b[313])^(a[131] & b[314])^(a[130] & b[315])^(a[129] & b[316])^(a[128] & b[317])^(a[127] & b[318])^(a[126] & b[319])^(a[125] & b[320])^(a[124] & b[321])^(a[123] & b[322])^(a[122] & b[323])^(a[121] & b[324])^(a[120] & b[325])^(a[119] & b[326])^(a[118] & b[327])^(a[117] & b[328])^(a[116] & b[329])^(a[115] & b[330])^(a[114] & b[331])^(a[113] & b[332])^(a[112] & b[333])^(a[111] & b[334])^(a[110] & b[335])^(a[109] & b[336])^(a[108] & b[337])^(a[107] & b[338])^(a[106] & b[339])^(a[105] & b[340])^(a[104] & b[341])^(a[103] & b[342])^(a[102] & b[343])^(a[101] & b[344])^(a[100] & b[345])^(a[99] & b[346])^(a[98] & b[347])^(a[97] & b[348])^(a[96] & b[349])^(a[95] & b[350])^(a[94] & b[351])^(a[93] & b[352])^(a[92] & b[353])^(a[91] & b[354])^(a[90] & b[355])^(a[89] & b[356])^(a[88] & b[357])^(a[87] & b[358])^(a[86] & b[359])^(a[85] & b[360])^(a[84] & b[361])^(a[83] & b[362])^(a[82] & b[363])^(a[81] & b[364])^(a[80] & b[365])^(a[79] & b[366])^(a[78] & b[367])^(a[77] & b[368])^(a[76] & b[369])^(a[75] & b[370])^(a[74] & b[371])^(a[73] & b[372])^(a[72] & b[373])^(a[71] & b[374])^(a[70] & b[375])^(a[69] & b[376])^(a[68] & b[377])^(a[67] & b[378])^(a[66] & b[379])^(a[65] & b[380])^(a[64] & b[381])^(a[63] & b[382])^(a[62] & b[383])^(a[61] & b[384])^(a[60] & b[385])^(a[59] & b[386])^(a[58] & b[387])^(a[57] & b[388])^(a[56] & b[389])^(a[55] & b[390])^(a[54] & b[391])^(a[53] & b[392])^(a[52] & b[393])^(a[51] & b[394])^(a[50] & b[395])^(a[49] & b[396])^(a[48] & b[397])^(a[47] & b[398])^(a[46] & b[399])^(a[45] & b[400])^(a[44] & b[401])^(a[43] & b[402])^(a[42] & b[403])^(a[41] & b[404])^(a[40] & b[405])^(a[39] & b[406])^(a[38] & b[407])^(a[37] & b[408]);
assign y[446] = (a[408] & b[38])^(a[407] & b[39])^(a[406] & b[40])^(a[405] & b[41])^(a[404] & b[42])^(a[403] & b[43])^(a[402] & b[44])^(a[401] & b[45])^(a[400] & b[46])^(a[399] & b[47])^(a[398] & b[48])^(a[397] & b[49])^(a[396] & b[50])^(a[395] & b[51])^(a[394] & b[52])^(a[393] & b[53])^(a[392] & b[54])^(a[391] & b[55])^(a[390] & b[56])^(a[389] & b[57])^(a[388] & b[58])^(a[387] & b[59])^(a[386] & b[60])^(a[385] & b[61])^(a[384] & b[62])^(a[383] & b[63])^(a[382] & b[64])^(a[381] & b[65])^(a[380] & b[66])^(a[379] & b[67])^(a[378] & b[68])^(a[377] & b[69])^(a[376] & b[70])^(a[375] & b[71])^(a[374] & b[72])^(a[373] & b[73])^(a[372] & b[74])^(a[371] & b[75])^(a[370] & b[76])^(a[369] & b[77])^(a[368] & b[78])^(a[367] & b[79])^(a[366] & b[80])^(a[365] & b[81])^(a[364] & b[82])^(a[363] & b[83])^(a[362] & b[84])^(a[361] & b[85])^(a[360] & b[86])^(a[359] & b[87])^(a[358] & b[88])^(a[357] & b[89])^(a[356] & b[90])^(a[355] & b[91])^(a[354] & b[92])^(a[353] & b[93])^(a[352] & b[94])^(a[351] & b[95])^(a[350] & b[96])^(a[349] & b[97])^(a[348] & b[98])^(a[347] & b[99])^(a[346] & b[100])^(a[345] & b[101])^(a[344] & b[102])^(a[343] & b[103])^(a[342] & b[104])^(a[341] & b[105])^(a[340] & b[106])^(a[339] & b[107])^(a[338] & b[108])^(a[337] & b[109])^(a[336] & b[110])^(a[335] & b[111])^(a[334] & b[112])^(a[333] & b[113])^(a[332] & b[114])^(a[331] & b[115])^(a[330] & b[116])^(a[329] & b[117])^(a[328] & b[118])^(a[327] & b[119])^(a[326] & b[120])^(a[325] & b[121])^(a[324] & b[122])^(a[323] & b[123])^(a[322] & b[124])^(a[321] & b[125])^(a[320] & b[126])^(a[319] & b[127])^(a[318] & b[128])^(a[317] & b[129])^(a[316] & b[130])^(a[315] & b[131])^(a[314] & b[132])^(a[313] & b[133])^(a[312] & b[134])^(a[311] & b[135])^(a[310] & b[136])^(a[309] & b[137])^(a[308] & b[138])^(a[307] & b[139])^(a[306] & b[140])^(a[305] & b[141])^(a[304] & b[142])^(a[303] & b[143])^(a[302] & b[144])^(a[301] & b[145])^(a[300] & b[146])^(a[299] & b[147])^(a[298] & b[148])^(a[297] & b[149])^(a[296] & b[150])^(a[295] & b[151])^(a[294] & b[152])^(a[293] & b[153])^(a[292] & b[154])^(a[291] & b[155])^(a[290] & b[156])^(a[289] & b[157])^(a[288] & b[158])^(a[287] & b[159])^(a[286] & b[160])^(a[285] & b[161])^(a[284] & b[162])^(a[283] & b[163])^(a[282] & b[164])^(a[281] & b[165])^(a[280] & b[166])^(a[279] & b[167])^(a[278] & b[168])^(a[277] & b[169])^(a[276] & b[170])^(a[275] & b[171])^(a[274] & b[172])^(a[273] & b[173])^(a[272] & b[174])^(a[271] & b[175])^(a[270] & b[176])^(a[269] & b[177])^(a[268] & b[178])^(a[267] & b[179])^(a[266] & b[180])^(a[265] & b[181])^(a[264] & b[182])^(a[263] & b[183])^(a[262] & b[184])^(a[261] & b[185])^(a[260] & b[186])^(a[259] & b[187])^(a[258] & b[188])^(a[257] & b[189])^(a[256] & b[190])^(a[255] & b[191])^(a[254] & b[192])^(a[253] & b[193])^(a[252] & b[194])^(a[251] & b[195])^(a[250] & b[196])^(a[249] & b[197])^(a[248] & b[198])^(a[247] & b[199])^(a[246] & b[200])^(a[245] & b[201])^(a[244] & b[202])^(a[243] & b[203])^(a[242] & b[204])^(a[241] & b[205])^(a[240] & b[206])^(a[239] & b[207])^(a[238] & b[208])^(a[237] & b[209])^(a[236] & b[210])^(a[235] & b[211])^(a[234] & b[212])^(a[233] & b[213])^(a[232] & b[214])^(a[231] & b[215])^(a[230] & b[216])^(a[229] & b[217])^(a[228] & b[218])^(a[227] & b[219])^(a[226] & b[220])^(a[225] & b[221])^(a[224] & b[222])^(a[223] & b[223])^(a[222] & b[224])^(a[221] & b[225])^(a[220] & b[226])^(a[219] & b[227])^(a[218] & b[228])^(a[217] & b[229])^(a[216] & b[230])^(a[215] & b[231])^(a[214] & b[232])^(a[213] & b[233])^(a[212] & b[234])^(a[211] & b[235])^(a[210] & b[236])^(a[209] & b[237])^(a[208] & b[238])^(a[207] & b[239])^(a[206] & b[240])^(a[205] & b[241])^(a[204] & b[242])^(a[203] & b[243])^(a[202] & b[244])^(a[201] & b[245])^(a[200] & b[246])^(a[199] & b[247])^(a[198] & b[248])^(a[197] & b[249])^(a[196] & b[250])^(a[195] & b[251])^(a[194] & b[252])^(a[193] & b[253])^(a[192] & b[254])^(a[191] & b[255])^(a[190] & b[256])^(a[189] & b[257])^(a[188] & b[258])^(a[187] & b[259])^(a[186] & b[260])^(a[185] & b[261])^(a[184] & b[262])^(a[183] & b[263])^(a[182] & b[264])^(a[181] & b[265])^(a[180] & b[266])^(a[179] & b[267])^(a[178] & b[268])^(a[177] & b[269])^(a[176] & b[270])^(a[175] & b[271])^(a[174] & b[272])^(a[173] & b[273])^(a[172] & b[274])^(a[171] & b[275])^(a[170] & b[276])^(a[169] & b[277])^(a[168] & b[278])^(a[167] & b[279])^(a[166] & b[280])^(a[165] & b[281])^(a[164] & b[282])^(a[163] & b[283])^(a[162] & b[284])^(a[161] & b[285])^(a[160] & b[286])^(a[159] & b[287])^(a[158] & b[288])^(a[157] & b[289])^(a[156] & b[290])^(a[155] & b[291])^(a[154] & b[292])^(a[153] & b[293])^(a[152] & b[294])^(a[151] & b[295])^(a[150] & b[296])^(a[149] & b[297])^(a[148] & b[298])^(a[147] & b[299])^(a[146] & b[300])^(a[145] & b[301])^(a[144] & b[302])^(a[143] & b[303])^(a[142] & b[304])^(a[141] & b[305])^(a[140] & b[306])^(a[139] & b[307])^(a[138] & b[308])^(a[137] & b[309])^(a[136] & b[310])^(a[135] & b[311])^(a[134] & b[312])^(a[133] & b[313])^(a[132] & b[314])^(a[131] & b[315])^(a[130] & b[316])^(a[129] & b[317])^(a[128] & b[318])^(a[127] & b[319])^(a[126] & b[320])^(a[125] & b[321])^(a[124] & b[322])^(a[123] & b[323])^(a[122] & b[324])^(a[121] & b[325])^(a[120] & b[326])^(a[119] & b[327])^(a[118] & b[328])^(a[117] & b[329])^(a[116] & b[330])^(a[115] & b[331])^(a[114] & b[332])^(a[113] & b[333])^(a[112] & b[334])^(a[111] & b[335])^(a[110] & b[336])^(a[109] & b[337])^(a[108] & b[338])^(a[107] & b[339])^(a[106] & b[340])^(a[105] & b[341])^(a[104] & b[342])^(a[103] & b[343])^(a[102] & b[344])^(a[101] & b[345])^(a[100] & b[346])^(a[99] & b[347])^(a[98] & b[348])^(a[97] & b[349])^(a[96] & b[350])^(a[95] & b[351])^(a[94] & b[352])^(a[93] & b[353])^(a[92] & b[354])^(a[91] & b[355])^(a[90] & b[356])^(a[89] & b[357])^(a[88] & b[358])^(a[87] & b[359])^(a[86] & b[360])^(a[85] & b[361])^(a[84] & b[362])^(a[83] & b[363])^(a[82] & b[364])^(a[81] & b[365])^(a[80] & b[366])^(a[79] & b[367])^(a[78] & b[368])^(a[77] & b[369])^(a[76] & b[370])^(a[75] & b[371])^(a[74] & b[372])^(a[73] & b[373])^(a[72] & b[374])^(a[71] & b[375])^(a[70] & b[376])^(a[69] & b[377])^(a[68] & b[378])^(a[67] & b[379])^(a[66] & b[380])^(a[65] & b[381])^(a[64] & b[382])^(a[63] & b[383])^(a[62] & b[384])^(a[61] & b[385])^(a[60] & b[386])^(a[59] & b[387])^(a[58] & b[388])^(a[57] & b[389])^(a[56] & b[390])^(a[55] & b[391])^(a[54] & b[392])^(a[53] & b[393])^(a[52] & b[394])^(a[51] & b[395])^(a[50] & b[396])^(a[49] & b[397])^(a[48] & b[398])^(a[47] & b[399])^(a[46] & b[400])^(a[45] & b[401])^(a[44] & b[402])^(a[43] & b[403])^(a[42] & b[404])^(a[41] & b[405])^(a[40] & b[406])^(a[39] & b[407])^(a[38] & b[408]);
assign y[447] = (a[408] & b[39])^(a[407] & b[40])^(a[406] & b[41])^(a[405] & b[42])^(a[404] & b[43])^(a[403] & b[44])^(a[402] & b[45])^(a[401] & b[46])^(a[400] & b[47])^(a[399] & b[48])^(a[398] & b[49])^(a[397] & b[50])^(a[396] & b[51])^(a[395] & b[52])^(a[394] & b[53])^(a[393] & b[54])^(a[392] & b[55])^(a[391] & b[56])^(a[390] & b[57])^(a[389] & b[58])^(a[388] & b[59])^(a[387] & b[60])^(a[386] & b[61])^(a[385] & b[62])^(a[384] & b[63])^(a[383] & b[64])^(a[382] & b[65])^(a[381] & b[66])^(a[380] & b[67])^(a[379] & b[68])^(a[378] & b[69])^(a[377] & b[70])^(a[376] & b[71])^(a[375] & b[72])^(a[374] & b[73])^(a[373] & b[74])^(a[372] & b[75])^(a[371] & b[76])^(a[370] & b[77])^(a[369] & b[78])^(a[368] & b[79])^(a[367] & b[80])^(a[366] & b[81])^(a[365] & b[82])^(a[364] & b[83])^(a[363] & b[84])^(a[362] & b[85])^(a[361] & b[86])^(a[360] & b[87])^(a[359] & b[88])^(a[358] & b[89])^(a[357] & b[90])^(a[356] & b[91])^(a[355] & b[92])^(a[354] & b[93])^(a[353] & b[94])^(a[352] & b[95])^(a[351] & b[96])^(a[350] & b[97])^(a[349] & b[98])^(a[348] & b[99])^(a[347] & b[100])^(a[346] & b[101])^(a[345] & b[102])^(a[344] & b[103])^(a[343] & b[104])^(a[342] & b[105])^(a[341] & b[106])^(a[340] & b[107])^(a[339] & b[108])^(a[338] & b[109])^(a[337] & b[110])^(a[336] & b[111])^(a[335] & b[112])^(a[334] & b[113])^(a[333] & b[114])^(a[332] & b[115])^(a[331] & b[116])^(a[330] & b[117])^(a[329] & b[118])^(a[328] & b[119])^(a[327] & b[120])^(a[326] & b[121])^(a[325] & b[122])^(a[324] & b[123])^(a[323] & b[124])^(a[322] & b[125])^(a[321] & b[126])^(a[320] & b[127])^(a[319] & b[128])^(a[318] & b[129])^(a[317] & b[130])^(a[316] & b[131])^(a[315] & b[132])^(a[314] & b[133])^(a[313] & b[134])^(a[312] & b[135])^(a[311] & b[136])^(a[310] & b[137])^(a[309] & b[138])^(a[308] & b[139])^(a[307] & b[140])^(a[306] & b[141])^(a[305] & b[142])^(a[304] & b[143])^(a[303] & b[144])^(a[302] & b[145])^(a[301] & b[146])^(a[300] & b[147])^(a[299] & b[148])^(a[298] & b[149])^(a[297] & b[150])^(a[296] & b[151])^(a[295] & b[152])^(a[294] & b[153])^(a[293] & b[154])^(a[292] & b[155])^(a[291] & b[156])^(a[290] & b[157])^(a[289] & b[158])^(a[288] & b[159])^(a[287] & b[160])^(a[286] & b[161])^(a[285] & b[162])^(a[284] & b[163])^(a[283] & b[164])^(a[282] & b[165])^(a[281] & b[166])^(a[280] & b[167])^(a[279] & b[168])^(a[278] & b[169])^(a[277] & b[170])^(a[276] & b[171])^(a[275] & b[172])^(a[274] & b[173])^(a[273] & b[174])^(a[272] & b[175])^(a[271] & b[176])^(a[270] & b[177])^(a[269] & b[178])^(a[268] & b[179])^(a[267] & b[180])^(a[266] & b[181])^(a[265] & b[182])^(a[264] & b[183])^(a[263] & b[184])^(a[262] & b[185])^(a[261] & b[186])^(a[260] & b[187])^(a[259] & b[188])^(a[258] & b[189])^(a[257] & b[190])^(a[256] & b[191])^(a[255] & b[192])^(a[254] & b[193])^(a[253] & b[194])^(a[252] & b[195])^(a[251] & b[196])^(a[250] & b[197])^(a[249] & b[198])^(a[248] & b[199])^(a[247] & b[200])^(a[246] & b[201])^(a[245] & b[202])^(a[244] & b[203])^(a[243] & b[204])^(a[242] & b[205])^(a[241] & b[206])^(a[240] & b[207])^(a[239] & b[208])^(a[238] & b[209])^(a[237] & b[210])^(a[236] & b[211])^(a[235] & b[212])^(a[234] & b[213])^(a[233] & b[214])^(a[232] & b[215])^(a[231] & b[216])^(a[230] & b[217])^(a[229] & b[218])^(a[228] & b[219])^(a[227] & b[220])^(a[226] & b[221])^(a[225] & b[222])^(a[224] & b[223])^(a[223] & b[224])^(a[222] & b[225])^(a[221] & b[226])^(a[220] & b[227])^(a[219] & b[228])^(a[218] & b[229])^(a[217] & b[230])^(a[216] & b[231])^(a[215] & b[232])^(a[214] & b[233])^(a[213] & b[234])^(a[212] & b[235])^(a[211] & b[236])^(a[210] & b[237])^(a[209] & b[238])^(a[208] & b[239])^(a[207] & b[240])^(a[206] & b[241])^(a[205] & b[242])^(a[204] & b[243])^(a[203] & b[244])^(a[202] & b[245])^(a[201] & b[246])^(a[200] & b[247])^(a[199] & b[248])^(a[198] & b[249])^(a[197] & b[250])^(a[196] & b[251])^(a[195] & b[252])^(a[194] & b[253])^(a[193] & b[254])^(a[192] & b[255])^(a[191] & b[256])^(a[190] & b[257])^(a[189] & b[258])^(a[188] & b[259])^(a[187] & b[260])^(a[186] & b[261])^(a[185] & b[262])^(a[184] & b[263])^(a[183] & b[264])^(a[182] & b[265])^(a[181] & b[266])^(a[180] & b[267])^(a[179] & b[268])^(a[178] & b[269])^(a[177] & b[270])^(a[176] & b[271])^(a[175] & b[272])^(a[174] & b[273])^(a[173] & b[274])^(a[172] & b[275])^(a[171] & b[276])^(a[170] & b[277])^(a[169] & b[278])^(a[168] & b[279])^(a[167] & b[280])^(a[166] & b[281])^(a[165] & b[282])^(a[164] & b[283])^(a[163] & b[284])^(a[162] & b[285])^(a[161] & b[286])^(a[160] & b[287])^(a[159] & b[288])^(a[158] & b[289])^(a[157] & b[290])^(a[156] & b[291])^(a[155] & b[292])^(a[154] & b[293])^(a[153] & b[294])^(a[152] & b[295])^(a[151] & b[296])^(a[150] & b[297])^(a[149] & b[298])^(a[148] & b[299])^(a[147] & b[300])^(a[146] & b[301])^(a[145] & b[302])^(a[144] & b[303])^(a[143] & b[304])^(a[142] & b[305])^(a[141] & b[306])^(a[140] & b[307])^(a[139] & b[308])^(a[138] & b[309])^(a[137] & b[310])^(a[136] & b[311])^(a[135] & b[312])^(a[134] & b[313])^(a[133] & b[314])^(a[132] & b[315])^(a[131] & b[316])^(a[130] & b[317])^(a[129] & b[318])^(a[128] & b[319])^(a[127] & b[320])^(a[126] & b[321])^(a[125] & b[322])^(a[124] & b[323])^(a[123] & b[324])^(a[122] & b[325])^(a[121] & b[326])^(a[120] & b[327])^(a[119] & b[328])^(a[118] & b[329])^(a[117] & b[330])^(a[116] & b[331])^(a[115] & b[332])^(a[114] & b[333])^(a[113] & b[334])^(a[112] & b[335])^(a[111] & b[336])^(a[110] & b[337])^(a[109] & b[338])^(a[108] & b[339])^(a[107] & b[340])^(a[106] & b[341])^(a[105] & b[342])^(a[104] & b[343])^(a[103] & b[344])^(a[102] & b[345])^(a[101] & b[346])^(a[100] & b[347])^(a[99] & b[348])^(a[98] & b[349])^(a[97] & b[350])^(a[96] & b[351])^(a[95] & b[352])^(a[94] & b[353])^(a[93] & b[354])^(a[92] & b[355])^(a[91] & b[356])^(a[90] & b[357])^(a[89] & b[358])^(a[88] & b[359])^(a[87] & b[360])^(a[86] & b[361])^(a[85] & b[362])^(a[84] & b[363])^(a[83] & b[364])^(a[82] & b[365])^(a[81] & b[366])^(a[80] & b[367])^(a[79] & b[368])^(a[78] & b[369])^(a[77] & b[370])^(a[76] & b[371])^(a[75] & b[372])^(a[74] & b[373])^(a[73] & b[374])^(a[72] & b[375])^(a[71] & b[376])^(a[70] & b[377])^(a[69] & b[378])^(a[68] & b[379])^(a[67] & b[380])^(a[66] & b[381])^(a[65] & b[382])^(a[64] & b[383])^(a[63] & b[384])^(a[62] & b[385])^(a[61] & b[386])^(a[60] & b[387])^(a[59] & b[388])^(a[58] & b[389])^(a[57] & b[390])^(a[56] & b[391])^(a[55] & b[392])^(a[54] & b[393])^(a[53] & b[394])^(a[52] & b[395])^(a[51] & b[396])^(a[50] & b[397])^(a[49] & b[398])^(a[48] & b[399])^(a[47] & b[400])^(a[46] & b[401])^(a[45] & b[402])^(a[44] & b[403])^(a[43] & b[404])^(a[42] & b[405])^(a[41] & b[406])^(a[40] & b[407])^(a[39] & b[408]);
assign y[448] = (a[408] & b[40])^(a[407] & b[41])^(a[406] & b[42])^(a[405] & b[43])^(a[404] & b[44])^(a[403] & b[45])^(a[402] & b[46])^(a[401] & b[47])^(a[400] & b[48])^(a[399] & b[49])^(a[398] & b[50])^(a[397] & b[51])^(a[396] & b[52])^(a[395] & b[53])^(a[394] & b[54])^(a[393] & b[55])^(a[392] & b[56])^(a[391] & b[57])^(a[390] & b[58])^(a[389] & b[59])^(a[388] & b[60])^(a[387] & b[61])^(a[386] & b[62])^(a[385] & b[63])^(a[384] & b[64])^(a[383] & b[65])^(a[382] & b[66])^(a[381] & b[67])^(a[380] & b[68])^(a[379] & b[69])^(a[378] & b[70])^(a[377] & b[71])^(a[376] & b[72])^(a[375] & b[73])^(a[374] & b[74])^(a[373] & b[75])^(a[372] & b[76])^(a[371] & b[77])^(a[370] & b[78])^(a[369] & b[79])^(a[368] & b[80])^(a[367] & b[81])^(a[366] & b[82])^(a[365] & b[83])^(a[364] & b[84])^(a[363] & b[85])^(a[362] & b[86])^(a[361] & b[87])^(a[360] & b[88])^(a[359] & b[89])^(a[358] & b[90])^(a[357] & b[91])^(a[356] & b[92])^(a[355] & b[93])^(a[354] & b[94])^(a[353] & b[95])^(a[352] & b[96])^(a[351] & b[97])^(a[350] & b[98])^(a[349] & b[99])^(a[348] & b[100])^(a[347] & b[101])^(a[346] & b[102])^(a[345] & b[103])^(a[344] & b[104])^(a[343] & b[105])^(a[342] & b[106])^(a[341] & b[107])^(a[340] & b[108])^(a[339] & b[109])^(a[338] & b[110])^(a[337] & b[111])^(a[336] & b[112])^(a[335] & b[113])^(a[334] & b[114])^(a[333] & b[115])^(a[332] & b[116])^(a[331] & b[117])^(a[330] & b[118])^(a[329] & b[119])^(a[328] & b[120])^(a[327] & b[121])^(a[326] & b[122])^(a[325] & b[123])^(a[324] & b[124])^(a[323] & b[125])^(a[322] & b[126])^(a[321] & b[127])^(a[320] & b[128])^(a[319] & b[129])^(a[318] & b[130])^(a[317] & b[131])^(a[316] & b[132])^(a[315] & b[133])^(a[314] & b[134])^(a[313] & b[135])^(a[312] & b[136])^(a[311] & b[137])^(a[310] & b[138])^(a[309] & b[139])^(a[308] & b[140])^(a[307] & b[141])^(a[306] & b[142])^(a[305] & b[143])^(a[304] & b[144])^(a[303] & b[145])^(a[302] & b[146])^(a[301] & b[147])^(a[300] & b[148])^(a[299] & b[149])^(a[298] & b[150])^(a[297] & b[151])^(a[296] & b[152])^(a[295] & b[153])^(a[294] & b[154])^(a[293] & b[155])^(a[292] & b[156])^(a[291] & b[157])^(a[290] & b[158])^(a[289] & b[159])^(a[288] & b[160])^(a[287] & b[161])^(a[286] & b[162])^(a[285] & b[163])^(a[284] & b[164])^(a[283] & b[165])^(a[282] & b[166])^(a[281] & b[167])^(a[280] & b[168])^(a[279] & b[169])^(a[278] & b[170])^(a[277] & b[171])^(a[276] & b[172])^(a[275] & b[173])^(a[274] & b[174])^(a[273] & b[175])^(a[272] & b[176])^(a[271] & b[177])^(a[270] & b[178])^(a[269] & b[179])^(a[268] & b[180])^(a[267] & b[181])^(a[266] & b[182])^(a[265] & b[183])^(a[264] & b[184])^(a[263] & b[185])^(a[262] & b[186])^(a[261] & b[187])^(a[260] & b[188])^(a[259] & b[189])^(a[258] & b[190])^(a[257] & b[191])^(a[256] & b[192])^(a[255] & b[193])^(a[254] & b[194])^(a[253] & b[195])^(a[252] & b[196])^(a[251] & b[197])^(a[250] & b[198])^(a[249] & b[199])^(a[248] & b[200])^(a[247] & b[201])^(a[246] & b[202])^(a[245] & b[203])^(a[244] & b[204])^(a[243] & b[205])^(a[242] & b[206])^(a[241] & b[207])^(a[240] & b[208])^(a[239] & b[209])^(a[238] & b[210])^(a[237] & b[211])^(a[236] & b[212])^(a[235] & b[213])^(a[234] & b[214])^(a[233] & b[215])^(a[232] & b[216])^(a[231] & b[217])^(a[230] & b[218])^(a[229] & b[219])^(a[228] & b[220])^(a[227] & b[221])^(a[226] & b[222])^(a[225] & b[223])^(a[224] & b[224])^(a[223] & b[225])^(a[222] & b[226])^(a[221] & b[227])^(a[220] & b[228])^(a[219] & b[229])^(a[218] & b[230])^(a[217] & b[231])^(a[216] & b[232])^(a[215] & b[233])^(a[214] & b[234])^(a[213] & b[235])^(a[212] & b[236])^(a[211] & b[237])^(a[210] & b[238])^(a[209] & b[239])^(a[208] & b[240])^(a[207] & b[241])^(a[206] & b[242])^(a[205] & b[243])^(a[204] & b[244])^(a[203] & b[245])^(a[202] & b[246])^(a[201] & b[247])^(a[200] & b[248])^(a[199] & b[249])^(a[198] & b[250])^(a[197] & b[251])^(a[196] & b[252])^(a[195] & b[253])^(a[194] & b[254])^(a[193] & b[255])^(a[192] & b[256])^(a[191] & b[257])^(a[190] & b[258])^(a[189] & b[259])^(a[188] & b[260])^(a[187] & b[261])^(a[186] & b[262])^(a[185] & b[263])^(a[184] & b[264])^(a[183] & b[265])^(a[182] & b[266])^(a[181] & b[267])^(a[180] & b[268])^(a[179] & b[269])^(a[178] & b[270])^(a[177] & b[271])^(a[176] & b[272])^(a[175] & b[273])^(a[174] & b[274])^(a[173] & b[275])^(a[172] & b[276])^(a[171] & b[277])^(a[170] & b[278])^(a[169] & b[279])^(a[168] & b[280])^(a[167] & b[281])^(a[166] & b[282])^(a[165] & b[283])^(a[164] & b[284])^(a[163] & b[285])^(a[162] & b[286])^(a[161] & b[287])^(a[160] & b[288])^(a[159] & b[289])^(a[158] & b[290])^(a[157] & b[291])^(a[156] & b[292])^(a[155] & b[293])^(a[154] & b[294])^(a[153] & b[295])^(a[152] & b[296])^(a[151] & b[297])^(a[150] & b[298])^(a[149] & b[299])^(a[148] & b[300])^(a[147] & b[301])^(a[146] & b[302])^(a[145] & b[303])^(a[144] & b[304])^(a[143] & b[305])^(a[142] & b[306])^(a[141] & b[307])^(a[140] & b[308])^(a[139] & b[309])^(a[138] & b[310])^(a[137] & b[311])^(a[136] & b[312])^(a[135] & b[313])^(a[134] & b[314])^(a[133] & b[315])^(a[132] & b[316])^(a[131] & b[317])^(a[130] & b[318])^(a[129] & b[319])^(a[128] & b[320])^(a[127] & b[321])^(a[126] & b[322])^(a[125] & b[323])^(a[124] & b[324])^(a[123] & b[325])^(a[122] & b[326])^(a[121] & b[327])^(a[120] & b[328])^(a[119] & b[329])^(a[118] & b[330])^(a[117] & b[331])^(a[116] & b[332])^(a[115] & b[333])^(a[114] & b[334])^(a[113] & b[335])^(a[112] & b[336])^(a[111] & b[337])^(a[110] & b[338])^(a[109] & b[339])^(a[108] & b[340])^(a[107] & b[341])^(a[106] & b[342])^(a[105] & b[343])^(a[104] & b[344])^(a[103] & b[345])^(a[102] & b[346])^(a[101] & b[347])^(a[100] & b[348])^(a[99] & b[349])^(a[98] & b[350])^(a[97] & b[351])^(a[96] & b[352])^(a[95] & b[353])^(a[94] & b[354])^(a[93] & b[355])^(a[92] & b[356])^(a[91] & b[357])^(a[90] & b[358])^(a[89] & b[359])^(a[88] & b[360])^(a[87] & b[361])^(a[86] & b[362])^(a[85] & b[363])^(a[84] & b[364])^(a[83] & b[365])^(a[82] & b[366])^(a[81] & b[367])^(a[80] & b[368])^(a[79] & b[369])^(a[78] & b[370])^(a[77] & b[371])^(a[76] & b[372])^(a[75] & b[373])^(a[74] & b[374])^(a[73] & b[375])^(a[72] & b[376])^(a[71] & b[377])^(a[70] & b[378])^(a[69] & b[379])^(a[68] & b[380])^(a[67] & b[381])^(a[66] & b[382])^(a[65] & b[383])^(a[64] & b[384])^(a[63] & b[385])^(a[62] & b[386])^(a[61] & b[387])^(a[60] & b[388])^(a[59] & b[389])^(a[58] & b[390])^(a[57] & b[391])^(a[56] & b[392])^(a[55] & b[393])^(a[54] & b[394])^(a[53] & b[395])^(a[52] & b[396])^(a[51] & b[397])^(a[50] & b[398])^(a[49] & b[399])^(a[48] & b[400])^(a[47] & b[401])^(a[46] & b[402])^(a[45] & b[403])^(a[44] & b[404])^(a[43] & b[405])^(a[42] & b[406])^(a[41] & b[407])^(a[40] & b[408]);
assign y[449] = (a[408] & b[41])^(a[407] & b[42])^(a[406] & b[43])^(a[405] & b[44])^(a[404] & b[45])^(a[403] & b[46])^(a[402] & b[47])^(a[401] & b[48])^(a[400] & b[49])^(a[399] & b[50])^(a[398] & b[51])^(a[397] & b[52])^(a[396] & b[53])^(a[395] & b[54])^(a[394] & b[55])^(a[393] & b[56])^(a[392] & b[57])^(a[391] & b[58])^(a[390] & b[59])^(a[389] & b[60])^(a[388] & b[61])^(a[387] & b[62])^(a[386] & b[63])^(a[385] & b[64])^(a[384] & b[65])^(a[383] & b[66])^(a[382] & b[67])^(a[381] & b[68])^(a[380] & b[69])^(a[379] & b[70])^(a[378] & b[71])^(a[377] & b[72])^(a[376] & b[73])^(a[375] & b[74])^(a[374] & b[75])^(a[373] & b[76])^(a[372] & b[77])^(a[371] & b[78])^(a[370] & b[79])^(a[369] & b[80])^(a[368] & b[81])^(a[367] & b[82])^(a[366] & b[83])^(a[365] & b[84])^(a[364] & b[85])^(a[363] & b[86])^(a[362] & b[87])^(a[361] & b[88])^(a[360] & b[89])^(a[359] & b[90])^(a[358] & b[91])^(a[357] & b[92])^(a[356] & b[93])^(a[355] & b[94])^(a[354] & b[95])^(a[353] & b[96])^(a[352] & b[97])^(a[351] & b[98])^(a[350] & b[99])^(a[349] & b[100])^(a[348] & b[101])^(a[347] & b[102])^(a[346] & b[103])^(a[345] & b[104])^(a[344] & b[105])^(a[343] & b[106])^(a[342] & b[107])^(a[341] & b[108])^(a[340] & b[109])^(a[339] & b[110])^(a[338] & b[111])^(a[337] & b[112])^(a[336] & b[113])^(a[335] & b[114])^(a[334] & b[115])^(a[333] & b[116])^(a[332] & b[117])^(a[331] & b[118])^(a[330] & b[119])^(a[329] & b[120])^(a[328] & b[121])^(a[327] & b[122])^(a[326] & b[123])^(a[325] & b[124])^(a[324] & b[125])^(a[323] & b[126])^(a[322] & b[127])^(a[321] & b[128])^(a[320] & b[129])^(a[319] & b[130])^(a[318] & b[131])^(a[317] & b[132])^(a[316] & b[133])^(a[315] & b[134])^(a[314] & b[135])^(a[313] & b[136])^(a[312] & b[137])^(a[311] & b[138])^(a[310] & b[139])^(a[309] & b[140])^(a[308] & b[141])^(a[307] & b[142])^(a[306] & b[143])^(a[305] & b[144])^(a[304] & b[145])^(a[303] & b[146])^(a[302] & b[147])^(a[301] & b[148])^(a[300] & b[149])^(a[299] & b[150])^(a[298] & b[151])^(a[297] & b[152])^(a[296] & b[153])^(a[295] & b[154])^(a[294] & b[155])^(a[293] & b[156])^(a[292] & b[157])^(a[291] & b[158])^(a[290] & b[159])^(a[289] & b[160])^(a[288] & b[161])^(a[287] & b[162])^(a[286] & b[163])^(a[285] & b[164])^(a[284] & b[165])^(a[283] & b[166])^(a[282] & b[167])^(a[281] & b[168])^(a[280] & b[169])^(a[279] & b[170])^(a[278] & b[171])^(a[277] & b[172])^(a[276] & b[173])^(a[275] & b[174])^(a[274] & b[175])^(a[273] & b[176])^(a[272] & b[177])^(a[271] & b[178])^(a[270] & b[179])^(a[269] & b[180])^(a[268] & b[181])^(a[267] & b[182])^(a[266] & b[183])^(a[265] & b[184])^(a[264] & b[185])^(a[263] & b[186])^(a[262] & b[187])^(a[261] & b[188])^(a[260] & b[189])^(a[259] & b[190])^(a[258] & b[191])^(a[257] & b[192])^(a[256] & b[193])^(a[255] & b[194])^(a[254] & b[195])^(a[253] & b[196])^(a[252] & b[197])^(a[251] & b[198])^(a[250] & b[199])^(a[249] & b[200])^(a[248] & b[201])^(a[247] & b[202])^(a[246] & b[203])^(a[245] & b[204])^(a[244] & b[205])^(a[243] & b[206])^(a[242] & b[207])^(a[241] & b[208])^(a[240] & b[209])^(a[239] & b[210])^(a[238] & b[211])^(a[237] & b[212])^(a[236] & b[213])^(a[235] & b[214])^(a[234] & b[215])^(a[233] & b[216])^(a[232] & b[217])^(a[231] & b[218])^(a[230] & b[219])^(a[229] & b[220])^(a[228] & b[221])^(a[227] & b[222])^(a[226] & b[223])^(a[225] & b[224])^(a[224] & b[225])^(a[223] & b[226])^(a[222] & b[227])^(a[221] & b[228])^(a[220] & b[229])^(a[219] & b[230])^(a[218] & b[231])^(a[217] & b[232])^(a[216] & b[233])^(a[215] & b[234])^(a[214] & b[235])^(a[213] & b[236])^(a[212] & b[237])^(a[211] & b[238])^(a[210] & b[239])^(a[209] & b[240])^(a[208] & b[241])^(a[207] & b[242])^(a[206] & b[243])^(a[205] & b[244])^(a[204] & b[245])^(a[203] & b[246])^(a[202] & b[247])^(a[201] & b[248])^(a[200] & b[249])^(a[199] & b[250])^(a[198] & b[251])^(a[197] & b[252])^(a[196] & b[253])^(a[195] & b[254])^(a[194] & b[255])^(a[193] & b[256])^(a[192] & b[257])^(a[191] & b[258])^(a[190] & b[259])^(a[189] & b[260])^(a[188] & b[261])^(a[187] & b[262])^(a[186] & b[263])^(a[185] & b[264])^(a[184] & b[265])^(a[183] & b[266])^(a[182] & b[267])^(a[181] & b[268])^(a[180] & b[269])^(a[179] & b[270])^(a[178] & b[271])^(a[177] & b[272])^(a[176] & b[273])^(a[175] & b[274])^(a[174] & b[275])^(a[173] & b[276])^(a[172] & b[277])^(a[171] & b[278])^(a[170] & b[279])^(a[169] & b[280])^(a[168] & b[281])^(a[167] & b[282])^(a[166] & b[283])^(a[165] & b[284])^(a[164] & b[285])^(a[163] & b[286])^(a[162] & b[287])^(a[161] & b[288])^(a[160] & b[289])^(a[159] & b[290])^(a[158] & b[291])^(a[157] & b[292])^(a[156] & b[293])^(a[155] & b[294])^(a[154] & b[295])^(a[153] & b[296])^(a[152] & b[297])^(a[151] & b[298])^(a[150] & b[299])^(a[149] & b[300])^(a[148] & b[301])^(a[147] & b[302])^(a[146] & b[303])^(a[145] & b[304])^(a[144] & b[305])^(a[143] & b[306])^(a[142] & b[307])^(a[141] & b[308])^(a[140] & b[309])^(a[139] & b[310])^(a[138] & b[311])^(a[137] & b[312])^(a[136] & b[313])^(a[135] & b[314])^(a[134] & b[315])^(a[133] & b[316])^(a[132] & b[317])^(a[131] & b[318])^(a[130] & b[319])^(a[129] & b[320])^(a[128] & b[321])^(a[127] & b[322])^(a[126] & b[323])^(a[125] & b[324])^(a[124] & b[325])^(a[123] & b[326])^(a[122] & b[327])^(a[121] & b[328])^(a[120] & b[329])^(a[119] & b[330])^(a[118] & b[331])^(a[117] & b[332])^(a[116] & b[333])^(a[115] & b[334])^(a[114] & b[335])^(a[113] & b[336])^(a[112] & b[337])^(a[111] & b[338])^(a[110] & b[339])^(a[109] & b[340])^(a[108] & b[341])^(a[107] & b[342])^(a[106] & b[343])^(a[105] & b[344])^(a[104] & b[345])^(a[103] & b[346])^(a[102] & b[347])^(a[101] & b[348])^(a[100] & b[349])^(a[99] & b[350])^(a[98] & b[351])^(a[97] & b[352])^(a[96] & b[353])^(a[95] & b[354])^(a[94] & b[355])^(a[93] & b[356])^(a[92] & b[357])^(a[91] & b[358])^(a[90] & b[359])^(a[89] & b[360])^(a[88] & b[361])^(a[87] & b[362])^(a[86] & b[363])^(a[85] & b[364])^(a[84] & b[365])^(a[83] & b[366])^(a[82] & b[367])^(a[81] & b[368])^(a[80] & b[369])^(a[79] & b[370])^(a[78] & b[371])^(a[77] & b[372])^(a[76] & b[373])^(a[75] & b[374])^(a[74] & b[375])^(a[73] & b[376])^(a[72] & b[377])^(a[71] & b[378])^(a[70] & b[379])^(a[69] & b[380])^(a[68] & b[381])^(a[67] & b[382])^(a[66] & b[383])^(a[65] & b[384])^(a[64] & b[385])^(a[63] & b[386])^(a[62] & b[387])^(a[61] & b[388])^(a[60] & b[389])^(a[59] & b[390])^(a[58] & b[391])^(a[57] & b[392])^(a[56] & b[393])^(a[55] & b[394])^(a[54] & b[395])^(a[53] & b[396])^(a[52] & b[397])^(a[51] & b[398])^(a[50] & b[399])^(a[49] & b[400])^(a[48] & b[401])^(a[47] & b[402])^(a[46] & b[403])^(a[45] & b[404])^(a[44] & b[405])^(a[43] & b[406])^(a[42] & b[407])^(a[41] & b[408]);
assign y[450] = (a[408] & b[42])^(a[407] & b[43])^(a[406] & b[44])^(a[405] & b[45])^(a[404] & b[46])^(a[403] & b[47])^(a[402] & b[48])^(a[401] & b[49])^(a[400] & b[50])^(a[399] & b[51])^(a[398] & b[52])^(a[397] & b[53])^(a[396] & b[54])^(a[395] & b[55])^(a[394] & b[56])^(a[393] & b[57])^(a[392] & b[58])^(a[391] & b[59])^(a[390] & b[60])^(a[389] & b[61])^(a[388] & b[62])^(a[387] & b[63])^(a[386] & b[64])^(a[385] & b[65])^(a[384] & b[66])^(a[383] & b[67])^(a[382] & b[68])^(a[381] & b[69])^(a[380] & b[70])^(a[379] & b[71])^(a[378] & b[72])^(a[377] & b[73])^(a[376] & b[74])^(a[375] & b[75])^(a[374] & b[76])^(a[373] & b[77])^(a[372] & b[78])^(a[371] & b[79])^(a[370] & b[80])^(a[369] & b[81])^(a[368] & b[82])^(a[367] & b[83])^(a[366] & b[84])^(a[365] & b[85])^(a[364] & b[86])^(a[363] & b[87])^(a[362] & b[88])^(a[361] & b[89])^(a[360] & b[90])^(a[359] & b[91])^(a[358] & b[92])^(a[357] & b[93])^(a[356] & b[94])^(a[355] & b[95])^(a[354] & b[96])^(a[353] & b[97])^(a[352] & b[98])^(a[351] & b[99])^(a[350] & b[100])^(a[349] & b[101])^(a[348] & b[102])^(a[347] & b[103])^(a[346] & b[104])^(a[345] & b[105])^(a[344] & b[106])^(a[343] & b[107])^(a[342] & b[108])^(a[341] & b[109])^(a[340] & b[110])^(a[339] & b[111])^(a[338] & b[112])^(a[337] & b[113])^(a[336] & b[114])^(a[335] & b[115])^(a[334] & b[116])^(a[333] & b[117])^(a[332] & b[118])^(a[331] & b[119])^(a[330] & b[120])^(a[329] & b[121])^(a[328] & b[122])^(a[327] & b[123])^(a[326] & b[124])^(a[325] & b[125])^(a[324] & b[126])^(a[323] & b[127])^(a[322] & b[128])^(a[321] & b[129])^(a[320] & b[130])^(a[319] & b[131])^(a[318] & b[132])^(a[317] & b[133])^(a[316] & b[134])^(a[315] & b[135])^(a[314] & b[136])^(a[313] & b[137])^(a[312] & b[138])^(a[311] & b[139])^(a[310] & b[140])^(a[309] & b[141])^(a[308] & b[142])^(a[307] & b[143])^(a[306] & b[144])^(a[305] & b[145])^(a[304] & b[146])^(a[303] & b[147])^(a[302] & b[148])^(a[301] & b[149])^(a[300] & b[150])^(a[299] & b[151])^(a[298] & b[152])^(a[297] & b[153])^(a[296] & b[154])^(a[295] & b[155])^(a[294] & b[156])^(a[293] & b[157])^(a[292] & b[158])^(a[291] & b[159])^(a[290] & b[160])^(a[289] & b[161])^(a[288] & b[162])^(a[287] & b[163])^(a[286] & b[164])^(a[285] & b[165])^(a[284] & b[166])^(a[283] & b[167])^(a[282] & b[168])^(a[281] & b[169])^(a[280] & b[170])^(a[279] & b[171])^(a[278] & b[172])^(a[277] & b[173])^(a[276] & b[174])^(a[275] & b[175])^(a[274] & b[176])^(a[273] & b[177])^(a[272] & b[178])^(a[271] & b[179])^(a[270] & b[180])^(a[269] & b[181])^(a[268] & b[182])^(a[267] & b[183])^(a[266] & b[184])^(a[265] & b[185])^(a[264] & b[186])^(a[263] & b[187])^(a[262] & b[188])^(a[261] & b[189])^(a[260] & b[190])^(a[259] & b[191])^(a[258] & b[192])^(a[257] & b[193])^(a[256] & b[194])^(a[255] & b[195])^(a[254] & b[196])^(a[253] & b[197])^(a[252] & b[198])^(a[251] & b[199])^(a[250] & b[200])^(a[249] & b[201])^(a[248] & b[202])^(a[247] & b[203])^(a[246] & b[204])^(a[245] & b[205])^(a[244] & b[206])^(a[243] & b[207])^(a[242] & b[208])^(a[241] & b[209])^(a[240] & b[210])^(a[239] & b[211])^(a[238] & b[212])^(a[237] & b[213])^(a[236] & b[214])^(a[235] & b[215])^(a[234] & b[216])^(a[233] & b[217])^(a[232] & b[218])^(a[231] & b[219])^(a[230] & b[220])^(a[229] & b[221])^(a[228] & b[222])^(a[227] & b[223])^(a[226] & b[224])^(a[225] & b[225])^(a[224] & b[226])^(a[223] & b[227])^(a[222] & b[228])^(a[221] & b[229])^(a[220] & b[230])^(a[219] & b[231])^(a[218] & b[232])^(a[217] & b[233])^(a[216] & b[234])^(a[215] & b[235])^(a[214] & b[236])^(a[213] & b[237])^(a[212] & b[238])^(a[211] & b[239])^(a[210] & b[240])^(a[209] & b[241])^(a[208] & b[242])^(a[207] & b[243])^(a[206] & b[244])^(a[205] & b[245])^(a[204] & b[246])^(a[203] & b[247])^(a[202] & b[248])^(a[201] & b[249])^(a[200] & b[250])^(a[199] & b[251])^(a[198] & b[252])^(a[197] & b[253])^(a[196] & b[254])^(a[195] & b[255])^(a[194] & b[256])^(a[193] & b[257])^(a[192] & b[258])^(a[191] & b[259])^(a[190] & b[260])^(a[189] & b[261])^(a[188] & b[262])^(a[187] & b[263])^(a[186] & b[264])^(a[185] & b[265])^(a[184] & b[266])^(a[183] & b[267])^(a[182] & b[268])^(a[181] & b[269])^(a[180] & b[270])^(a[179] & b[271])^(a[178] & b[272])^(a[177] & b[273])^(a[176] & b[274])^(a[175] & b[275])^(a[174] & b[276])^(a[173] & b[277])^(a[172] & b[278])^(a[171] & b[279])^(a[170] & b[280])^(a[169] & b[281])^(a[168] & b[282])^(a[167] & b[283])^(a[166] & b[284])^(a[165] & b[285])^(a[164] & b[286])^(a[163] & b[287])^(a[162] & b[288])^(a[161] & b[289])^(a[160] & b[290])^(a[159] & b[291])^(a[158] & b[292])^(a[157] & b[293])^(a[156] & b[294])^(a[155] & b[295])^(a[154] & b[296])^(a[153] & b[297])^(a[152] & b[298])^(a[151] & b[299])^(a[150] & b[300])^(a[149] & b[301])^(a[148] & b[302])^(a[147] & b[303])^(a[146] & b[304])^(a[145] & b[305])^(a[144] & b[306])^(a[143] & b[307])^(a[142] & b[308])^(a[141] & b[309])^(a[140] & b[310])^(a[139] & b[311])^(a[138] & b[312])^(a[137] & b[313])^(a[136] & b[314])^(a[135] & b[315])^(a[134] & b[316])^(a[133] & b[317])^(a[132] & b[318])^(a[131] & b[319])^(a[130] & b[320])^(a[129] & b[321])^(a[128] & b[322])^(a[127] & b[323])^(a[126] & b[324])^(a[125] & b[325])^(a[124] & b[326])^(a[123] & b[327])^(a[122] & b[328])^(a[121] & b[329])^(a[120] & b[330])^(a[119] & b[331])^(a[118] & b[332])^(a[117] & b[333])^(a[116] & b[334])^(a[115] & b[335])^(a[114] & b[336])^(a[113] & b[337])^(a[112] & b[338])^(a[111] & b[339])^(a[110] & b[340])^(a[109] & b[341])^(a[108] & b[342])^(a[107] & b[343])^(a[106] & b[344])^(a[105] & b[345])^(a[104] & b[346])^(a[103] & b[347])^(a[102] & b[348])^(a[101] & b[349])^(a[100] & b[350])^(a[99] & b[351])^(a[98] & b[352])^(a[97] & b[353])^(a[96] & b[354])^(a[95] & b[355])^(a[94] & b[356])^(a[93] & b[357])^(a[92] & b[358])^(a[91] & b[359])^(a[90] & b[360])^(a[89] & b[361])^(a[88] & b[362])^(a[87] & b[363])^(a[86] & b[364])^(a[85] & b[365])^(a[84] & b[366])^(a[83] & b[367])^(a[82] & b[368])^(a[81] & b[369])^(a[80] & b[370])^(a[79] & b[371])^(a[78] & b[372])^(a[77] & b[373])^(a[76] & b[374])^(a[75] & b[375])^(a[74] & b[376])^(a[73] & b[377])^(a[72] & b[378])^(a[71] & b[379])^(a[70] & b[380])^(a[69] & b[381])^(a[68] & b[382])^(a[67] & b[383])^(a[66] & b[384])^(a[65] & b[385])^(a[64] & b[386])^(a[63] & b[387])^(a[62] & b[388])^(a[61] & b[389])^(a[60] & b[390])^(a[59] & b[391])^(a[58] & b[392])^(a[57] & b[393])^(a[56] & b[394])^(a[55] & b[395])^(a[54] & b[396])^(a[53] & b[397])^(a[52] & b[398])^(a[51] & b[399])^(a[50] & b[400])^(a[49] & b[401])^(a[48] & b[402])^(a[47] & b[403])^(a[46] & b[404])^(a[45] & b[405])^(a[44] & b[406])^(a[43] & b[407])^(a[42] & b[408]);
assign y[451] = (a[408] & b[43])^(a[407] & b[44])^(a[406] & b[45])^(a[405] & b[46])^(a[404] & b[47])^(a[403] & b[48])^(a[402] & b[49])^(a[401] & b[50])^(a[400] & b[51])^(a[399] & b[52])^(a[398] & b[53])^(a[397] & b[54])^(a[396] & b[55])^(a[395] & b[56])^(a[394] & b[57])^(a[393] & b[58])^(a[392] & b[59])^(a[391] & b[60])^(a[390] & b[61])^(a[389] & b[62])^(a[388] & b[63])^(a[387] & b[64])^(a[386] & b[65])^(a[385] & b[66])^(a[384] & b[67])^(a[383] & b[68])^(a[382] & b[69])^(a[381] & b[70])^(a[380] & b[71])^(a[379] & b[72])^(a[378] & b[73])^(a[377] & b[74])^(a[376] & b[75])^(a[375] & b[76])^(a[374] & b[77])^(a[373] & b[78])^(a[372] & b[79])^(a[371] & b[80])^(a[370] & b[81])^(a[369] & b[82])^(a[368] & b[83])^(a[367] & b[84])^(a[366] & b[85])^(a[365] & b[86])^(a[364] & b[87])^(a[363] & b[88])^(a[362] & b[89])^(a[361] & b[90])^(a[360] & b[91])^(a[359] & b[92])^(a[358] & b[93])^(a[357] & b[94])^(a[356] & b[95])^(a[355] & b[96])^(a[354] & b[97])^(a[353] & b[98])^(a[352] & b[99])^(a[351] & b[100])^(a[350] & b[101])^(a[349] & b[102])^(a[348] & b[103])^(a[347] & b[104])^(a[346] & b[105])^(a[345] & b[106])^(a[344] & b[107])^(a[343] & b[108])^(a[342] & b[109])^(a[341] & b[110])^(a[340] & b[111])^(a[339] & b[112])^(a[338] & b[113])^(a[337] & b[114])^(a[336] & b[115])^(a[335] & b[116])^(a[334] & b[117])^(a[333] & b[118])^(a[332] & b[119])^(a[331] & b[120])^(a[330] & b[121])^(a[329] & b[122])^(a[328] & b[123])^(a[327] & b[124])^(a[326] & b[125])^(a[325] & b[126])^(a[324] & b[127])^(a[323] & b[128])^(a[322] & b[129])^(a[321] & b[130])^(a[320] & b[131])^(a[319] & b[132])^(a[318] & b[133])^(a[317] & b[134])^(a[316] & b[135])^(a[315] & b[136])^(a[314] & b[137])^(a[313] & b[138])^(a[312] & b[139])^(a[311] & b[140])^(a[310] & b[141])^(a[309] & b[142])^(a[308] & b[143])^(a[307] & b[144])^(a[306] & b[145])^(a[305] & b[146])^(a[304] & b[147])^(a[303] & b[148])^(a[302] & b[149])^(a[301] & b[150])^(a[300] & b[151])^(a[299] & b[152])^(a[298] & b[153])^(a[297] & b[154])^(a[296] & b[155])^(a[295] & b[156])^(a[294] & b[157])^(a[293] & b[158])^(a[292] & b[159])^(a[291] & b[160])^(a[290] & b[161])^(a[289] & b[162])^(a[288] & b[163])^(a[287] & b[164])^(a[286] & b[165])^(a[285] & b[166])^(a[284] & b[167])^(a[283] & b[168])^(a[282] & b[169])^(a[281] & b[170])^(a[280] & b[171])^(a[279] & b[172])^(a[278] & b[173])^(a[277] & b[174])^(a[276] & b[175])^(a[275] & b[176])^(a[274] & b[177])^(a[273] & b[178])^(a[272] & b[179])^(a[271] & b[180])^(a[270] & b[181])^(a[269] & b[182])^(a[268] & b[183])^(a[267] & b[184])^(a[266] & b[185])^(a[265] & b[186])^(a[264] & b[187])^(a[263] & b[188])^(a[262] & b[189])^(a[261] & b[190])^(a[260] & b[191])^(a[259] & b[192])^(a[258] & b[193])^(a[257] & b[194])^(a[256] & b[195])^(a[255] & b[196])^(a[254] & b[197])^(a[253] & b[198])^(a[252] & b[199])^(a[251] & b[200])^(a[250] & b[201])^(a[249] & b[202])^(a[248] & b[203])^(a[247] & b[204])^(a[246] & b[205])^(a[245] & b[206])^(a[244] & b[207])^(a[243] & b[208])^(a[242] & b[209])^(a[241] & b[210])^(a[240] & b[211])^(a[239] & b[212])^(a[238] & b[213])^(a[237] & b[214])^(a[236] & b[215])^(a[235] & b[216])^(a[234] & b[217])^(a[233] & b[218])^(a[232] & b[219])^(a[231] & b[220])^(a[230] & b[221])^(a[229] & b[222])^(a[228] & b[223])^(a[227] & b[224])^(a[226] & b[225])^(a[225] & b[226])^(a[224] & b[227])^(a[223] & b[228])^(a[222] & b[229])^(a[221] & b[230])^(a[220] & b[231])^(a[219] & b[232])^(a[218] & b[233])^(a[217] & b[234])^(a[216] & b[235])^(a[215] & b[236])^(a[214] & b[237])^(a[213] & b[238])^(a[212] & b[239])^(a[211] & b[240])^(a[210] & b[241])^(a[209] & b[242])^(a[208] & b[243])^(a[207] & b[244])^(a[206] & b[245])^(a[205] & b[246])^(a[204] & b[247])^(a[203] & b[248])^(a[202] & b[249])^(a[201] & b[250])^(a[200] & b[251])^(a[199] & b[252])^(a[198] & b[253])^(a[197] & b[254])^(a[196] & b[255])^(a[195] & b[256])^(a[194] & b[257])^(a[193] & b[258])^(a[192] & b[259])^(a[191] & b[260])^(a[190] & b[261])^(a[189] & b[262])^(a[188] & b[263])^(a[187] & b[264])^(a[186] & b[265])^(a[185] & b[266])^(a[184] & b[267])^(a[183] & b[268])^(a[182] & b[269])^(a[181] & b[270])^(a[180] & b[271])^(a[179] & b[272])^(a[178] & b[273])^(a[177] & b[274])^(a[176] & b[275])^(a[175] & b[276])^(a[174] & b[277])^(a[173] & b[278])^(a[172] & b[279])^(a[171] & b[280])^(a[170] & b[281])^(a[169] & b[282])^(a[168] & b[283])^(a[167] & b[284])^(a[166] & b[285])^(a[165] & b[286])^(a[164] & b[287])^(a[163] & b[288])^(a[162] & b[289])^(a[161] & b[290])^(a[160] & b[291])^(a[159] & b[292])^(a[158] & b[293])^(a[157] & b[294])^(a[156] & b[295])^(a[155] & b[296])^(a[154] & b[297])^(a[153] & b[298])^(a[152] & b[299])^(a[151] & b[300])^(a[150] & b[301])^(a[149] & b[302])^(a[148] & b[303])^(a[147] & b[304])^(a[146] & b[305])^(a[145] & b[306])^(a[144] & b[307])^(a[143] & b[308])^(a[142] & b[309])^(a[141] & b[310])^(a[140] & b[311])^(a[139] & b[312])^(a[138] & b[313])^(a[137] & b[314])^(a[136] & b[315])^(a[135] & b[316])^(a[134] & b[317])^(a[133] & b[318])^(a[132] & b[319])^(a[131] & b[320])^(a[130] & b[321])^(a[129] & b[322])^(a[128] & b[323])^(a[127] & b[324])^(a[126] & b[325])^(a[125] & b[326])^(a[124] & b[327])^(a[123] & b[328])^(a[122] & b[329])^(a[121] & b[330])^(a[120] & b[331])^(a[119] & b[332])^(a[118] & b[333])^(a[117] & b[334])^(a[116] & b[335])^(a[115] & b[336])^(a[114] & b[337])^(a[113] & b[338])^(a[112] & b[339])^(a[111] & b[340])^(a[110] & b[341])^(a[109] & b[342])^(a[108] & b[343])^(a[107] & b[344])^(a[106] & b[345])^(a[105] & b[346])^(a[104] & b[347])^(a[103] & b[348])^(a[102] & b[349])^(a[101] & b[350])^(a[100] & b[351])^(a[99] & b[352])^(a[98] & b[353])^(a[97] & b[354])^(a[96] & b[355])^(a[95] & b[356])^(a[94] & b[357])^(a[93] & b[358])^(a[92] & b[359])^(a[91] & b[360])^(a[90] & b[361])^(a[89] & b[362])^(a[88] & b[363])^(a[87] & b[364])^(a[86] & b[365])^(a[85] & b[366])^(a[84] & b[367])^(a[83] & b[368])^(a[82] & b[369])^(a[81] & b[370])^(a[80] & b[371])^(a[79] & b[372])^(a[78] & b[373])^(a[77] & b[374])^(a[76] & b[375])^(a[75] & b[376])^(a[74] & b[377])^(a[73] & b[378])^(a[72] & b[379])^(a[71] & b[380])^(a[70] & b[381])^(a[69] & b[382])^(a[68] & b[383])^(a[67] & b[384])^(a[66] & b[385])^(a[65] & b[386])^(a[64] & b[387])^(a[63] & b[388])^(a[62] & b[389])^(a[61] & b[390])^(a[60] & b[391])^(a[59] & b[392])^(a[58] & b[393])^(a[57] & b[394])^(a[56] & b[395])^(a[55] & b[396])^(a[54] & b[397])^(a[53] & b[398])^(a[52] & b[399])^(a[51] & b[400])^(a[50] & b[401])^(a[49] & b[402])^(a[48] & b[403])^(a[47] & b[404])^(a[46] & b[405])^(a[45] & b[406])^(a[44] & b[407])^(a[43] & b[408]);
assign y[452] = (a[408] & b[44])^(a[407] & b[45])^(a[406] & b[46])^(a[405] & b[47])^(a[404] & b[48])^(a[403] & b[49])^(a[402] & b[50])^(a[401] & b[51])^(a[400] & b[52])^(a[399] & b[53])^(a[398] & b[54])^(a[397] & b[55])^(a[396] & b[56])^(a[395] & b[57])^(a[394] & b[58])^(a[393] & b[59])^(a[392] & b[60])^(a[391] & b[61])^(a[390] & b[62])^(a[389] & b[63])^(a[388] & b[64])^(a[387] & b[65])^(a[386] & b[66])^(a[385] & b[67])^(a[384] & b[68])^(a[383] & b[69])^(a[382] & b[70])^(a[381] & b[71])^(a[380] & b[72])^(a[379] & b[73])^(a[378] & b[74])^(a[377] & b[75])^(a[376] & b[76])^(a[375] & b[77])^(a[374] & b[78])^(a[373] & b[79])^(a[372] & b[80])^(a[371] & b[81])^(a[370] & b[82])^(a[369] & b[83])^(a[368] & b[84])^(a[367] & b[85])^(a[366] & b[86])^(a[365] & b[87])^(a[364] & b[88])^(a[363] & b[89])^(a[362] & b[90])^(a[361] & b[91])^(a[360] & b[92])^(a[359] & b[93])^(a[358] & b[94])^(a[357] & b[95])^(a[356] & b[96])^(a[355] & b[97])^(a[354] & b[98])^(a[353] & b[99])^(a[352] & b[100])^(a[351] & b[101])^(a[350] & b[102])^(a[349] & b[103])^(a[348] & b[104])^(a[347] & b[105])^(a[346] & b[106])^(a[345] & b[107])^(a[344] & b[108])^(a[343] & b[109])^(a[342] & b[110])^(a[341] & b[111])^(a[340] & b[112])^(a[339] & b[113])^(a[338] & b[114])^(a[337] & b[115])^(a[336] & b[116])^(a[335] & b[117])^(a[334] & b[118])^(a[333] & b[119])^(a[332] & b[120])^(a[331] & b[121])^(a[330] & b[122])^(a[329] & b[123])^(a[328] & b[124])^(a[327] & b[125])^(a[326] & b[126])^(a[325] & b[127])^(a[324] & b[128])^(a[323] & b[129])^(a[322] & b[130])^(a[321] & b[131])^(a[320] & b[132])^(a[319] & b[133])^(a[318] & b[134])^(a[317] & b[135])^(a[316] & b[136])^(a[315] & b[137])^(a[314] & b[138])^(a[313] & b[139])^(a[312] & b[140])^(a[311] & b[141])^(a[310] & b[142])^(a[309] & b[143])^(a[308] & b[144])^(a[307] & b[145])^(a[306] & b[146])^(a[305] & b[147])^(a[304] & b[148])^(a[303] & b[149])^(a[302] & b[150])^(a[301] & b[151])^(a[300] & b[152])^(a[299] & b[153])^(a[298] & b[154])^(a[297] & b[155])^(a[296] & b[156])^(a[295] & b[157])^(a[294] & b[158])^(a[293] & b[159])^(a[292] & b[160])^(a[291] & b[161])^(a[290] & b[162])^(a[289] & b[163])^(a[288] & b[164])^(a[287] & b[165])^(a[286] & b[166])^(a[285] & b[167])^(a[284] & b[168])^(a[283] & b[169])^(a[282] & b[170])^(a[281] & b[171])^(a[280] & b[172])^(a[279] & b[173])^(a[278] & b[174])^(a[277] & b[175])^(a[276] & b[176])^(a[275] & b[177])^(a[274] & b[178])^(a[273] & b[179])^(a[272] & b[180])^(a[271] & b[181])^(a[270] & b[182])^(a[269] & b[183])^(a[268] & b[184])^(a[267] & b[185])^(a[266] & b[186])^(a[265] & b[187])^(a[264] & b[188])^(a[263] & b[189])^(a[262] & b[190])^(a[261] & b[191])^(a[260] & b[192])^(a[259] & b[193])^(a[258] & b[194])^(a[257] & b[195])^(a[256] & b[196])^(a[255] & b[197])^(a[254] & b[198])^(a[253] & b[199])^(a[252] & b[200])^(a[251] & b[201])^(a[250] & b[202])^(a[249] & b[203])^(a[248] & b[204])^(a[247] & b[205])^(a[246] & b[206])^(a[245] & b[207])^(a[244] & b[208])^(a[243] & b[209])^(a[242] & b[210])^(a[241] & b[211])^(a[240] & b[212])^(a[239] & b[213])^(a[238] & b[214])^(a[237] & b[215])^(a[236] & b[216])^(a[235] & b[217])^(a[234] & b[218])^(a[233] & b[219])^(a[232] & b[220])^(a[231] & b[221])^(a[230] & b[222])^(a[229] & b[223])^(a[228] & b[224])^(a[227] & b[225])^(a[226] & b[226])^(a[225] & b[227])^(a[224] & b[228])^(a[223] & b[229])^(a[222] & b[230])^(a[221] & b[231])^(a[220] & b[232])^(a[219] & b[233])^(a[218] & b[234])^(a[217] & b[235])^(a[216] & b[236])^(a[215] & b[237])^(a[214] & b[238])^(a[213] & b[239])^(a[212] & b[240])^(a[211] & b[241])^(a[210] & b[242])^(a[209] & b[243])^(a[208] & b[244])^(a[207] & b[245])^(a[206] & b[246])^(a[205] & b[247])^(a[204] & b[248])^(a[203] & b[249])^(a[202] & b[250])^(a[201] & b[251])^(a[200] & b[252])^(a[199] & b[253])^(a[198] & b[254])^(a[197] & b[255])^(a[196] & b[256])^(a[195] & b[257])^(a[194] & b[258])^(a[193] & b[259])^(a[192] & b[260])^(a[191] & b[261])^(a[190] & b[262])^(a[189] & b[263])^(a[188] & b[264])^(a[187] & b[265])^(a[186] & b[266])^(a[185] & b[267])^(a[184] & b[268])^(a[183] & b[269])^(a[182] & b[270])^(a[181] & b[271])^(a[180] & b[272])^(a[179] & b[273])^(a[178] & b[274])^(a[177] & b[275])^(a[176] & b[276])^(a[175] & b[277])^(a[174] & b[278])^(a[173] & b[279])^(a[172] & b[280])^(a[171] & b[281])^(a[170] & b[282])^(a[169] & b[283])^(a[168] & b[284])^(a[167] & b[285])^(a[166] & b[286])^(a[165] & b[287])^(a[164] & b[288])^(a[163] & b[289])^(a[162] & b[290])^(a[161] & b[291])^(a[160] & b[292])^(a[159] & b[293])^(a[158] & b[294])^(a[157] & b[295])^(a[156] & b[296])^(a[155] & b[297])^(a[154] & b[298])^(a[153] & b[299])^(a[152] & b[300])^(a[151] & b[301])^(a[150] & b[302])^(a[149] & b[303])^(a[148] & b[304])^(a[147] & b[305])^(a[146] & b[306])^(a[145] & b[307])^(a[144] & b[308])^(a[143] & b[309])^(a[142] & b[310])^(a[141] & b[311])^(a[140] & b[312])^(a[139] & b[313])^(a[138] & b[314])^(a[137] & b[315])^(a[136] & b[316])^(a[135] & b[317])^(a[134] & b[318])^(a[133] & b[319])^(a[132] & b[320])^(a[131] & b[321])^(a[130] & b[322])^(a[129] & b[323])^(a[128] & b[324])^(a[127] & b[325])^(a[126] & b[326])^(a[125] & b[327])^(a[124] & b[328])^(a[123] & b[329])^(a[122] & b[330])^(a[121] & b[331])^(a[120] & b[332])^(a[119] & b[333])^(a[118] & b[334])^(a[117] & b[335])^(a[116] & b[336])^(a[115] & b[337])^(a[114] & b[338])^(a[113] & b[339])^(a[112] & b[340])^(a[111] & b[341])^(a[110] & b[342])^(a[109] & b[343])^(a[108] & b[344])^(a[107] & b[345])^(a[106] & b[346])^(a[105] & b[347])^(a[104] & b[348])^(a[103] & b[349])^(a[102] & b[350])^(a[101] & b[351])^(a[100] & b[352])^(a[99] & b[353])^(a[98] & b[354])^(a[97] & b[355])^(a[96] & b[356])^(a[95] & b[357])^(a[94] & b[358])^(a[93] & b[359])^(a[92] & b[360])^(a[91] & b[361])^(a[90] & b[362])^(a[89] & b[363])^(a[88] & b[364])^(a[87] & b[365])^(a[86] & b[366])^(a[85] & b[367])^(a[84] & b[368])^(a[83] & b[369])^(a[82] & b[370])^(a[81] & b[371])^(a[80] & b[372])^(a[79] & b[373])^(a[78] & b[374])^(a[77] & b[375])^(a[76] & b[376])^(a[75] & b[377])^(a[74] & b[378])^(a[73] & b[379])^(a[72] & b[380])^(a[71] & b[381])^(a[70] & b[382])^(a[69] & b[383])^(a[68] & b[384])^(a[67] & b[385])^(a[66] & b[386])^(a[65] & b[387])^(a[64] & b[388])^(a[63] & b[389])^(a[62] & b[390])^(a[61] & b[391])^(a[60] & b[392])^(a[59] & b[393])^(a[58] & b[394])^(a[57] & b[395])^(a[56] & b[396])^(a[55] & b[397])^(a[54] & b[398])^(a[53] & b[399])^(a[52] & b[400])^(a[51] & b[401])^(a[50] & b[402])^(a[49] & b[403])^(a[48] & b[404])^(a[47] & b[405])^(a[46] & b[406])^(a[45] & b[407])^(a[44] & b[408]);
assign y[453] = (a[408] & b[45])^(a[407] & b[46])^(a[406] & b[47])^(a[405] & b[48])^(a[404] & b[49])^(a[403] & b[50])^(a[402] & b[51])^(a[401] & b[52])^(a[400] & b[53])^(a[399] & b[54])^(a[398] & b[55])^(a[397] & b[56])^(a[396] & b[57])^(a[395] & b[58])^(a[394] & b[59])^(a[393] & b[60])^(a[392] & b[61])^(a[391] & b[62])^(a[390] & b[63])^(a[389] & b[64])^(a[388] & b[65])^(a[387] & b[66])^(a[386] & b[67])^(a[385] & b[68])^(a[384] & b[69])^(a[383] & b[70])^(a[382] & b[71])^(a[381] & b[72])^(a[380] & b[73])^(a[379] & b[74])^(a[378] & b[75])^(a[377] & b[76])^(a[376] & b[77])^(a[375] & b[78])^(a[374] & b[79])^(a[373] & b[80])^(a[372] & b[81])^(a[371] & b[82])^(a[370] & b[83])^(a[369] & b[84])^(a[368] & b[85])^(a[367] & b[86])^(a[366] & b[87])^(a[365] & b[88])^(a[364] & b[89])^(a[363] & b[90])^(a[362] & b[91])^(a[361] & b[92])^(a[360] & b[93])^(a[359] & b[94])^(a[358] & b[95])^(a[357] & b[96])^(a[356] & b[97])^(a[355] & b[98])^(a[354] & b[99])^(a[353] & b[100])^(a[352] & b[101])^(a[351] & b[102])^(a[350] & b[103])^(a[349] & b[104])^(a[348] & b[105])^(a[347] & b[106])^(a[346] & b[107])^(a[345] & b[108])^(a[344] & b[109])^(a[343] & b[110])^(a[342] & b[111])^(a[341] & b[112])^(a[340] & b[113])^(a[339] & b[114])^(a[338] & b[115])^(a[337] & b[116])^(a[336] & b[117])^(a[335] & b[118])^(a[334] & b[119])^(a[333] & b[120])^(a[332] & b[121])^(a[331] & b[122])^(a[330] & b[123])^(a[329] & b[124])^(a[328] & b[125])^(a[327] & b[126])^(a[326] & b[127])^(a[325] & b[128])^(a[324] & b[129])^(a[323] & b[130])^(a[322] & b[131])^(a[321] & b[132])^(a[320] & b[133])^(a[319] & b[134])^(a[318] & b[135])^(a[317] & b[136])^(a[316] & b[137])^(a[315] & b[138])^(a[314] & b[139])^(a[313] & b[140])^(a[312] & b[141])^(a[311] & b[142])^(a[310] & b[143])^(a[309] & b[144])^(a[308] & b[145])^(a[307] & b[146])^(a[306] & b[147])^(a[305] & b[148])^(a[304] & b[149])^(a[303] & b[150])^(a[302] & b[151])^(a[301] & b[152])^(a[300] & b[153])^(a[299] & b[154])^(a[298] & b[155])^(a[297] & b[156])^(a[296] & b[157])^(a[295] & b[158])^(a[294] & b[159])^(a[293] & b[160])^(a[292] & b[161])^(a[291] & b[162])^(a[290] & b[163])^(a[289] & b[164])^(a[288] & b[165])^(a[287] & b[166])^(a[286] & b[167])^(a[285] & b[168])^(a[284] & b[169])^(a[283] & b[170])^(a[282] & b[171])^(a[281] & b[172])^(a[280] & b[173])^(a[279] & b[174])^(a[278] & b[175])^(a[277] & b[176])^(a[276] & b[177])^(a[275] & b[178])^(a[274] & b[179])^(a[273] & b[180])^(a[272] & b[181])^(a[271] & b[182])^(a[270] & b[183])^(a[269] & b[184])^(a[268] & b[185])^(a[267] & b[186])^(a[266] & b[187])^(a[265] & b[188])^(a[264] & b[189])^(a[263] & b[190])^(a[262] & b[191])^(a[261] & b[192])^(a[260] & b[193])^(a[259] & b[194])^(a[258] & b[195])^(a[257] & b[196])^(a[256] & b[197])^(a[255] & b[198])^(a[254] & b[199])^(a[253] & b[200])^(a[252] & b[201])^(a[251] & b[202])^(a[250] & b[203])^(a[249] & b[204])^(a[248] & b[205])^(a[247] & b[206])^(a[246] & b[207])^(a[245] & b[208])^(a[244] & b[209])^(a[243] & b[210])^(a[242] & b[211])^(a[241] & b[212])^(a[240] & b[213])^(a[239] & b[214])^(a[238] & b[215])^(a[237] & b[216])^(a[236] & b[217])^(a[235] & b[218])^(a[234] & b[219])^(a[233] & b[220])^(a[232] & b[221])^(a[231] & b[222])^(a[230] & b[223])^(a[229] & b[224])^(a[228] & b[225])^(a[227] & b[226])^(a[226] & b[227])^(a[225] & b[228])^(a[224] & b[229])^(a[223] & b[230])^(a[222] & b[231])^(a[221] & b[232])^(a[220] & b[233])^(a[219] & b[234])^(a[218] & b[235])^(a[217] & b[236])^(a[216] & b[237])^(a[215] & b[238])^(a[214] & b[239])^(a[213] & b[240])^(a[212] & b[241])^(a[211] & b[242])^(a[210] & b[243])^(a[209] & b[244])^(a[208] & b[245])^(a[207] & b[246])^(a[206] & b[247])^(a[205] & b[248])^(a[204] & b[249])^(a[203] & b[250])^(a[202] & b[251])^(a[201] & b[252])^(a[200] & b[253])^(a[199] & b[254])^(a[198] & b[255])^(a[197] & b[256])^(a[196] & b[257])^(a[195] & b[258])^(a[194] & b[259])^(a[193] & b[260])^(a[192] & b[261])^(a[191] & b[262])^(a[190] & b[263])^(a[189] & b[264])^(a[188] & b[265])^(a[187] & b[266])^(a[186] & b[267])^(a[185] & b[268])^(a[184] & b[269])^(a[183] & b[270])^(a[182] & b[271])^(a[181] & b[272])^(a[180] & b[273])^(a[179] & b[274])^(a[178] & b[275])^(a[177] & b[276])^(a[176] & b[277])^(a[175] & b[278])^(a[174] & b[279])^(a[173] & b[280])^(a[172] & b[281])^(a[171] & b[282])^(a[170] & b[283])^(a[169] & b[284])^(a[168] & b[285])^(a[167] & b[286])^(a[166] & b[287])^(a[165] & b[288])^(a[164] & b[289])^(a[163] & b[290])^(a[162] & b[291])^(a[161] & b[292])^(a[160] & b[293])^(a[159] & b[294])^(a[158] & b[295])^(a[157] & b[296])^(a[156] & b[297])^(a[155] & b[298])^(a[154] & b[299])^(a[153] & b[300])^(a[152] & b[301])^(a[151] & b[302])^(a[150] & b[303])^(a[149] & b[304])^(a[148] & b[305])^(a[147] & b[306])^(a[146] & b[307])^(a[145] & b[308])^(a[144] & b[309])^(a[143] & b[310])^(a[142] & b[311])^(a[141] & b[312])^(a[140] & b[313])^(a[139] & b[314])^(a[138] & b[315])^(a[137] & b[316])^(a[136] & b[317])^(a[135] & b[318])^(a[134] & b[319])^(a[133] & b[320])^(a[132] & b[321])^(a[131] & b[322])^(a[130] & b[323])^(a[129] & b[324])^(a[128] & b[325])^(a[127] & b[326])^(a[126] & b[327])^(a[125] & b[328])^(a[124] & b[329])^(a[123] & b[330])^(a[122] & b[331])^(a[121] & b[332])^(a[120] & b[333])^(a[119] & b[334])^(a[118] & b[335])^(a[117] & b[336])^(a[116] & b[337])^(a[115] & b[338])^(a[114] & b[339])^(a[113] & b[340])^(a[112] & b[341])^(a[111] & b[342])^(a[110] & b[343])^(a[109] & b[344])^(a[108] & b[345])^(a[107] & b[346])^(a[106] & b[347])^(a[105] & b[348])^(a[104] & b[349])^(a[103] & b[350])^(a[102] & b[351])^(a[101] & b[352])^(a[100] & b[353])^(a[99] & b[354])^(a[98] & b[355])^(a[97] & b[356])^(a[96] & b[357])^(a[95] & b[358])^(a[94] & b[359])^(a[93] & b[360])^(a[92] & b[361])^(a[91] & b[362])^(a[90] & b[363])^(a[89] & b[364])^(a[88] & b[365])^(a[87] & b[366])^(a[86] & b[367])^(a[85] & b[368])^(a[84] & b[369])^(a[83] & b[370])^(a[82] & b[371])^(a[81] & b[372])^(a[80] & b[373])^(a[79] & b[374])^(a[78] & b[375])^(a[77] & b[376])^(a[76] & b[377])^(a[75] & b[378])^(a[74] & b[379])^(a[73] & b[380])^(a[72] & b[381])^(a[71] & b[382])^(a[70] & b[383])^(a[69] & b[384])^(a[68] & b[385])^(a[67] & b[386])^(a[66] & b[387])^(a[65] & b[388])^(a[64] & b[389])^(a[63] & b[390])^(a[62] & b[391])^(a[61] & b[392])^(a[60] & b[393])^(a[59] & b[394])^(a[58] & b[395])^(a[57] & b[396])^(a[56] & b[397])^(a[55] & b[398])^(a[54] & b[399])^(a[53] & b[400])^(a[52] & b[401])^(a[51] & b[402])^(a[50] & b[403])^(a[49] & b[404])^(a[48] & b[405])^(a[47] & b[406])^(a[46] & b[407])^(a[45] & b[408]);
assign y[454] = (a[408] & b[46])^(a[407] & b[47])^(a[406] & b[48])^(a[405] & b[49])^(a[404] & b[50])^(a[403] & b[51])^(a[402] & b[52])^(a[401] & b[53])^(a[400] & b[54])^(a[399] & b[55])^(a[398] & b[56])^(a[397] & b[57])^(a[396] & b[58])^(a[395] & b[59])^(a[394] & b[60])^(a[393] & b[61])^(a[392] & b[62])^(a[391] & b[63])^(a[390] & b[64])^(a[389] & b[65])^(a[388] & b[66])^(a[387] & b[67])^(a[386] & b[68])^(a[385] & b[69])^(a[384] & b[70])^(a[383] & b[71])^(a[382] & b[72])^(a[381] & b[73])^(a[380] & b[74])^(a[379] & b[75])^(a[378] & b[76])^(a[377] & b[77])^(a[376] & b[78])^(a[375] & b[79])^(a[374] & b[80])^(a[373] & b[81])^(a[372] & b[82])^(a[371] & b[83])^(a[370] & b[84])^(a[369] & b[85])^(a[368] & b[86])^(a[367] & b[87])^(a[366] & b[88])^(a[365] & b[89])^(a[364] & b[90])^(a[363] & b[91])^(a[362] & b[92])^(a[361] & b[93])^(a[360] & b[94])^(a[359] & b[95])^(a[358] & b[96])^(a[357] & b[97])^(a[356] & b[98])^(a[355] & b[99])^(a[354] & b[100])^(a[353] & b[101])^(a[352] & b[102])^(a[351] & b[103])^(a[350] & b[104])^(a[349] & b[105])^(a[348] & b[106])^(a[347] & b[107])^(a[346] & b[108])^(a[345] & b[109])^(a[344] & b[110])^(a[343] & b[111])^(a[342] & b[112])^(a[341] & b[113])^(a[340] & b[114])^(a[339] & b[115])^(a[338] & b[116])^(a[337] & b[117])^(a[336] & b[118])^(a[335] & b[119])^(a[334] & b[120])^(a[333] & b[121])^(a[332] & b[122])^(a[331] & b[123])^(a[330] & b[124])^(a[329] & b[125])^(a[328] & b[126])^(a[327] & b[127])^(a[326] & b[128])^(a[325] & b[129])^(a[324] & b[130])^(a[323] & b[131])^(a[322] & b[132])^(a[321] & b[133])^(a[320] & b[134])^(a[319] & b[135])^(a[318] & b[136])^(a[317] & b[137])^(a[316] & b[138])^(a[315] & b[139])^(a[314] & b[140])^(a[313] & b[141])^(a[312] & b[142])^(a[311] & b[143])^(a[310] & b[144])^(a[309] & b[145])^(a[308] & b[146])^(a[307] & b[147])^(a[306] & b[148])^(a[305] & b[149])^(a[304] & b[150])^(a[303] & b[151])^(a[302] & b[152])^(a[301] & b[153])^(a[300] & b[154])^(a[299] & b[155])^(a[298] & b[156])^(a[297] & b[157])^(a[296] & b[158])^(a[295] & b[159])^(a[294] & b[160])^(a[293] & b[161])^(a[292] & b[162])^(a[291] & b[163])^(a[290] & b[164])^(a[289] & b[165])^(a[288] & b[166])^(a[287] & b[167])^(a[286] & b[168])^(a[285] & b[169])^(a[284] & b[170])^(a[283] & b[171])^(a[282] & b[172])^(a[281] & b[173])^(a[280] & b[174])^(a[279] & b[175])^(a[278] & b[176])^(a[277] & b[177])^(a[276] & b[178])^(a[275] & b[179])^(a[274] & b[180])^(a[273] & b[181])^(a[272] & b[182])^(a[271] & b[183])^(a[270] & b[184])^(a[269] & b[185])^(a[268] & b[186])^(a[267] & b[187])^(a[266] & b[188])^(a[265] & b[189])^(a[264] & b[190])^(a[263] & b[191])^(a[262] & b[192])^(a[261] & b[193])^(a[260] & b[194])^(a[259] & b[195])^(a[258] & b[196])^(a[257] & b[197])^(a[256] & b[198])^(a[255] & b[199])^(a[254] & b[200])^(a[253] & b[201])^(a[252] & b[202])^(a[251] & b[203])^(a[250] & b[204])^(a[249] & b[205])^(a[248] & b[206])^(a[247] & b[207])^(a[246] & b[208])^(a[245] & b[209])^(a[244] & b[210])^(a[243] & b[211])^(a[242] & b[212])^(a[241] & b[213])^(a[240] & b[214])^(a[239] & b[215])^(a[238] & b[216])^(a[237] & b[217])^(a[236] & b[218])^(a[235] & b[219])^(a[234] & b[220])^(a[233] & b[221])^(a[232] & b[222])^(a[231] & b[223])^(a[230] & b[224])^(a[229] & b[225])^(a[228] & b[226])^(a[227] & b[227])^(a[226] & b[228])^(a[225] & b[229])^(a[224] & b[230])^(a[223] & b[231])^(a[222] & b[232])^(a[221] & b[233])^(a[220] & b[234])^(a[219] & b[235])^(a[218] & b[236])^(a[217] & b[237])^(a[216] & b[238])^(a[215] & b[239])^(a[214] & b[240])^(a[213] & b[241])^(a[212] & b[242])^(a[211] & b[243])^(a[210] & b[244])^(a[209] & b[245])^(a[208] & b[246])^(a[207] & b[247])^(a[206] & b[248])^(a[205] & b[249])^(a[204] & b[250])^(a[203] & b[251])^(a[202] & b[252])^(a[201] & b[253])^(a[200] & b[254])^(a[199] & b[255])^(a[198] & b[256])^(a[197] & b[257])^(a[196] & b[258])^(a[195] & b[259])^(a[194] & b[260])^(a[193] & b[261])^(a[192] & b[262])^(a[191] & b[263])^(a[190] & b[264])^(a[189] & b[265])^(a[188] & b[266])^(a[187] & b[267])^(a[186] & b[268])^(a[185] & b[269])^(a[184] & b[270])^(a[183] & b[271])^(a[182] & b[272])^(a[181] & b[273])^(a[180] & b[274])^(a[179] & b[275])^(a[178] & b[276])^(a[177] & b[277])^(a[176] & b[278])^(a[175] & b[279])^(a[174] & b[280])^(a[173] & b[281])^(a[172] & b[282])^(a[171] & b[283])^(a[170] & b[284])^(a[169] & b[285])^(a[168] & b[286])^(a[167] & b[287])^(a[166] & b[288])^(a[165] & b[289])^(a[164] & b[290])^(a[163] & b[291])^(a[162] & b[292])^(a[161] & b[293])^(a[160] & b[294])^(a[159] & b[295])^(a[158] & b[296])^(a[157] & b[297])^(a[156] & b[298])^(a[155] & b[299])^(a[154] & b[300])^(a[153] & b[301])^(a[152] & b[302])^(a[151] & b[303])^(a[150] & b[304])^(a[149] & b[305])^(a[148] & b[306])^(a[147] & b[307])^(a[146] & b[308])^(a[145] & b[309])^(a[144] & b[310])^(a[143] & b[311])^(a[142] & b[312])^(a[141] & b[313])^(a[140] & b[314])^(a[139] & b[315])^(a[138] & b[316])^(a[137] & b[317])^(a[136] & b[318])^(a[135] & b[319])^(a[134] & b[320])^(a[133] & b[321])^(a[132] & b[322])^(a[131] & b[323])^(a[130] & b[324])^(a[129] & b[325])^(a[128] & b[326])^(a[127] & b[327])^(a[126] & b[328])^(a[125] & b[329])^(a[124] & b[330])^(a[123] & b[331])^(a[122] & b[332])^(a[121] & b[333])^(a[120] & b[334])^(a[119] & b[335])^(a[118] & b[336])^(a[117] & b[337])^(a[116] & b[338])^(a[115] & b[339])^(a[114] & b[340])^(a[113] & b[341])^(a[112] & b[342])^(a[111] & b[343])^(a[110] & b[344])^(a[109] & b[345])^(a[108] & b[346])^(a[107] & b[347])^(a[106] & b[348])^(a[105] & b[349])^(a[104] & b[350])^(a[103] & b[351])^(a[102] & b[352])^(a[101] & b[353])^(a[100] & b[354])^(a[99] & b[355])^(a[98] & b[356])^(a[97] & b[357])^(a[96] & b[358])^(a[95] & b[359])^(a[94] & b[360])^(a[93] & b[361])^(a[92] & b[362])^(a[91] & b[363])^(a[90] & b[364])^(a[89] & b[365])^(a[88] & b[366])^(a[87] & b[367])^(a[86] & b[368])^(a[85] & b[369])^(a[84] & b[370])^(a[83] & b[371])^(a[82] & b[372])^(a[81] & b[373])^(a[80] & b[374])^(a[79] & b[375])^(a[78] & b[376])^(a[77] & b[377])^(a[76] & b[378])^(a[75] & b[379])^(a[74] & b[380])^(a[73] & b[381])^(a[72] & b[382])^(a[71] & b[383])^(a[70] & b[384])^(a[69] & b[385])^(a[68] & b[386])^(a[67] & b[387])^(a[66] & b[388])^(a[65] & b[389])^(a[64] & b[390])^(a[63] & b[391])^(a[62] & b[392])^(a[61] & b[393])^(a[60] & b[394])^(a[59] & b[395])^(a[58] & b[396])^(a[57] & b[397])^(a[56] & b[398])^(a[55] & b[399])^(a[54] & b[400])^(a[53] & b[401])^(a[52] & b[402])^(a[51] & b[403])^(a[50] & b[404])^(a[49] & b[405])^(a[48] & b[406])^(a[47] & b[407])^(a[46] & b[408]);
assign y[455] = (a[408] & b[47])^(a[407] & b[48])^(a[406] & b[49])^(a[405] & b[50])^(a[404] & b[51])^(a[403] & b[52])^(a[402] & b[53])^(a[401] & b[54])^(a[400] & b[55])^(a[399] & b[56])^(a[398] & b[57])^(a[397] & b[58])^(a[396] & b[59])^(a[395] & b[60])^(a[394] & b[61])^(a[393] & b[62])^(a[392] & b[63])^(a[391] & b[64])^(a[390] & b[65])^(a[389] & b[66])^(a[388] & b[67])^(a[387] & b[68])^(a[386] & b[69])^(a[385] & b[70])^(a[384] & b[71])^(a[383] & b[72])^(a[382] & b[73])^(a[381] & b[74])^(a[380] & b[75])^(a[379] & b[76])^(a[378] & b[77])^(a[377] & b[78])^(a[376] & b[79])^(a[375] & b[80])^(a[374] & b[81])^(a[373] & b[82])^(a[372] & b[83])^(a[371] & b[84])^(a[370] & b[85])^(a[369] & b[86])^(a[368] & b[87])^(a[367] & b[88])^(a[366] & b[89])^(a[365] & b[90])^(a[364] & b[91])^(a[363] & b[92])^(a[362] & b[93])^(a[361] & b[94])^(a[360] & b[95])^(a[359] & b[96])^(a[358] & b[97])^(a[357] & b[98])^(a[356] & b[99])^(a[355] & b[100])^(a[354] & b[101])^(a[353] & b[102])^(a[352] & b[103])^(a[351] & b[104])^(a[350] & b[105])^(a[349] & b[106])^(a[348] & b[107])^(a[347] & b[108])^(a[346] & b[109])^(a[345] & b[110])^(a[344] & b[111])^(a[343] & b[112])^(a[342] & b[113])^(a[341] & b[114])^(a[340] & b[115])^(a[339] & b[116])^(a[338] & b[117])^(a[337] & b[118])^(a[336] & b[119])^(a[335] & b[120])^(a[334] & b[121])^(a[333] & b[122])^(a[332] & b[123])^(a[331] & b[124])^(a[330] & b[125])^(a[329] & b[126])^(a[328] & b[127])^(a[327] & b[128])^(a[326] & b[129])^(a[325] & b[130])^(a[324] & b[131])^(a[323] & b[132])^(a[322] & b[133])^(a[321] & b[134])^(a[320] & b[135])^(a[319] & b[136])^(a[318] & b[137])^(a[317] & b[138])^(a[316] & b[139])^(a[315] & b[140])^(a[314] & b[141])^(a[313] & b[142])^(a[312] & b[143])^(a[311] & b[144])^(a[310] & b[145])^(a[309] & b[146])^(a[308] & b[147])^(a[307] & b[148])^(a[306] & b[149])^(a[305] & b[150])^(a[304] & b[151])^(a[303] & b[152])^(a[302] & b[153])^(a[301] & b[154])^(a[300] & b[155])^(a[299] & b[156])^(a[298] & b[157])^(a[297] & b[158])^(a[296] & b[159])^(a[295] & b[160])^(a[294] & b[161])^(a[293] & b[162])^(a[292] & b[163])^(a[291] & b[164])^(a[290] & b[165])^(a[289] & b[166])^(a[288] & b[167])^(a[287] & b[168])^(a[286] & b[169])^(a[285] & b[170])^(a[284] & b[171])^(a[283] & b[172])^(a[282] & b[173])^(a[281] & b[174])^(a[280] & b[175])^(a[279] & b[176])^(a[278] & b[177])^(a[277] & b[178])^(a[276] & b[179])^(a[275] & b[180])^(a[274] & b[181])^(a[273] & b[182])^(a[272] & b[183])^(a[271] & b[184])^(a[270] & b[185])^(a[269] & b[186])^(a[268] & b[187])^(a[267] & b[188])^(a[266] & b[189])^(a[265] & b[190])^(a[264] & b[191])^(a[263] & b[192])^(a[262] & b[193])^(a[261] & b[194])^(a[260] & b[195])^(a[259] & b[196])^(a[258] & b[197])^(a[257] & b[198])^(a[256] & b[199])^(a[255] & b[200])^(a[254] & b[201])^(a[253] & b[202])^(a[252] & b[203])^(a[251] & b[204])^(a[250] & b[205])^(a[249] & b[206])^(a[248] & b[207])^(a[247] & b[208])^(a[246] & b[209])^(a[245] & b[210])^(a[244] & b[211])^(a[243] & b[212])^(a[242] & b[213])^(a[241] & b[214])^(a[240] & b[215])^(a[239] & b[216])^(a[238] & b[217])^(a[237] & b[218])^(a[236] & b[219])^(a[235] & b[220])^(a[234] & b[221])^(a[233] & b[222])^(a[232] & b[223])^(a[231] & b[224])^(a[230] & b[225])^(a[229] & b[226])^(a[228] & b[227])^(a[227] & b[228])^(a[226] & b[229])^(a[225] & b[230])^(a[224] & b[231])^(a[223] & b[232])^(a[222] & b[233])^(a[221] & b[234])^(a[220] & b[235])^(a[219] & b[236])^(a[218] & b[237])^(a[217] & b[238])^(a[216] & b[239])^(a[215] & b[240])^(a[214] & b[241])^(a[213] & b[242])^(a[212] & b[243])^(a[211] & b[244])^(a[210] & b[245])^(a[209] & b[246])^(a[208] & b[247])^(a[207] & b[248])^(a[206] & b[249])^(a[205] & b[250])^(a[204] & b[251])^(a[203] & b[252])^(a[202] & b[253])^(a[201] & b[254])^(a[200] & b[255])^(a[199] & b[256])^(a[198] & b[257])^(a[197] & b[258])^(a[196] & b[259])^(a[195] & b[260])^(a[194] & b[261])^(a[193] & b[262])^(a[192] & b[263])^(a[191] & b[264])^(a[190] & b[265])^(a[189] & b[266])^(a[188] & b[267])^(a[187] & b[268])^(a[186] & b[269])^(a[185] & b[270])^(a[184] & b[271])^(a[183] & b[272])^(a[182] & b[273])^(a[181] & b[274])^(a[180] & b[275])^(a[179] & b[276])^(a[178] & b[277])^(a[177] & b[278])^(a[176] & b[279])^(a[175] & b[280])^(a[174] & b[281])^(a[173] & b[282])^(a[172] & b[283])^(a[171] & b[284])^(a[170] & b[285])^(a[169] & b[286])^(a[168] & b[287])^(a[167] & b[288])^(a[166] & b[289])^(a[165] & b[290])^(a[164] & b[291])^(a[163] & b[292])^(a[162] & b[293])^(a[161] & b[294])^(a[160] & b[295])^(a[159] & b[296])^(a[158] & b[297])^(a[157] & b[298])^(a[156] & b[299])^(a[155] & b[300])^(a[154] & b[301])^(a[153] & b[302])^(a[152] & b[303])^(a[151] & b[304])^(a[150] & b[305])^(a[149] & b[306])^(a[148] & b[307])^(a[147] & b[308])^(a[146] & b[309])^(a[145] & b[310])^(a[144] & b[311])^(a[143] & b[312])^(a[142] & b[313])^(a[141] & b[314])^(a[140] & b[315])^(a[139] & b[316])^(a[138] & b[317])^(a[137] & b[318])^(a[136] & b[319])^(a[135] & b[320])^(a[134] & b[321])^(a[133] & b[322])^(a[132] & b[323])^(a[131] & b[324])^(a[130] & b[325])^(a[129] & b[326])^(a[128] & b[327])^(a[127] & b[328])^(a[126] & b[329])^(a[125] & b[330])^(a[124] & b[331])^(a[123] & b[332])^(a[122] & b[333])^(a[121] & b[334])^(a[120] & b[335])^(a[119] & b[336])^(a[118] & b[337])^(a[117] & b[338])^(a[116] & b[339])^(a[115] & b[340])^(a[114] & b[341])^(a[113] & b[342])^(a[112] & b[343])^(a[111] & b[344])^(a[110] & b[345])^(a[109] & b[346])^(a[108] & b[347])^(a[107] & b[348])^(a[106] & b[349])^(a[105] & b[350])^(a[104] & b[351])^(a[103] & b[352])^(a[102] & b[353])^(a[101] & b[354])^(a[100] & b[355])^(a[99] & b[356])^(a[98] & b[357])^(a[97] & b[358])^(a[96] & b[359])^(a[95] & b[360])^(a[94] & b[361])^(a[93] & b[362])^(a[92] & b[363])^(a[91] & b[364])^(a[90] & b[365])^(a[89] & b[366])^(a[88] & b[367])^(a[87] & b[368])^(a[86] & b[369])^(a[85] & b[370])^(a[84] & b[371])^(a[83] & b[372])^(a[82] & b[373])^(a[81] & b[374])^(a[80] & b[375])^(a[79] & b[376])^(a[78] & b[377])^(a[77] & b[378])^(a[76] & b[379])^(a[75] & b[380])^(a[74] & b[381])^(a[73] & b[382])^(a[72] & b[383])^(a[71] & b[384])^(a[70] & b[385])^(a[69] & b[386])^(a[68] & b[387])^(a[67] & b[388])^(a[66] & b[389])^(a[65] & b[390])^(a[64] & b[391])^(a[63] & b[392])^(a[62] & b[393])^(a[61] & b[394])^(a[60] & b[395])^(a[59] & b[396])^(a[58] & b[397])^(a[57] & b[398])^(a[56] & b[399])^(a[55] & b[400])^(a[54] & b[401])^(a[53] & b[402])^(a[52] & b[403])^(a[51] & b[404])^(a[50] & b[405])^(a[49] & b[406])^(a[48] & b[407])^(a[47] & b[408]);
assign y[456] = (a[408] & b[48])^(a[407] & b[49])^(a[406] & b[50])^(a[405] & b[51])^(a[404] & b[52])^(a[403] & b[53])^(a[402] & b[54])^(a[401] & b[55])^(a[400] & b[56])^(a[399] & b[57])^(a[398] & b[58])^(a[397] & b[59])^(a[396] & b[60])^(a[395] & b[61])^(a[394] & b[62])^(a[393] & b[63])^(a[392] & b[64])^(a[391] & b[65])^(a[390] & b[66])^(a[389] & b[67])^(a[388] & b[68])^(a[387] & b[69])^(a[386] & b[70])^(a[385] & b[71])^(a[384] & b[72])^(a[383] & b[73])^(a[382] & b[74])^(a[381] & b[75])^(a[380] & b[76])^(a[379] & b[77])^(a[378] & b[78])^(a[377] & b[79])^(a[376] & b[80])^(a[375] & b[81])^(a[374] & b[82])^(a[373] & b[83])^(a[372] & b[84])^(a[371] & b[85])^(a[370] & b[86])^(a[369] & b[87])^(a[368] & b[88])^(a[367] & b[89])^(a[366] & b[90])^(a[365] & b[91])^(a[364] & b[92])^(a[363] & b[93])^(a[362] & b[94])^(a[361] & b[95])^(a[360] & b[96])^(a[359] & b[97])^(a[358] & b[98])^(a[357] & b[99])^(a[356] & b[100])^(a[355] & b[101])^(a[354] & b[102])^(a[353] & b[103])^(a[352] & b[104])^(a[351] & b[105])^(a[350] & b[106])^(a[349] & b[107])^(a[348] & b[108])^(a[347] & b[109])^(a[346] & b[110])^(a[345] & b[111])^(a[344] & b[112])^(a[343] & b[113])^(a[342] & b[114])^(a[341] & b[115])^(a[340] & b[116])^(a[339] & b[117])^(a[338] & b[118])^(a[337] & b[119])^(a[336] & b[120])^(a[335] & b[121])^(a[334] & b[122])^(a[333] & b[123])^(a[332] & b[124])^(a[331] & b[125])^(a[330] & b[126])^(a[329] & b[127])^(a[328] & b[128])^(a[327] & b[129])^(a[326] & b[130])^(a[325] & b[131])^(a[324] & b[132])^(a[323] & b[133])^(a[322] & b[134])^(a[321] & b[135])^(a[320] & b[136])^(a[319] & b[137])^(a[318] & b[138])^(a[317] & b[139])^(a[316] & b[140])^(a[315] & b[141])^(a[314] & b[142])^(a[313] & b[143])^(a[312] & b[144])^(a[311] & b[145])^(a[310] & b[146])^(a[309] & b[147])^(a[308] & b[148])^(a[307] & b[149])^(a[306] & b[150])^(a[305] & b[151])^(a[304] & b[152])^(a[303] & b[153])^(a[302] & b[154])^(a[301] & b[155])^(a[300] & b[156])^(a[299] & b[157])^(a[298] & b[158])^(a[297] & b[159])^(a[296] & b[160])^(a[295] & b[161])^(a[294] & b[162])^(a[293] & b[163])^(a[292] & b[164])^(a[291] & b[165])^(a[290] & b[166])^(a[289] & b[167])^(a[288] & b[168])^(a[287] & b[169])^(a[286] & b[170])^(a[285] & b[171])^(a[284] & b[172])^(a[283] & b[173])^(a[282] & b[174])^(a[281] & b[175])^(a[280] & b[176])^(a[279] & b[177])^(a[278] & b[178])^(a[277] & b[179])^(a[276] & b[180])^(a[275] & b[181])^(a[274] & b[182])^(a[273] & b[183])^(a[272] & b[184])^(a[271] & b[185])^(a[270] & b[186])^(a[269] & b[187])^(a[268] & b[188])^(a[267] & b[189])^(a[266] & b[190])^(a[265] & b[191])^(a[264] & b[192])^(a[263] & b[193])^(a[262] & b[194])^(a[261] & b[195])^(a[260] & b[196])^(a[259] & b[197])^(a[258] & b[198])^(a[257] & b[199])^(a[256] & b[200])^(a[255] & b[201])^(a[254] & b[202])^(a[253] & b[203])^(a[252] & b[204])^(a[251] & b[205])^(a[250] & b[206])^(a[249] & b[207])^(a[248] & b[208])^(a[247] & b[209])^(a[246] & b[210])^(a[245] & b[211])^(a[244] & b[212])^(a[243] & b[213])^(a[242] & b[214])^(a[241] & b[215])^(a[240] & b[216])^(a[239] & b[217])^(a[238] & b[218])^(a[237] & b[219])^(a[236] & b[220])^(a[235] & b[221])^(a[234] & b[222])^(a[233] & b[223])^(a[232] & b[224])^(a[231] & b[225])^(a[230] & b[226])^(a[229] & b[227])^(a[228] & b[228])^(a[227] & b[229])^(a[226] & b[230])^(a[225] & b[231])^(a[224] & b[232])^(a[223] & b[233])^(a[222] & b[234])^(a[221] & b[235])^(a[220] & b[236])^(a[219] & b[237])^(a[218] & b[238])^(a[217] & b[239])^(a[216] & b[240])^(a[215] & b[241])^(a[214] & b[242])^(a[213] & b[243])^(a[212] & b[244])^(a[211] & b[245])^(a[210] & b[246])^(a[209] & b[247])^(a[208] & b[248])^(a[207] & b[249])^(a[206] & b[250])^(a[205] & b[251])^(a[204] & b[252])^(a[203] & b[253])^(a[202] & b[254])^(a[201] & b[255])^(a[200] & b[256])^(a[199] & b[257])^(a[198] & b[258])^(a[197] & b[259])^(a[196] & b[260])^(a[195] & b[261])^(a[194] & b[262])^(a[193] & b[263])^(a[192] & b[264])^(a[191] & b[265])^(a[190] & b[266])^(a[189] & b[267])^(a[188] & b[268])^(a[187] & b[269])^(a[186] & b[270])^(a[185] & b[271])^(a[184] & b[272])^(a[183] & b[273])^(a[182] & b[274])^(a[181] & b[275])^(a[180] & b[276])^(a[179] & b[277])^(a[178] & b[278])^(a[177] & b[279])^(a[176] & b[280])^(a[175] & b[281])^(a[174] & b[282])^(a[173] & b[283])^(a[172] & b[284])^(a[171] & b[285])^(a[170] & b[286])^(a[169] & b[287])^(a[168] & b[288])^(a[167] & b[289])^(a[166] & b[290])^(a[165] & b[291])^(a[164] & b[292])^(a[163] & b[293])^(a[162] & b[294])^(a[161] & b[295])^(a[160] & b[296])^(a[159] & b[297])^(a[158] & b[298])^(a[157] & b[299])^(a[156] & b[300])^(a[155] & b[301])^(a[154] & b[302])^(a[153] & b[303])^(a[152] & b[304])^(a[151] & b[305])^(a[150] & b[306])^(a[149] & b[307])^(a[148] & b[308])^(a[147] & b[309])^(a[146] & b[310])^(a[145] & b[311])^(a[144] & b[312])^(a[143] & b[313])^(a[142] & b[314])^(a[141] & b[315])^(a[140] & b[316])^(a[139] & b[317])^(a[138] & b[318])^(a[137] & b[319])^(a[136] & b[320])^(a[135] & b[321])^(a[134] & b[322])^(a[133] & b[323])^(a[132] & b[324])^(a[131] & b[325])^(a[130] & b[326])^(a[129] & b[327])^(a[128] & b[328])^(a[127] & b[329])^(a[126] & b[330])^(a[125] & b[331])^(a[124] & b[332])^(a[123] & b[333])^(a[122] & b[334])^(a[121] & b[335])^(a[120] & b[336])^(a[119] & b[337])^(a[118] & b[338])^(a[117] & b[339])^(a[116] & b[340])^(a[115] & b[341])^(a[114] & b[342])^(a[113] & b[343])^(a[112] & b[344])^(a[111] & b[345])^(a[110] & b[346])^(a[109] & b[347])^(a[108] & b[348])^(a[107] & b[349])^(a[106] & b[350])^(a[105] & b[351])^(a[104] & b[352])^(a[103] & b[353])^(a[102] & b[354])^(a[101] & b[355])^(a[100] & b[356])^(a[99] & b[357])^(a[98] & b[358])^(a[97] & b[359])^(a[96] & b[360])^(a[95] & b[361])^(a[94] & b[362])^(a[93] & b[363])^(a[92] & b[364])^(a[91] & b[365])^(a[90] & b[366])^(a[89] & b[367])^(a[88] & b[368])^(a[87] & b[369])^(a[86] & b[370])^(a[85] & b[371])^(a[84] & b[372])^(a[83] & b[373])^(a[82] & b[374])^(a[81] & b[375])^(a[80] & b[376])^(a[79] & b[377])^(a[78] & b[378])^(a[77] & b[379])^(a[76] & b[380])^(a[75] & b[381])^(a[74] & b[382])^(a[73] & b[383])^(a[72] & b[384])^(a[71] & b[385])^(a[70] & b[386])^(a[69] & b[387])^(a[68] & b[388])^(a[67] & b[389])^(a[66] & b[390])^(a[65] & b[391])^(a[64] & b[392])^(a[63] & b[393])^(a[62] & b[394])^(a[61] & b[395])^(a[60] & b[396])^(a[59] & b[397])^(a[58] & b[398])^(a[57] & b[399])^(a[56] & b[400])^(a[55] & b[401])^(a[54] & b[402])^(a[53] & b[403])^(a[52] & b[404])^(a[51] & b[405])^(a[50] & b[406])^(a[49] & b[407])^(a[48] & b[408]);
assign y[457] = (a[408] & b[49])^(a[407] & b[50])^(a[406] & b[51])^(a[405] & b[52])^(a[404] & b[53])^(a[403] & b[54])^(a[402] & b[55])^(a[401] & b[56])^(a[400] & b[57])^(a[399] & b[58])^(a[398] & b[59])^(a[397] & b[60])^(a[396] & b[61])^(a[395] & b[62])^(a[394] & b[63])^(a[393] & b[64])^(a[392] & b[65])^(a[391] & b[66])^(a[390] & b[67])^(a[389] & b[68])^(a[388] & b[69])^(a[387] & b[70])^(a[386] & b[71])^(a[385] & b[72])^(a[384] & b[73])^(a[383] & b[74])^(a[382] & b[75])^(a[381] & b[76])^(a[380] & b[77])^(a[379] & b[78])^(a[378] & b[79])^(a[377] & b[80])^(a[376] & b[81])^(a[375] & b[82])^(a[374] & b[83])^(a[373] & b[84])^(a[372] & b[85])^(a[371] & b[86])^(a[370] & b[87])^(a[369] & b[88])^(a[368] & b[89])^(a[367] & b[90])^(a[366] & b[91])^(a[365] & b[92])^(a[364] & b[93])^(a[363] & b[94])^(a[362] & b[95])^(a[361] & b[96])^(a[360] & b[97])^(a[359] & b[98])^(a[358] & b[99])^(a[357] & b[100])^(a[356] & b[101])^(a[355] & b[102])^(a[354] & b[103])^(a[353] & b[104])^(a[352] & b[105])^(a[351] & b[106])^(a[350] & b[107])^(a[349] & b[108])^(a[348] & b[109])^(a[347] & b[110])^(a[346] & b[111])^(a[345] & b[112])^(a[344] & b[113])^(a[343] & b[114])^(a[342] & b[115])^(a[341] & b[116])^(a[340] & b[117])^(a[339] & b[118])^(a[338] & b[119])^(a[337] & b[120])^(a[336] & b[121])^(a[335] & b[122])^(a[334] & b[123])^(a[333] & b[124])^(a[332] & b[125])^(a[331] & b[126])^(a[330] & b[127])^(a[329] & b[128])^(a[328] & b[129])^(a[327] & b[130])^(a[326] & b[131])^(a[325] & b[132])^(a[324] & b[133])^(a[323] & b[134])^(a[322] & b[135])^(a[321] & b[136])^(a[320] & b[137])^(a[319] & b[138])^(a[318] & b[139])^(a[317] & b[140])^(a[316] & b[141])^(a[315] & b[142])^(a[314] & b[143])^(a[313] & b[144])^(a[312] & b[145])^(a[311] & b[146])^(a[310] & b[147])^(a[309] & b[148])^(a[308] & b[149])^(a[307] & b[150])^(a[306] & b[151])^(a[305] & b[152])^(a[304] & b[153])^(a[303] & b[154])^(a[302] & b[155])^(a[301] & b[156])^(a[300] & b[157])^(a[299] & b[158])^(a[298] & b[159])^(a[297] & b[160])^(a[296] & b[161])^(a[295] & b[162])^(a[294] & b[163])^(a[293] & b[164])^(a[292] & b[165])^(a[291] & b[166])^(a[290] & b[167])^(a[289] & b[168])^(a[288] & b[169])^(a[287] & b[170])^(a[286] & b[171])^(a[285] & b[172])^(a[284] & b[173])^(a[283] & b[174])^(a[282] & b[175])^(a[281] & b[176])^(a[280] & b[177])^(a[279] & b[178])^(a[278] & b[179])^(a[277] & b[180])^(a[276] & b[181])^(a[275] & b[182])^(a[274] & b[183])^(a[273] & b[184])^(a[272] & b[185])^(a[271] & b[186])^(a[270] & b[187])^(a[269] & b[188])^(a[268] & b[189])^(a[267] & b[190])^(a[266] & b[191])^(a[265] & b[192])^(a[264] & b[193])^(a[263] & b[194])^(a[262] & b[195])^(a[261] & b[196])^(a[260] & b[197])^(a[259] & b[198])^(a[258] & b[199])^(a[257] & b[200])^(a[256] & b[201])^(a[255] & b[202])^(a[254] & b[203])^(a[253] & b[204])^(a[252] & b[205])^(a[251] & b[206])^(a[250] & b[207])^(a[249] & b[208])^(a[248] & b[209])^(a[247] & b[210])^(a[246] & b[211])^(a[245] & b[212])^(a[244] & b[213])^(a[243] & b[214])^(a[242] & b[215])^(a[241] & b[216])^(a[240] & b[217])^(a[239] & b[218])^(a[238] & b[219])^(a[237] & b[220])^(a[236] & b[221])^(a[235] & b[222])^(a[234] & b[223])^(a[233] & b[224])^(a[232] & b[225])^(a[231] & b[226])^(a[230] & b[227])^(a[229] & b[228])^(a[228] & b[229])^(a[227] & b[230])^(a[226] & b[231])^(a[225] & b[232])^(a[224] & b[233])^(a[223] & b[234])^(a[222] & b[235])^(a[221] & b[236])^(a[220] & b[237])^(a[219] & b[238])^(a[218] & b[239])^(a[217] & b[240])^(a[216] & b[241])^(a[215] & b[242])^(a[214] & b[243])^(a[213] & b[244])^(a[212] & b[245])^(a[211] & b[246])^(a[210] & b[247])^(a[209] & b[248])^(a[208] & b[249])^(a[207] & b[250])^(a[206] & b[251])^(a[205] & b[252])^(a[204] & b[253])^(a[203] & b[254])^(a[202] & b[255])^(a[201] & b[256])^(a[200] & b[257])^(a[199] & b[258])^(a[198] & b[259])^(a[197] & b[260])^(a[196] & b[261])^(a[195] & b[262])^(a[194] & b[263])^(a[193] & b[264])^(a[192] & b[265])^(a[191] & b[266])^(a[190] & b[267])^(a[189] & b[268])^(a[188] & b[269])^(a[187] & b[270])^(a[186] & b[271])^(a[185] & b[272])^(a[184] & b[273])^(a[183] & b[274])^(a[182] & b[275])^(a[181] & b[276])^(a[180] & b[277])^(a[179] & b[278])^(a[178] & b[279])^(a[177] & b[280])^(a[176] & b[281])^(a[175] & b[282])^(a[174] & b[283])^(a[173] & b[284])^(a[172] & b[285])^(a[171] & b[286])^(a[170] & b[287])^(a[169] & b[288])^(a[168] & b[289])^(a[167] & b[290])^(a[166] & b[291])^(a[165] & b[292])^(a[164] & b[293])^(a[163] & b[294])^(a[162] & b[295])^(a[161] & b[296])^(a[160] & b[297])^(a[159] & b[298])^(a[158] & b[299])^(a[157] & b[300])^(a[156] & b[301])^(a[155] & b[302])^(a[154] & b[303])^(a[153] & b[304])^(a[152] & b[305])^(a[151] & b[306])^(a[150] & b[307])^(a[149] & b[308])^(a[148] & b[309])^(a[147] & b[310])^(a[146] & b[311])^(a[145] & b[312])^(a[144] & b[313])^(a[143] & b[314])^(a[142] & b[315])^(a[141] & b[316])^(a[140] & b[317])^(a[139] & b[318])^(a[138] & b[319])^(a[137] & b[320])^(a[136] & b[321])^(a[135] & b[322])^(a[134] & b[323])^(a[133] & b[324])^(a[132] & b[325])^(a[131] & b[326])^(a[130] & b[327])^(a[129] & b[328])^(a[128] & b[329])^(a[127] & b[330])^(a[126] & b[331])^(a[125] & b[332])^(a[124] & b[333])^(a[123] & b[334])^(a[122] & b[335])^(a[121] & b[336])^(a[120] & b[337])^(a[119] & b[338])^(a[118] & b[339])^(a[117] & b[340])^(a[116] & b[341])^(a[115] & b[342])^(a[114] & b[343])^(a[113] & b[344])^(a[112] & b[345])^(a[111] & b[346])^(a[110] & b[347])^(a[109] & b[348])^(a[108] & b[349])^(a[107] & b[350])^(a[106] & b[351])^(a[105] & b[352])^(a[104] & b[353])^(a[103] & b[354])^(a[102] & b[355])^(a[101] & b[356])^(a[100] & b[357])^(a[99] & b[358])^(a[98] & b[359])^(a[97] & b[360])^(a[96] & b[361])^(a[95] & b[362])^(a[94] & b[363])^(a[93] & b[364])^(a[92] & b[365])^(a[91] & b[366])^(a[90] & b[367])^(a[89] & b[368])^(a[88] & b[369])^(a[87] & b[370])^(a[86] & b[371])^(a[85] & b[372])^(a[84] & b[373])^(a[83] & b[374])^(a[82] & b[375])^(a[81] & b[376])^(a[80] & b[377])^(a[79] & b[378])^(a[78] & b[379])^(a[77] & b[380])^(a[76] & b[381])^(a[75] & b[382])^(a[74] & b[383])^(a[73] & b[384])^(a[72] & b[385])^(a[71] & b[386])^(a[70] & b[387])^(a[69] & b[388])^(a[68] & b[389])^(a[67] & b[390])^(a[66] & b[391])^(a[65] & b[392])^(a[64] & b[393])^(a[63] & b[394])^(a[62] & b[395])^(a[61] & b[396])^(a[60] & b[397])^(a[59] & b[398])^(a[58] & b[399])^(a[57] & b[400])^(a[56] & b[401])^(a[55] & b[402])^(a[54] & b[403])^(a[53] & b[404])^(a[52] & b[405])^(a[51] & b[406])^(a[50] & b[407])^(a[49] & b[408]);
assign y[458] = (a[408] & b[50])^(a[407] & b[51])^(a[406] & b[52])^(a[405] & b[53])^(a[404] & b[54])^(a[403] & b[55])^(a[402] & b[56])^(a[401] & b[57])^(a[400] & b[58])^(a[399] & b[59])^(a[398] & b[60])^(a[397] & b[61])^(a[396] & b[62])^(a[395] & b[63])^(a[394] & b[64])^(a[393] & b[65])^(a[392] & b[66])^(a[391] & b[67])^(a[390] & b[68])^(a[389] & b[69])^(a[388] & b[70])^(a[387] & b[71])^(a[386] & b[72])^(a[385] & b[73])^(a[384] & b[74])^(a[383] & b[75])^(a[382] & b[76])^(a[381] & b[77])^(a[380] & b[78])^(a[379] & b[79])^(a[378] & b[80])^(a[377] & b[81])^(a[376] & b[82])^(a[375] & b[83])^(a[374] & b[84])^(a[373] & b[85])^(a[372] & b[86])^(a[371] & b[87])^(a[370] & b[88])^(a[369] & b[89])^(a[368] & b[90])^(a[367] & b[91])^(a[366] & b[92])^(a[365] & b[93])^(a[364] & b[94])^(a[363] & b[95])^(a[362] & b[96])^(a[361] & b[97])^(a[360] & b[98])^(a[359] & b[99])^(a[358] & b[100])^(a[357] & b[101])^(a[356] & b[102])^(a[355] & b[103])^(a[354] & b[104])^(a[353] & b[105])^(a[352] & b[106])^(a[351] & b[107])^(a[350] & b[108])^(a[349] & b[109])^(a[348] & b[110])^(a[347] & b[111])^(a[346] & b[112])^(a[345] & b[113])^(a[344] & b[114])^(a[343] & b[115])^(a[342] & b[116])^(a[341] & b[117])^(a[340] & b[118])^(a[339] & b[119])^(a[338] & b[120])^(a[337] & b[121])^(a[336] & b[122])^(a[335] & b[123])^(a[334] & b[124])^(a[333] & b[125])^(a[332] & b[126])^(a[331] & b[127])^(a[330] & b[128])^(a[329] & b[129])^(a[328] & b[130])^(a[327] & b[131])^(a[326] & b[132])^(a[325] & b[133])^(a[324] & b[134])^(a[323] & b[135])^(a[322] & b[136])^(a[321] & b[137])^(a[320] & b[138])^(a[319] & b[139])^(a[318] & b[140])^(a[317] & b[141])^(a[316] & b[142])^(a[315] & b[143])^(a[314] & b[144])^(a[313] & b[145])^(a[312] & b[146])^(a[311] & b[147])^(a[310] & b[148])^(a[309] & b[149])^(a[308] & b[150])^(a[307] & b[151])^(a[306] & b[152])^(a[305] & b[153])^(a[304] & b[154])^(a[303] & b[155])^(a[302] & b[156])^(a[301] & b[157])^(a[300] & b[158])^(a[299] & b[159])^(a[298] & b[160])^(a[297] & b[161])^(a[296] & b[162])^(a[295] & b[163])^(a[294] & b[164])^(a[293] & b[165])^(a[292] & b[166])^(a[291] & b[167])^(a[290] & b[168])^(a[289] & b[169])^(a[288] & b[170])^(a[287] & b[171])^(a[286] & b[172])^(a[285] & b[173])^(a[284] & b[174])^(a[283] & b[175])^(a[282] & b[176])^(a[281] & b[177])^(a[280] & b[178])^(a[279] & b[179])^(a[278] & b[180])^(a[277] & b[181])^(a[276] & b[182])^(a[275] & b[183])^(a[274] & b[184])^(a[273] & b[185])^(a[272] & b[186])^(a[271] & b[187])^(a[270] & b[188])^(a[269] & b[189])^(a[268] & b[190])^(a[267] & b[191])^(a[266] & b[192])^(a[265] & b[193])^(a[264] & b[194])^(a[263] & b[195])^(a[262] & b[196])^(a[261] & b[197])^(a[260] & b[198])^(a[259] & b[199])^(a[258] & b[200])^(a[257] & b[201])^(a[256] & b[202])^(a[255] & b[203])^(a[254] & b[204])^(a[253] & b[205])^(a[252] & b[206])^(a[251] & b[207])^(a[250] & b[208])^(a[249] & b[209])^(a[248] & b[210])^(a[247] & b[211])^(a[246] & b[212])^(a[245] & b[213])^(a[244] & b[214])^(a[243] & b[215])^(a[242] & b[216])^(a[241] & b[217])^(a[240] & b[218])^(a[239] & b[219])^(a[238] & b[220])^(a[237] & b[221])^(a[236] & b[222])^(a[235] & b[223])^(a[234] & b[224])^(a[233] & b[225])^(a[232] & b[226])^(a[231] & b[227])^(a[230] & b[228])^(a[229] & b[229])^(a[228] & b[230])^(a[227] & b[231])^(a[226] & b[232])^(a[225] & b[233])^(a[224] & b[234])^(a[223] & b[235])^(a[222] & b[236])^(a[221] & b[237])^(a[220] & b[238])^(a[219] & b[239])^(a[218] & b[240])^(a[217] & b[241])^(a[216] & b[242])^(a[215] & b[243])^(a[214] & b[244])^(a[213] & b[245])^(a[212] & b[246])^(a[211] & b[247])^(a[210] & b[248])^(a[209] & b[249])^(a[208] & b[250])^(a[207] & b[251])^(a[206] & b[252])^(a[205] & b[253])^(a[204] & b[254])^(a[203] & b[255])^(a[202] & b[256])^(a[201] & b[257])^(a[200] & b[258])^(a[199] & b[259])^(a[198] & b[260])^(a[197] & b[261])^(a[196] & b[262])^(a[195] & b[263])^(a[194] & b[264])^(a[193] & b[265])^(a[192] & b[266])^(a[191] & b[267])^(a[190] & b[268])^(a[189] & b[269])^(a[188] & b[270])^(a[187] & b[271])^(a[186] & b[272])^(a[185] & b[273])^(a[184] & b[274])^(a[183] & b[275])^(a[182] & b[276])^(a[181] & b[277])^(a[180] & b[278])^(a[179] & b[279])^(a[178] & b[280])^(a[177] & b[281])^(a[176] & b[282])^(a[175] & b[283])^(a[174] & b[284])^(a[173] & b[285])^(a[172] & b[286])^(a[171] & b[287])^(a[170] & b[288])^(a[169] & b[289])^(a[168] & b[290])^(a[167] & b[291])^(a[166] & b[292])^(a[165] & b[293])^(a[164] & b[294])^(a[163] & b[295])^(a[162] & b[296])^(a[161] & b[297])^(a[160] & b[298])^(a[159] & b[299])^(a[158] & b[300])^(a[157] & b[301])^(a[156] & b[302])^(a[155] & b[303])^(a[154] & b[304])^(a[153] & b[305])^(a[152] & b[306])^(a[151] & b[307])^(a[150] & b[308])^(a[149] & b[309])^(a[148] & b[310])^(a[147] & b[311])^(a[146] & b[312])^(a[145] & b[313])^(a[144] & b[314])^(a[143] & b[315])^(a[142] & b[316])^(a[141] & b[317])^(a[140] & b[318])^(a[139] & b[319])^(a[138] & b[320])^(a[137] & b[321])^(a[136] & b[322])^(a[135] & b[323])^(a[134] & b[324])^(a[133] & b[325])^(a[132] & b[326])^(a[131] & b[327])^(a[130] & b[328])^(a[129] & b[329])^(a[128] & b[330])^(a[127] & b[331])^(a[126] & b[332])^(a[125] & b[333])^(a[124] & b[334])^(a[123] & b[335])^(a[122] & b[336])^(a[121] & b[337])^(a[120] & b[338])^(a[119] & b[339])^(a[118] & b[340])^(a[117] & b[341])^(a[116] & b[342])^(a[115] & b[343])^(a[114] & b[344])^(a[113] & b[345])^(a[112] & b[346])^(a[111] & b[347])^(a[110] & b[348])^(a[109] & b[349])^(a[108] & b[350])^(a[107] & b[351])^(a[106] & b[352])^(a[105] & b[353])^(a[104] & b[354])^(a[103] & b[355])^(a[102] & b[356])^(a[101] & b[357])^(a[100] & b[358])^(a[99] & b[359])^(a[98] & b[360])^(a[97] & b[361])^(a[96] & b[362])^(a[95] & b[363])^(a[94] & b[364])^(a[93] & b[365])^(a[92] & b[366])^(a[91] & b[367])^(a[90] & b[368])^(a[89] & b[369])^(a[88] & b[370])^(a[87] & b[371])^(a[86] & b[372])^(a[85] & b[373])^(a[84] & b[374])^(a[83] & b[375])^(a[82] & b[376])^(a[81] & b[377])^(a[80] & b[378])^(a[79] & b[379])^(a[78] & b[380])^(a[77] & b[381])^(a[76] & b[382])^(a[75] & b[383])^(a[74] & b[384])^(a[73] & b[385])^(a[72] & b[386])^(a[71] & b[387])^(a[70] & b[388])^(a[69] & b[389])^(a[68] & b[390])^(a[67] & b[391])^(a[66] & b[392])^(a[65] & b[393])^(a[64] & b[394])^(a[63] & b[395])^(a[62] & b[396])^(a[61] & b[397])^(a[60] & b[398])^(a[59] & b[399])^(a[58] & b[400])^(a[57] & b[401])^(a[56] & b[402])^(a[55] & b[403])^(a[54] & b[404])^(a[53] & b[405])^(a[52] & b[406])^(a[51] & b[407])^(a[50] & b[408]);
assign y[459] = (a[408] & b[51])^(a[407] & b[52])^(a[406] & b[53])^(a[405] & b[54])^(a[404] & b[55])^(a[403] & b[56])^(a[402] & b[57])^(a[401] & b[58])^(a[400] & b[59])^(a[399] & b[60])^(a[398] & b[61])^(a[397] & b[62])^(a[396] & b[63])^(a[395] & b[64])^(a[394] & b[65])^(a[393] & b[66])^(a[392] & b[67])^(a[391] & b[68])^(a[390] & b[69])^(a[389] & b[70])^(a[388] & b[71])^(a[387] & b[72])^(a[386] & b[73])^(a[385] & b[74])^(a[384] & b[75])^(a[383] & b[76])^(a[382] & b[77])^(a[381] & b[78])^(a[380] & b[79])^(a[379] & b[80])^(a[378] & b[81])^(a[377] & b[82])^(a[376] & b[83])^(a[375] & b[84])^(a[374] & b[85])^(a[373] & b[86])^(a[372] & b[87])^(a[371] & b[88])^(a[370] & b[89])^(a[369] & b[90])^(a[368] & b[91])^(a[367] & b[92])^(a[366] & b[93])^(a[365] & b[94])^(a[364] & b[95])^(a[363] & b[96])^(a[362] & b[97])^(a[361] & b[98])^(a[360] & b[99])^(a[359] & b[100])^(a[358] & b[101])^(a[357] & b[102])^(a[356] & b[103])^(a[355] & b[104])^(a[354] & b[105])^(a[353] & b[106])^(a[352] & b[107])^(a[351] & b[108])^(a[350] & b[109])^(a[349] & b[110])^(a[348] & b[111])^(a[347] & b[112])^(a[346] & b[113])^(a[345] & b[114])^(a[344] & b[115])^(a[343] & b[116])^(a[342] & b[117])^(a[341] & b[118])^(a[340] & b[119])^(a[339] & b[120])^(a[338] & b[121])^(a[337] & b[122])^(a[336] & b[123])^(a[335] & b[124])^(a[334] & b[125])^(a[333] & b[126])^(a[332] & b[127])^(a[331] & b[128])^(a[330] & b[129])^(a[329] & b[130])^(a[328] & b[131])^(a[327] & b[132])^(a[326] & b[133])^(a[325] & b[134])^(a[324] & b[135])^(a[323] & b[136])^(a[322] & b[137])^(a[321] & b[138])^(a[320] & b[139])^(a[319] & b[140])^(a[318] & b[141])^(a[317] & b[142])^(a[316] & b[143])^(a[315] & b[144])^(a[314] & b[145])^(a[313] & b[146])^(a[312] & b[147])^(a[311] & b[148])^(a[310] & b[149])^(a[309] & b[150])^(a[308] & b[151])^(a[307] & b[152])^(a[306] & b[153])^(a[305] & b[154])^(a[304] & b[155])^(a[303] & b[156])^(a[302] & b[157])^(a[301] & b[158])^(a[300] & b[159])^(a[299] & b[160])^(a[298] & b[161])^(a[297] & b[162])^(a[296] & b[163])^(a[295] & b[164])^(a[294] & b[165])^(a[293] & b[166])^(a[292] & b[167])^(a[291] & b[168])^(a[290] & b[169])^(a[289] & b[170])^(a[288] & b[171])^(a[287] & b[172])^(a[286] & b[173])^(a[285] & b[174])^(a[284] & b[175])^(a[283] & b[176])^(a[282] & b[177])^(a[281] & b[178])^(a[280] & b[179])^(a[279] & b[180])^(a[278] & b[181])^(a[277] & b[182])^(a[276] & b[183])^(a[275] & b[184])^(a[274] & b[185])^(a[273] & b[186])^(a[272] & b[187])^(a[271] & b[188])^(a[270] & b[189])^(a[269] & b[190])^(a[268] & b[191])^(a[267] & b[192])^(a[266] & b[193])^(a[265] & b[194])^(a[264] & b[195])^(a[263] & b[196])^(a[262] & b[197])^(a[261] & b[198])^(a[260] & b[199])^(a[259] & b[200])^(a[258] & b[201])^(a[257] & b[202])^(a[256] & b[203])^(a[255] & b[204])^(a[254] & b[205])^(a[253] & b[206])^(a[252] & b[207])^(a[251] & b[208])^(a[250] & b[209])^(a[249] & b[210])^(a[248] & b[211])^(a[247] & b[212])^(a[246] & b[213])^(a[245] & b[214])^(a[244] & b[215])^(a[243] & b[216])^(a[242] & b[217])^(a[241] & b[218])^(a[240] & b[219])^(a[239] & b[220])^(a[238] & b[221])^(a[237] & b[222])^(a[236] & b[223])^(a[235] & b[224])^(a[234] & b[225])^(a[233] & b[226])^(a[232] & b[227])^(a[231] & b[228])^(a[230] & b[229])^(a[229] & b[230])^(a[228] & b[231])^(a[227] & b[232])^(a[226] & b[233])^(a[225] & b[234])^(a[224] & b[235])^(a[223] & b[236])^(a[222] & b[237])^(a[221] & b[238])^(a[220] & b[239])^(a[219] & b[240])^(a[218] & b[241])^(a[217] & b[242])^(a[216] & b[243])^(a[215] & b[244])^(a[214] & b[245])^(a[213] & b[246])^(a[212] & b[247])^(a[211] & b[248])^(a[210] & b[249])^(a[209] & b[250])^(a[208] & b[251])^(a[207] & b[252])^(a[206] & b[253])^(a[205] & b[254])^(a[204] & b[255])^(a[203] & b[256])^(a[202] & b[257])^(a[201] & b[258])^(a[200] & b[259])^(a[199] & b[260])^(a[198] & b[261])^(a[197] & b[262])^(a[196] & b[263])^(a[195] & b[264])^(a[194] & b[265])^(a[193] & b[266])^(a[192] & b[267])^(a[191] & b[268])^(a[190] & b[269])^(a[189] & b[270])^(a[188] & b[271])^(a[187] & b[272])^(a[186] & b[273])^(a[185] & b[274])^(a[184] & b[275])^(a[183] & b[276])^(a[182] & b[277])^(a[181] & b[278])^(a[180] & b[279])^(a[179] & b[280])^(a[178] & b[281])^(a[177] & b[282])^(a[176] & b[283])^(a[175] & b[284])^(a[174] & b[285])^(a[173] & b[286])^(a[172] & b[287])^(a[171] & b[288])^(a[170] & b[289])^(a[169] & b[290])^(a[168] & b[291])^(a[167] & b[292])^(a[166] & b[293])^(a[165] & b[294])^(a[164] & b[295])^(a[163] & b[296])^(a[162] & b[297])^(a[161] & b[298])^(a[160] & b[299])^(a[159] & b[300])^(a[158] & b[301])^(a[157] & b[302])^(a[156] & b[303])^(a[155] & b[304])^(a[154] & b[305])^(a[153] & b[306])^(a[152] & b[307])^(a[151] & b[308])^(a[150] & b[309])^(a[149] & b[310])^(a[148] & b[311])^(a[147] & b[312])^(a[146] & b[313])^(a[145] & b[314])^(a[144] & b[315])^(a[143] & b[316])^(a[142] & b[317])^(a[141] & b[318])^(a[140] & b[319])^(a[139] & b[320])^(a[138] & b[321])^(a[137] & b[322])^(a[136] & b[323])^(a[135] & b[324])^(a[134] & b[325])^(a[133] & b[326])^(a[132] & b[327])^(a[131] & b[328])^(a[130] & b[329])^(a[129] & b[330])^(a[128] & b[331])^(a[127] & b[332])^(a[126] & b[333])^(a[125] & b[334])^(a[124] & b[335])^(a[123] & b[336])^(a[122] & b[337])^(a[121] & b[338])^(a[120] & b[339])^(a[119] & b[340])^(a[118] & b[341])^(a[117] & b[342])^(a[116] & b[343])^(a[115] & b[344])^(a[114] & b[345])^(a[113] & b[346])^(a[112] & b[347])^(a[111] & b[348])^(a[110] & b[349])^(a[109] & b[350])^(a[108] & b[351])^(a[107] & b[352])^(a[106] & b[353])^(a[105] & b[354])^(a[104] & b[355])^(a[103] & b[356])^(a[102] & b[357])^(a[101] & b[358])^(a[100] & b[359])^(a[99] & b[360])^(a[98] & b[361])^(a[97] & b[362])^(a[96] & b[363])^(a[95] & b[364])^(a[94] & b[365])^(a[93] & b[366])^(a[92] & b[367])^(a[91] & b[368])^(a[90] & b[369])^(a[89] & b[370])^(a[88] & b[371])^(a[87] & b[372])^(a[86] & b[373])^(a[85] & b[374])^(a[84] & b[375])^(a[83] & b[376])^(a[82] & b[377])^(a[81] & b[378])^(a[80] & b[379])^(a[79] & b[380])^(a[78] & b[381])^(a[77] & b[382])^(a[76] & b[383])^(a[75] & b[384])^(a[74] & b[385])^(a[73] & b[386])^(a[72] & b[387])^(a[71] & b[388])^(a[70] & b[389])^(a[69] & b[390])^(a[68] & b[391])^(a[67] & b[392])^(a[66] & b[393])^(a[65] & b[394])^(a[64] & b[395])^(a[63] & b[396])^(a[62] & b[397])^(a[61] & b[398])^(a[60] & b[399])^(a[59] & b[400])^(a[58] & b[401])^(a[57] & b[402])^(a[56] & b[403])^(a[55] & b[404])^(a[54] & b[405])^(a[53] & b[406])^(a[52] & b[407])^(a[51] & b[408]);
assign y[460] = (a[408] & b[52])^(a[407] & b[53])^(a[406] & b[54])^(a[405] & b[55])^(a[404] & b[56])^(a[403] & b[57])^(a[402] & b[58])^(a[401] & b[59])^(a[400] & b[60])^(a[399] & b[61])^(a[398] & b[62])^(a[397] & b[63])^(a[396] & b[64])^(a[395] & b[65])^(a[394] & b[66])^(a[393] & b[67])^(a[392] & b[68])^(a[391] & b[69])^(a[390] & b[70])^(a[389] & b[71])^(a[388] & b[72])^(a[387] & b[73])^(a[386] & b[74])^(a[385] & b[75])^(a[384] & b[76])^(a[383] & b[77])^(a[382] & b[78])^(a[381] & b[79])^(a[380] & b[80])^(a[379] & b[81])^(a[378] & b[82])^(a[377] & b[83])^(a[376] & b[84])^(a[375] & b[85])^(a[374] & b[86])^(a[373] & b[87])^(a[372] & b[88])^(a[371] & b[89])^(a[370] & b[90])^(a[369] & b[91])^(a[368] & b[92])^(a[367] & b[93])^(a[366] & b[94])^(a[365] & b[95])^(a[364] & b[96])^(a[363] & b[97])^(a[362] & b[98])^(a[361] & b[99])^(a[360] & b[100])^(a[359] & b[101])^(a[358] & b[102])^(a[357] & b[103])^(a[356] & b[104])^(a[355] & b[105])^(a[354] & b[106])^(a[353] & b[107])^(a[352] & b[108])^(a[351] & b[109])^(a[350] & b[110])^(a[349] & b[111])^(a[348] & b[112])^(a[347] & b[113])^(a[346] & b[114])^(a[345] & b[115])^(a[344] & b[116])^(a[343] & b[117])^(a[342] & b[118])^(a[341] & b[119])^(a[340] & b[120])^(a[339] & b[121])^(a[338] & b[122])^(a[337] & b[123])^(a[336] & b[124])^(a[335] & b[125])^(a[334] & b[126])^(a[333] & b[127])^(a[332] & b[128])^(a[331] & b[129])^(a[330] & b[130])^(a[329] & b[131])^(a[328] & b[132])^(a[327] & b[133])^(a[326] & b[134])^(a[325] & b[135])^(a[324] & b[136])^(a[323] & b[137])^(a[322] & b[138])^(a[321] & b[139])^(a[320] & b[140])^(a[319] & b[141])^(a[318] & b[142])^(a[317] & b[143])^(a[316] & b[144])^(a[315] & b[145])^(a[314] & b[146])^(a[313] & b[147])^(a[312] & b[148])^(a[311] & b[149])^(a[310] & b[150])^(a[309] & b[151])^(a[308] & b[152])^(a[307] & b[153])^(a[306] & b[154])^(a[305] & b[155])^(a[304] & b[156])^(a[303] & b[157])^(a[302] & b[158])^(a[301] & b[159])^(a[300] & b[160])^(a[299] & b[161])^(a[298] & b[162])^(a[297] & b[163])^(a[296] & b[164])^(a[295] & b[165])^(a[294] & b[166])^(a[293] & b[167])^(a[292] & b[168])^(a[291] & b[169])^(a[290] & b[170])^(a[289] & b[171])^(a[288] & b[172])^(a[287] & b[173])^(a[286] & b[174])^(a[285] & b[175])^(a[284] & b[176])^(a[283] & b[177])^(a[282] & b[178])^(a[281] & b[179])^(a[280] & b[180])^(a[279] & b[181])^(a[278] & b[182])^(a[277] & b[183])^(a[276] & b[184])^(a[275] & b[185])^(a[274] & b[186])^(a[273] & b[187])^(a[272] & b[188])^(a[271] & b[189])^(a[270] & b[190])^(a[269] & b[191])^(a[268] & b[192])^(a[267] & b[193])^(a[266] & b[194])^(a[265] & b[195])^(a[264] & b[196])^(a[263] & b[197])^(a[262] & b[198])^(a[261] & b[199])^(a[260] & b[200])^(a[259] & b[201])^(a[258] & b[202])^(a[257] & b[203])^(a[256] & b[204])^(a[255] & b[205])^(a[254] & b[206])^(a[253] & b[207])^(a[252] & b[208])^(a[251] & b[209])^(a[250] & b[210])^(a[249] & b[211])^(a[248] & b[212])^(a[247] & b[213])^(a[246] & b[214])^(a[245] & b[215])^(a[244] & b[216])^(a[243] & b[217])^(a[242] & b[218])^(a[241] & b[219])^(a[240] & b[220])^(a[239] & b[221])^(a[238] & b[222])^(a[237] & b[223])^(a[236] & b[224])^(a[235] & b[225])^(a[234] & b[226])^(a[233] & b[227])^(a[232] & b[228])^(a[231] & b[229])^(a[230] & b[230])^(a[229] & b[231])^(a[228] & b[232])^(a[227] & b[233])^(a[226] & b[234])^(a[225] & b[235])^(a[224] & b[236])^(a[223] & b[237])^(a[222] & b[238])^(a[221] & b[239])^(a[220] & b[240])^(a[219] & b[241])^(a[218] & b[242])^(a[217] & b[243])^(a[216] & b[244])^(a[215] & b[245])^(a[214] & b[246])^(a[213] & b[247])^(a[212] & b[248])^(a[211] & b[249])^(a[210] & b[250])^(a[209] & b[251])^(a[208] & b[252])^(a[207] & b[253])^(a[206] & b[254])^(a[205] & b[255])^(a[204] & b[256])^(a[203] & b[257])^(a[202] & b[258])^(a[201] & b[259])^(a[200] & b[260])^(a[199] & b[261])^(a[198] & b[262])^(a[197] & b[263])^(a[196] & b[264])^(a[195] & b[265])^(a[194] & b[266])^(a[193] & b[267])^(a[192] & b[268])^(a[191] & b[269])^(a[190] & b[270])^(a[189] & b[271])^(a[188] & b[272])^(a[187] & b[273])^(a[186] & b[274])^(a[185] & b[275])^(a[184] & b[276])^(a[183] & b[277])^(a[182] & b[278])^(a[181] & b[279])^(a[180] & b[280])^(a[179] & b[281])^(a[178] & b[282])^(a[177] & b[283])^(a[176] & b[284])^(a[175] & b[285])^(a[174] & b[286])^(a[173] & b[287])^(a[172] & b[288])^(a[171] & b[289])^(a[170] & b[290])^(a[169] & b[291])^(a[168] & b[292])^(a[167] & b[293])^(a[166] & b[294])^(a[165] & b[295])^(a[164] & b[296])^(a[163] & b[297])^(a[162] & b[298])^(a[161] & b[299])^(a[160] & b[300])^(a[159] & b[301])^(a[158] & b[302])^(a[157] & b[303])^(a[156] & b[304])^(a[155] & b[305])^(a[154] & b[306])^(a[153] & b[307])^(a[152] & b[308])^(a[151] & b[309])^(a[150] & b[310])^(a[149] & b[311])^(a[148] & b[312])^(a[147] & b[313])^(a[146] & b[314])^(a[145] & b[315])^(a[144] & b[316])^(a[143] & b[317])^(a[142] & b[318])^(a[141] & b[319])^(a[140] & b[320])^(a[139] & b[321])^(a[138] & b[322])^(a[137] & b[323])^(a[136] & b[324])^(a[135] & b[325])^(a[134] & b[326])^(a[133] & b[327])^(a[132] & b[328])^(a[131] & b[329])^(a[130] & b[330])^(a[129] & b[331])^(a[128] & b[332])^(a[127] & b[333])^(a[126] & b[334])^(a[125] & b[335])^(a[124] & b[336])^(a[123] & b[337])^(a[122] & b[338])^(a[121] & b[339])^(a[120] & b[340])^(a[119] & b[341])^(a[118] & b[342])^(a[117] & b[343])^(a[116] & b[344])^(a[115] & b[345])^(a[114] & b[346])^(a[113] & b[347])^(a[112] & b[348])^(a[111] & b[349])^(a[110] & b[350])^(a[109] & b[351])^(a[108] & b[352])^(a[107] & b[353])^(a[106] & b[354])^(a[105] & b[355])^(a[104] & b[356])^(a[103] & b[357])^(a[102] & b[358])^(a[101] & b[359])^(a[100] & b[360])^(a[99] & b[361])^(a[98] & b[362])^(a[97] & b[363])^(a[96] & b[364])^(a[95] & b[365])^(a[94] & b[366])^(a[93] & b[367])^(a[92] & b[368])^(a[91] & b[369])^(a[90] & b[370])^(a[89] & b[371])^(a[88] & b[372])^(a[87] & b[373])^(a[86] & b[374])^(a[85] & b[375])^(a[84] & b[376])^(a[83] & b[377])^(a[82] & b[378])^(a[81] & b[379])^(a[80] & b[380])^(a[79] & b[381])^(a[78] & b[382])^(a[77] & b[383])^(a[76] & b[384])^(a[75] & b[385])^(a[74] & b[386])^(a[73] & b[387])^(a[72] & b[388])^(a[71] & b[389])^(a[70] & b[390])^(a[69] & b[391])^(a[68] & b[392])^(a[67] & b[393])^(a[66] & b[394])^(a[65] & b[395])^(a[64] & b[396])^(a[63] & b[397])^(a[62] & b[398])^(a[61] & b[399])^(a[60] & b[400])^(a[59] & b[401])^(a[58] & b[402])^(a[57] & b[403])^(a[56] & b[404])^(a[55] & b[405])^(a[54] & b[406])^(a[53] & b[407])^(a[52] & b[408]);
assign y[461] = (a[408] & b[53])^(a[407] & b[54])^(a[406] & b[55])^(a[405] & b[56])^(a[404] & b[57])^(a[403] & b[58])^(a[402] & b[59])^(a[401] & b[60])^(a[400] & b[61])^(a[399] & b[62])^(a[398] & b[63])^(a[397] & b[64])^(a[396] & b[65])^(a[395] & b[66])^(a[394] & b[67])^(a[393] & b[68])^(a[392] & b[69])^(a[391] & b[70])^(a[390] & b[71])^(a[389] & b[72])^(a[388] & b[73])^(a[387] & b[74])^(a[386] & b[75])^(a[385] & b[76])^(a[384] & b[77])^(a[383] & b[78])^(a[382] & b[79])^(a[381] & b[80])^(a[380] & b[81])^(a[379] & b[82])^(a[378] & b[83])^(a[377] & b[84])^(a[376] & b[85])^(a[375] & b[86])^(a[374] & b[87])^(a[373] & b[88])^(a[372] & b[89])^(a[371] & b[90])^(a[370] & b[91])^(a[369] & b[92])^(a[368] & b[93])^(a[367] & b[94])^(a[366] & b[95])^(a[365] & b[96])^(a[364] & b[97])^(a[363] & b[98])^(a[362] & b[99])^(a[361] & b[100])^(a[360] & b[101])^(a[359] & b[102])^(a[358] & b[103])^(a[357] & b[104])^(a[356] & b[105])^(a[355] & b[106])^(a[354] & b[107])^(a[353] & b[108])^(a[352] & b[109])^(a[351] & b[110])^(a[350] & b[111])^(a[349] & b[112])^(a[348] & b[113])^(a[347] & b[114])^(a[346] & b[115])^(a[345] & b[116])^(a[344] & b[117])^(a[343] & b[118])^(a[342] & b[119])^(a[341] & b[120])^(a[340] & b[121])^(a[339] & b[122])^(a[338] & b[123])^(a[337] & b[124])^(a[336] & b[125])^(a[335] & b[126])^(a[334] & b[127])^(a[333] & b[128])^(a[332] & b[129])^(a[331] & b[130])^(a[330] & b[131])^(a[329] & b[132])^(a[328] & b[133])^(a[327] & b[134])^(a[326] & b[135])^(a[325] & b[136])^(a[324] & b[137])^(a[323] & b[138])^(a[322] & b[139])^(a[321] & b[140])^(a[320] & b[141])^(a[319] & b[142])^(a[318] & b[143])^(a[317] & b[144])^(a[316] & b[145])^(a[315] & b[146])^(a[314] & b[147])^(a[313] & b[148])^(a[312] & b[149])^(a[311] & b[150])^(a[310] & b[151])^(a[309] & b[152])^(a[308] & b[153])^(a[307] & b[154])^(a[306] & b[155])^(a[305] & b[156])^(a[304] & b[157])^(a[303] & b[158])^(a[302] & b[159])^(a[301] & b[160])^(a[300] & b[161])^(a[299] & b[162])^(a[298] & b[163])^(a[297] & b[164])^(a[296] & b[165])^(a[295] & b[166])^(a[294] & b[167])^(a[293] & b[168])^(a[292] & b[169])^(a[291] & b[170])^(a[290] & b[171])^(a[289] & b[172])^(a[288] & b[173])^(a[287] & b[174])^(a[286] & b[175])^(a[285] & b[176])^(a[284] & b[177])^(a[283] & b[178])^(a[282] & b[179])^(a[281] & b[180])^(a[280] & b[181])^(a[279] & b[182])^(a[278] & b[183])^(a[277] & b[184])^(a[276] & b[185])^(a[275] & b[186])^(a[274] & b[187])^(a[273] & b[188])^(a[272] & b[189])^(a[271] & b[190])^(a[270] & b[191])^(a[269] & b[192])^(a[268] & b[193])^(a[267] & b[194])^(a[266] & b[195])^(a[265] & b[196])^(a[264] & b[197])^(a[263] & b[198])^(a[262] & b[199])^(a[261] & b[200])^(a[260] & b[201])^(a[259] & b[202])^(a[258] & b[203])^(a[257] & b[204])^(a[256] & b[205])^(a[255] & b[206])^(a[254] & b[207])^(a[253] & b[208])^(a[252] & b[209])^(a[251] & b[210])^(a[250] & b[211])^(a[249] & b[212])^(a[248] & b[213])^(a[247] & b[214])^(a[246] & b[215])^(a[245] & b[216])^(a[244] & b[217])^(a[243] & b[218])^(a[242] & b[219])^(a[241] & b[220])^(a[240] & b[221])^(a[239] & b[222])^(a[238] & b[223])^(a[237] & b[224])^(a[236] & b[225])^(a[235] & b[226])^(a[234] & b[227])^(a[233] & b[228])^(a[232] & b[229])^(a[231] & b[230])^(a[230] & b[231])^(a[229] & b[232])^(a[228] & b[233])^(a[227] & b[234])^(a[226] & b[235])^(a[225] & b[236])^(a[224] & b[237])^(a[223] & b[238])^(a[222] & b[239])^(a[221] & b[240])^(a[220] & b[241])^(a[219] & b[242])^(a[218] & b[243])^(a[217] & b[244])^(a[216] & b[245])^(a[215] & b[246])^(a[214] & b[247])^(a[213] & b[248])^(a[212] & b[249])^(a[211] & b[250])^(a[210] & b[251])^(a[209] & b[252])^(a[208] & b[253])^(a[207] & b[254])^(a[206] & b[255])^(a[205] & b[256])^(a[204] & b[257])^(a[203] & b[258])^(a[202] & b[259])^(a[201] & b[260])^(a[200] & b[261])^(a[199] & b[262])^(a[198] & b[263])^(a[197] & b[264])^(a[196] & b[265])^(a[195] & b[266])^(a[194] & b[267])^(a[193] & b[268])^(a[192] & b[269])^(a[191] & b[270])^(a[190] & b[271])^(a[189] & b[272])^(a[188] & b[273])^(a[187] & b[274])^(a[186] & b[275])^(a[185] & b[276])^(a[184] & b[277])^(a[183] & b[278])^(a[182] & b[279])^(a[181] & b[280])^(a[180] & b[281])^(a[179] & b[282])^(a[178] & b[283])^(a[177] & b[284])^(a[176] & b[285])^(a[175] & b[286])^(a[174] & b[287])^(a[173] & b[288])^(a[172] & b[289])^(a[171] & b[290])^(a[170] & b[291])^(a[169] & b[292])^(a[168] & b[293])^(a[167] & b[294])^(a[166] & b[295])^(a[165] & b[296])^(a[164] & b[297])^(a[163] & b[298])^(a[162] & b[299])^(a[161] & b[300])^(a[160] & b[301])^(a[159] & b[302])^(a[158] & b[303])^(a[157] & b[304])^(a[156] & b[305])^(a[155] & b[306])^(a[154] & b[307])^(a[153] & b[308])^(a[152] & b[309])^(a[151] & b[310])^(a[150] & b[311])^(a[149] & b[312])^(a[148] & b[313])^(a[147] & b[314])^(a[146] & b[315])^(a[145] & b[316])^(a[144] & b[317])^(a[143] & b[318])^(a[142] & b[319])^(a[141] & b[320])^(a[140] & b[321])^(a[139] & b[322])^(a[138] & b[323])^(a[137] & b[324])^(a[136] & b[325])^(a[135] & b[326])^(a[134] & b[327])^(a[133] & b[328])^(a[132] & b[329])^(a[131] & b[330])^(a[130] & b[331])^(a[129] & b[332])^(a[128] & b[333])^(a[127] & b[334])^(a[126] & b[335])^(a[125] & b[336])^(a[124] & b[337])^(a[123] & b[338])^(a[122] & b[339])^(a[121] & b[340])^(a[120] & b[341])^(a[119] & b[342])^(a[118] & b[343])^(a[117] & b[344])^(a[116] & b[345])^(a[115] & b[346])^(a[114] & b[347])^(a[113] & b[348])^(a[112] & b[349])^(a[111] & b[350])^(a[110] & b[351])^(a[109] & b[352])^(a[108] & b[353])^(a[107] & b[354])^(a[106] & b[355])^(a[105] & b[356])^(a[104] & b[357])^(a[103] & b[358])^(a[102] & b[359])^(a[101] & b[360])^(a[100] & b[361])^(a[99] & b[362])^(a[98] & b[363])^(a[97] & b[364])^(a[96] & b[365])^(a[95] & b[366])^(a[94] & b[367])^(a[93] & b[368])^(a[92] & b[369])^(a[91] & b[370])^(a[90] & b[371])^(a[89] & b[372])^(a[88] & b[373])^(a[87] & b[374])^(a[86] & b[375])^(a[85] & b[376])^(a[84] & b[377])^(a[83] & b[378])^(a[82] & b[379])^(a[81] & b[380])^(a[80] & b[381])^(a[79] & b[382])^(a[78] & b[383])^(a[77] & b[384])^(a[76] & b[385])^(a[75] & b[386])^(a[74] & b[387])^(a[73] & b[388])^(a[72] & b[389])^(a[71] & b[390])^(a[70] & b[391])^(a[69] & b[392])^(a[68] & b[393])^(a[67] & b[394])^(a[66] & b[395])^(a[65] & b[396])^(a[64] & b[397])^(a[63] & b[398])^(a[62] & b[399])^(a[61] & b[400])^(a[60] & b[401])^(a[59] & b[402])^(a[58] & b[403])^(a[57] & b[404])^(a[56] & b[405])^(a[55] & b[406])^(a[54] & b[407])^(a[53] & b[408]);
assign y[462] = (a[408] & b[54])^(a[407] & b[55])^(a[406] & b[56])^(a[405] & b[57])^(a[404] & b[58])^(a[403] & b[59])^(a[402] & b[60])^(a[401] & b[61])^(a[400] & b[62])^(a[399] & b[63])^(a[398] & b[64])^(a[397] & b[65])^(a[396] & b[66])^(a[395] & b[67])^(a[394] & b[68])^(a[393] & b[69])^(a[392] & b[70])^(a[391] & b[71])^(a[390] & b[72])^(a[389] & b[73])^(a[388] & b[74])^(a[387] & b[75])^(a[386] & b[76])^(a[385] & b[77])^(a[384] & b[78])^(a[383] & b[79])^(a[382] & b[80])^(a[381] & b[81])^(a[380] & b[82])^(a[379] & b[83])^(a[378] & b[84])^(a[377] & b[85])^(a[376] & b[86])^(a[375] & b[87])^(a[374] & b[88])^(a[373] & b[89])^(a[372] & b[90])^(a[371] & b[91])^(a[370] & b[92])^(a[369] & b[93])^(a[368] & b[94])^(a[367] & b[95])^(a[366] & b[96])^(a[365] & b[97])^(a[364] & b[98])^(a[363] & b[99])^(a[362] & b[100])^(a[361] & b[101])^(a[360] & b[102])^(a[359] & b[103])^(a[358] & b[104])^(a[357] & b[105])^(a[356] & b[106])^(a[355] & b[107])^(a[354] & b[108])^(a[353] & b[109])^(a[352] & b[110])^(a[351] & b[111])^(a[350] & b[112])^(a[349] & b[113])^(a[348] & b[114])^(a[347] & b[115])^(a[346] & b[116])^(a[345] & b[117])^(a[344] & b[118])^(a[343] & b[119])^(a[342] & b[120])^(a[341] & b[121])^(a[340] & b[122])^(a[339] & b[123])^(a[338] & b[124])^(a[337] & b[125])^(a[336] & b[126])^(a[335] & b[127])^(a[334] & b[128])^(a[333] & b[129])^(a[332] & b[130])^(a[331] & b[131])^(a[330] & b[132])^(a[329] & b[133])^(a[328] & b[134])^(a[327] & b[135])^(a[326] & b[136])^(a[325] & b[137])^(a[324] & b[138])^(a[323] & b[139])^(a[322] & b[140])^(a[321] & b[141])^(a[320] & b[142])^(a[319] & b[143])^(a[318] & b[144])^(a[317] & b[145])^(a[316] & b[146])^(a[315] & b[147])^(a[314] & b[148])^(a[313] & b[149])^(a[312] & b[150])^(a[311] & b[151])^(a[310] & b[152])^(a[309] & b[153])^(a[308] & b[154])^(a[307] & b[155])^(a[306] & b[156])^(a[305] & b[157])^(a[304] & b[158])^(a[303] & b[159])^(a[302] & b[160])^(a[301] & b[161])^(a[300] & b[162])^(a[299] & b[163])^(a[298] & b[164])^(a[297] & b[165])^(a[296] & b[166])^(a[295] & b[167])^(a[294] & b[168])^(a[293] & b[169])^(a[292] & b[170])^(a[291] & b[171])^(a[290] & b[172])^(a[289] & b[173])^(a[288] & b[174])^(a[287] & b[175])^(a[286] & b[176])^(a[285] & b[177])^(a[284] & b[178])^(a[283] & b[179])^(a[282] & b[180])^(a[281] & b[181])^(a[280] & b[182])^(a[279] & b[183])^(a[278] & b[184])^(a[277] & b[185])^(a[276] & b[186])^(a[275] & b[187])^(a[274] & b[188])^(a[273] & b[189])^(a[272] & b[190])^(a[271] & b[191])^(a[270] & b[192])^(a[269] & b[193])^(a[268] & b[194])^(a[267] & b[195])^(a[266] & b[196])^(a[265] & b[197])^(a[264] & b[198])^(a[263] & b[199])^(a[262] & b[200])^(a[261] & b[201])^(a[260] & b[202])^(a[259] & b[203])^(a[258] & b[204])^(a[257] & b[205])^(a[256] & b[206])^(a[255] & b[207])^(a[254] & b[208])^(a[253] & b[209])^(a[252] & b[210])^(a[251] & b[211])^(a[250] & b[212])^(a[249] & b[213])^(a[248] & b[214])^(a[247] & b[215])^(a[246] & b[216])^(a[245] & b[217])^(a[244] & b[218])^(a[243] & b[219])^(a[242] & b[220])^(a[241] & b[221])^(a[240] & b[222])^(a[239] & b[223])^(a[238] & b[224])^(a[237] & b[225])^(a[236] & b[226])^(a[235] & b[227])^(a[234] & b[228])^(a[233] & b[229])^(a[232] & b[230])^(a[231] & b[231])^(a[230] & b[232])^(a[229] & b[233])^(a[228] & b[234])^(a[227] & b[235])^(a[226] & b[236])^(a[225] & b[237])^(a[224] & b[238])^(a[223] & b[239])^(a[222] & b[240])^(a[221] & b[241])^(a[220] & b[242])^(a[219] & b[243])^(a[218] & b[244])^(a[217] & b[245])^(a[216] & b[246])^(a[215] & b[247])^(a[214] & b[248])^(a[213] & b[249])^(a[212] & b[250])^(a[211] & b[251])^(a[210] & b[252])^(a[209] & b[253])^(a[208] & b[254])^(a[207] & b[255])^(a[206] & b[256])^(a[205] & b[257])^(a[204] & b[258])^(a[203] & b[259])^(a[202] & b[260])^(a[201] & b[261])^(a[200] & b[262])^(a[199] & b[263])^(a[198] & b[264])^(a[197] & b[265])^(a[196] & b[266])^(a[195] & b[267])^(a[194] & b[268])^(a[193] & b[269])^(a[192] & b[270])^(a[191] & b[271])^(a[190] & b[272])^(a[189] & b[273])^(a[188] & b[274])^(a[187] & b[275])^(a[186] & b[276])^(a[185] & b[277])^(a[184] & b[278])^(a[183] & b[279])^(a[182] & b[280])^(a[181] & b[281])^(a[180] & b[282])^(a[179] & b[283])^(a[178] & b[284])^(a[177] & b[285])^(a[176] & b[286])^(a[175] & b[287])^(a[174] & b[288])^(a[173] & b[289])^(a[172] & b[290])^(a[171] & b[291])^(a[170] & b[292])^(a[169] & b[293])^(a[168] & b[294])^(a[167] & b[295])^(a[166] & b[296])^(a[165] & b[297])^(a[164] & b[298])^(a[163] & b[299])^(a[162] & b[300])^(a[161] & b[301])^(a[160] & b[302])^(a[159] & b[303])^(a[158] & b[304])^(a[157] & b[305])^(a[156] & b[306])^(a[155] & b[307])^(a[154] & b[308])^(a[153] & b[309])^(a[152] & b[310])^(a[151] & b[311])^(a[150] & b[312])^(a[149] & b[313])^(a[148] & b[314])^(a[147] & b[315])^(a[146] & b[316])^(a[145] & b[317])^(a[144] & b[318])^(a[143] & b[319])^(a[142] & b[320])^(a[141] & b[321])^(a[140] & b[322])^(a[139] & b[323])^(a[138] & b[324])^(a[137] & b[325])^(a[136] & b[326])^(a[135] & b[327])^(a[134] & b[328])^(a[133] & b[329])^(a[132] & b[330])^(a[131] & b[331])^(a[130] & b[332])^(a[129] & b[333])^(a[128] & b[334])^(a[127] & b[335])^(a[126] & b[336])^(a[125] & b[337])^(a[124] & b[338])^(a[123] & b[339])^(a[122] & b[340])^(a[121] & b[341])^(a[120] & b[342])^(a[119] & b[343])^(a[118] & b[344])^(a[117] & b[345])^(a[116] & b[346])^(a[115] & b[347])^(a[114] & b[348])^(a[113] & b[349])^(a[112] & b[350])^(a[111] & b[351])^(a[110] & b[352])^(a[109] & b[353])^(a[108] & b[354])^(a[107] & b[355])^(a[106] & b[356])^(a[105] & b[357])^(a[104] & b[358])^(a[103] & b[359])^(a[102] & b[360])^(a[101] & b[361])^(a[100] & b[362])^(a[99] & b[363])^(a[98] & b[364])^(a[97] & b[365])^(a[96] & b[366])^(a[95] & b[367])^(a[94] & b[368])^(a[93] & b[369])^(a[92] & b[370])^(a[91] & b[371])^(a[90] & b[372])^(a[89] & b[373])^(a[88] & b[374])^(a[87] & b[375])^(a[86] & b[376])^(a[85] & b[377])^(a[84] & b[378])^(a[83] & b[379])^(a[82] & b[380])^(a[81] & b[381])^(a[80] & b[382])^(a[79] & b[383])^(a[78] & b[384])^(a[77] & b[385])^(a[76] & b[386])^(a[75] & b[387])^(a[74] & b[388])^(a[73] & b[389])^(a[72] & b[390])^(a[71] & b[391])^(a[70] & b[392])^(a[69] & b[393])^(a[68] & b[394])^(a[67] & b[395])^(a[66] & b[396])^(a[65] & b[397])^(a[64] & b[398])^(a[63] & b[399])^(a[62] & b[400])^(a[61] & b[401])^(a[60] & b[402])^(a[59] & b[403])^(a[58] & b[404])^(a[57] & b[405])^(a[56] & b[406])^(a[55] & b[407])^(a[54] & b[408]);
assign y[463] = (a[408] & b[55])^(a[407] & b[56])^(a[406] & b[57])^(a[405] & b[58])^(a[404] & b[59])^(a[403] & b[60])^(a[402] & b[61])^(a[401] & b[62])^(a[400] & b[63])^(a[399] & b[64])^(a[398] & b[65])^(a[397] & b[66])^(a[396] & b[67])^(a[395] & b[68])^(a[394] & b[69])^(a[393] & b[70])^(a[392] & b[71])^(a[391] & b[72])^(a[390] & b[73])^(a[389] & b[74])^(a[388] & b[75])^(a[387] & b[76])^(a[386] & b[77])^(a[385] & b[78])^(a[384] & b[79])^(a[383] & b[80])^(a[382] & b[81])^(a[381] & b[82])^(a[380] & b[83])^(a[379] & b[84])^(a[378] & b[85])^(a[377] & b[86])^(a[376] & b[87])^(a[375] & b[88])^(a[374] & b[89])^(a[373] & b[90])^(a[372] & b[91])^(a[371] & b[92])^(a[370] & b[93])^(a[369] & b[94])^(a[368] & b[95])^(a[367] & b[96])^(a[366] & b[97])^(a[365] & b[98])^(a[364] & b[99])^(a[363] & b[100])^(a[362] & b[101])^(a[361] & b[102])^(a[360] & b[103])^(a[359] & b[104])^(a[358] & b[105])^(a[357] & b[106])^(a[356] & b[107])^(a[355] & b[108])^(a[354] & b[109])^(a[353] & b[110])^(a[352] & b[111])^(a[351] & b[112])^(a[350] & b[113])^(a[349] & b[114])^(a[348] & b[115])^(a[347] & b[116])^(a[346] & b[117])^(a[345] & b[118])^(a[344] & b[119])^(a[343] & b[120])^(a[342] & b[121])^(a[341] & b[122])^(a[340] & b[123])^(a[339] & b[124])^(a[338] & b[125])^(a[337] & b[126])^(a[336] & b[127])^(a[335] & b[128])^(a[334] & b[129])^(a[333] & b[130])^(a[332] & b[131])^(a[331] & b[132])^(a[330] & b[133])^(a[329] & b[134])^(a[328] & b[135])^(a[327] & b[136])^(a[326] & b[137])^(a[325] & b[138])^(a[324] & b[139])^(a[323] & b[140])^(a[322] & b[141])^(a[321] & b[142])^(a[320] & b[143])^(a[319] & b[144])^(a[318] & b[145])^(a[317] & b[146])^(a[316] & b[147])^(a[315] & b[148])^(a[314] & b[149])^(a[313] & b[150])^(a[312] & b[151])^(a[311] & b[152])^(a[310] & b[153])^(a[309] & b[154])^(a[308] & b[155])^(a[307] & b[156])^(a[306] & b[157])^(a[305] & b[158])^(a[304] & b[159])^(a[303] & b[160])^(a[302] & b[161])^(a[301] & b[162])^(a[300] & b[163])^(a[299] & b[164])^(a[298] & b[165])^(a[297] & b[166])^(a[296] & b[167])^(a[295] & b[168])^(a[294] & b[169])^(a[293] & b[170])^(a[292] & b[171])^(a[291] & b[172])^(a[290] & b[173])^(a[289] & b[174])^(a[288] & b[175])^(a[287] & b[176])^(a[286] & b[177])^(a[285] & b[178])^(a[284] & b[179])^(a[283] & b[180])^(a[282] & b[181])^(a[281] & b[182])^(a[280] & b[183])^(a[279] & b[184])^(a[278] & b[185])^(a[277] & b[186])^(a[276] & b[187])^(a[275] & b[188])^(a[274] & b[189])^(a[273] & b[190])^(a[272] & b[191])^(a[271] & b[192])^(a[270] & b[193])^(a[269] & b[194])^(a[268] & b[195])^(a[267] & b[196])^(a[266] & b[197])^(a[265] & b[198])^(a[264] & b[199])^(a[263] & b[200])^(a[262] & b[201])^(a[261] & b[202])^(a[260] & b[203])^(a[259] & b[204])^(a[258] & b[205])^(a[257] & b[206])^(a[256] & b[207])^(a[255] & b[208])^(a[254] & b[209])^(a[253] & b[210])^(a[252] & b[211])^(a[251] & b[212])^(a[250] & b[213])^(a[249] & b[214])^(a[248] & b[215])^(a[247] & b[216])^(a[246] & b[217])^(a[245] & b[218])^(a[244] & b[219])^(a[243] & b[220])^(a[242] & b[221])^(a[241] & b[222])^(a[240] & b[223])^(a[239] & b[224])^(a[238] & b[225])^(a[237] & b[226])^(a[236] & b[227])^(a[235] & b[228])^(a[234] & b[229])^(a[233] & b[230])^(a[232] & b[231])^(a[231] & b[232])^(a[230] & b[233])^(a[229] & b[234])^(a[228] & b[235])^(a[227] & b[236])^(a[226] & b[237])^(a[225] & b[238])^(a[224] & b[239])^(a[223] & b[240])^(a[222] & b[241])^(a[221] & b[242])^(a[220] & b[243])^(a[219] & b[244])^(a[218] & b[245])^(a[217] & b[246])^(a[216] & b[247])^(a[215] & b[248])^(a[214] & b[249])^(a[213] & b[250])^(a[212] & b[251])^(a[211] & b[252])^(a[210] & b[253])^(a[209] & b[254])^(a[208] & b[255])^(a[207] & b[256])^(a[206] & b[257])^(a[205] & b[258])^(a[204] & b[259])^(a[203] & b[260])^(a[202] & b[261])^(a[201] & b[262])^(a[200] & b[263])^(a[199] & b[264])^(a[198] & b[265])^(a[197] & b[266])^(a[196] & b[267])^(a[195] & b[268])^(a[194] & b[269])^(a[193] & b[270])^(a[192] & b[271])^(a[191] & b[272])^(a[190] & b[273])^(a[189] & b[274])^(a[188] & b[275])^(a[187] & b[276])^(a[186] & b[277])^(a[185] & b[278])^(a[184] & b[279])^(a[183] & b[280])^(a[182] & b[281])^(a[181] & b[282])^(a[180] & b[283])^(a[179] & b[284])^(a[178] & b[285])^(a[177] & b[286])^(a[176] & b[287])^(a[175] & b[288])^(a[174] & b[289])^(a[173] & b[290])^(a[172] & b[291])^(a[171] & b[292])^(a[170] & b[293])^(a[169] & b[294])^(a[168] & b[295])^(a[167] & b[296])^(a[166] & b[297])^(a[165] & b[298])^(a[164] & b[299])^(a[163] & b[300])^(a[162] & b[301])^(a[161] & b[302])^(a[160] & b[303])^(a[159] & b[304])^(a[158] & b[305])^(a[157] & b[306])^(a[156] & b[307])^(a[155] & b[308])^(a[154] & b[309])^(a[153] & b[310])^(a[152] & b[311])^(a[151] & b[312])^(a[150] & b[313])^(a[149] & b[314])^(a[148] & b[315])^(a[147] & b[316])^(a[146] & b[317])^(a[145] & b[318])^(a[144] & b[319])^(a[143] & b[320])^(a[142] & b[321])^(a[141] & b[322])^(a[140] & b[323])^(a[139] & b[324])^(a[138] & b[325])^(a[137] & b[326])^(a[136] & b[327])^(a[135] & b[328])^(a[134] & b[329])^(a[133] & b[330])^(a[132] & b[331])^(a[131] & b[332])^(a[130] & b[333])^(a[129] & b[334])^(a[128] & b[335])^(a[127] & b[336])^(a[126] & b[337])^(a[125] & b[338])^(a[124] & b[339])^(a[123] & b[340])^(a[122] & b[341])^(a[121] & b[342])^(a[120] & b[343])^(a[119] & b[344])^(a[118] & b[345])^(a[117] & b[346])^(a[116] & b[347])^(a[115] & b[348])^(a[114] & b[349])^(a[113] & b[350])^(a[112] & b[351])^(a[111] & b[352])^(a[110] & b[353])^(a[109] & b[354])^(a[108] & b[355])^(a[107] & b[356])^(a[106] & b[357])^(a[105] & b[358])^(a[104] & b[359])^(a[103] & b[360])^(a[102] & b[361])^(a[101] & b[362])^(a[100] & b[363])^(a[99] & b[364])^(a[98] & b[365])^(a[97] & b[366])^(a[96] & b[367])^(a[95] & b[368])^(a[94] & b[369])^(a[93] & b[370])^(a[92] & b[371])^(a[91] & b[372])^(a[90] & b[373])^(a[89] & b[374])^(a[88] & b[375])^(a[87] & b[376])^(a[86] & b[377])^(a[85] & b[378])^(a[84] & b[379])^(a[83] & b[380])^(a[82] & b[381])^(a[81] & b[382])^(a[80] & b[383])^(a[79] & b[384])^(a[78] & b[385])^(a[77] & b[386])^(a[76] & b[387])^(a[75] & b[388])^(a[74] & b[389])^(a[73] & b[390])^(a[72] & b[391])^(a[71] & b[392])^(a[70] & b[393])^(a[69] & b[394])^(a[68] & b[395])^(a[67] & b[396])^(a[66] & b[397])^(a[65] & b[398])^(a[64] & b[399])^(a[63] & b[400])^(a[62] & b[401])^(a[61] & b[402])^(a[60] & b[403])^(a[59] & b[404])^(a[58] & b[405])^(a[57] & b[406])^(a[56] & b[407])^(a[55] & b[408]);
assign y[464] = (a[408] & b[56])^(a[407] & b[57])^(a[406] & b[58])^(a[405] & b[59])^(a[404] & b[60])^(a[403] & b[61])^(a[402] & b[62])^(a[401] & b[63])^(a[400] & b[64])^(a[399] & b[65])^(a[398] & b[66])^(a[397] & b[67])^(a[396] & b[68])^(a[395] & b[69])^(a[394] & b[70])^(a[393] & b[71])^(a[392] & b[72])^(a[391] & b[73])^(a[390] & b[74])^(a[389] & b[75])^(a[388] & b[76])^(a[387] & b[77])^(a[386] & b[78])^(a[385] & b[79])^(a[384] & b[80])^(a[383] & b[81])^(a[382] & b[82])^(a[381] & b[83])^(a[380] & b[84])^(a[379] & b[85])^(a[378] & b[86])^(a[377] & b[87])^(a[376] & b[88])^(a[375] & b[89])^(a[374] & b[90])^(a[373] & b[91])^(a[372] & b[92])^(a[371] & b[93])^(a[370] & b[94])^(a[369] & b[95])^(a[368] & b[96])^(a[367] & b[97])^(a[366] & b[98])^(a[365] & b[99])^(a[364] & b[100])^(a[363] & b[101])^(a[362] & b[102])^(a[361] & b[103])^(a[360] & b[104])^(a[359] & b[105])^(a[358] & b[106])^(a[357] & b[107])^(a[356] & b[108])^(a[355] & b[109])^(a[354] & b[110])^(a[353] & b[111])^(a[352] & b[112])^(a[351] & b[113])^(a[350] & b[114])^(a[349] & b[115])^(a[348] & b[116])^(a[347] & b[117])^(a[346] & b[118])^(a[345] & b[119])^(a[344] & b[120])^(a[343] & b[121])^(a[342] & b[122])^(a[341] & b[123])^(a[340] & b[124])^(a[339] & b[125])^(a[338] & b[126])^(a[337] & b[127])^(a[336] & b[128])^(a[335] & b[129])^(a[334] & b[130])^(a[333] & b[131])^(a[332] & b[132])^(a[331] & b[133])^(a[330] & b[134])^(a[329] & b[135])^(a[328] & b[136])^(a[327] & b[137])^(a[326] & b[138])^(a[325] & b[139])^(a[324] & b[140])^(a[323] & b[141])^(a[322] & b[142])^(a[321] & b[143])^(a[320] & b[144])^(a[319] & b[145])^(a[318] & b[146])^(a[317] & b[147])^(a[316] & b[148])^(a[315] & b[149])^(a[314] & b[150])^(a[313] & b[151])^(a[312] & b[152])^(a[311] & b[153])^(a[310] & b[154])^(a[309] & b[155])^(a[308] & b[156])^(a[307] & b[157])^(a[306] & b[158])^(a[305] & b[159])^(a[304] & b[160])^(a[303] & b[161])^(a[302] & b[162])^(a[301] & b[163])^(a[300] & b[164])^(a[299] & b[165])^(a[298] & b[166])^(a[297] & b[167])^(a[296] & b[168])^(a[295] & b[169])^(a[294] & b[170])^(a[293] & b[171])^(a[292] & b[172])^(a[291] & b[173])^(a[290] & b[174])^(a[289] & b[175])^(a[288] & b[176])^(a[287] & b[177])^(a[286] & b[178])^(a[285] & b[179])^(a[284] & b[180])^(a[283] & b[181])^(a[282] & b[182])^(a[281] & b[183])^(a[280] & b[184])^(a[279] & b[185])^(a[278] & b[186])^(a[277] & b[187])^(a[276] & b[188])^(a[275] & b[189])^(a[274] & b[190])^(a[273] & b[191])^(a[272] & b[192])^(a[271] & b[193])^(a[270] & b[194])^(a[269] & b[195])^(a[268] & b[196])^(a[267] & b[197])^(a[266] & b[198])^(a[265] & b[199])^(a[264] & b[200])^(a[263] & b[201])^(a[262] & b[202])^(a[261] & b[203])^(a[260] & b[204])^(a[259] & b[205])^(a[258] & b[206])^(a[257] & b[207])^(a[256] & b[208])^(a[255] & b[209])^(a[254] & b[210])^(a[253] & b[211])^(a[252] & b[212])^(a[251] & b[213])^(a[250] & b[214])^(a[249] & b[215])^(a[248] & b[216])^(a[247] & b[217])^(a[246] & b[218])^(a[245] & b[219])^(a[244] & b[220])^(a[243] & b[221])^(a[242] & b[222])^(a[241] & b[223])^(a[240] & b[224])^(a[239] & b[225])^(a[238] & b[226])^(a[237] & b[227])^(a[236] & b[228])^(a[235] & b[229])^(a[234] & b[230])^(a[233] & b[231])^(a[232] & b[232])^(a[231] & b[233])^(a[230] & b[234])^(a[229] & b[235])^(a[228] & b[236])^(a[227] & b[237])^(a[226] & b[238])^(a[225] & b[239])^(a[224] & b[240])^(a[223] & b[241])^(a[222] & b[242])^(a[221] & b[243])^(a[220] & b[244])^(a[219] & b[245])^(a[218] & b[246])^(a[217] & b[247])^(a[216] & b[248])^(a[215] & b[249])^(a[214] & b[250])^(a[213] & b[251])^(a[212] & b[252])^(a[211] & b[253])^(a[210] & b[254])^(a[209] & b[255])^(a[208] & b[256])^(a[207] & b[257])^(a[206] & b[258])^(a[205] & b[259])^(a[204] & b[260])^(a[203] & b[261])^(a[202] & b[262])^(a[201] & b[263])^(a[200] & b[264])^(a[199] & b[265])^(a[198] & b[266])^(a[197] & b[267])^(a[196] & b[268])^(a[195] & b[269])^(a[194] & b[270])^(a[193] & b[271])^(a[192] & b[272])^(a[191] & b[273])^(a[190] & b[274])^(a[189] & b[275])^(a[188] & b[276])^(a[187] & b[277])^(a[186] & b[278])^(a[185] & b[279])^(a[184] & b[280])^(a[183] & b[281])^(a[182] & b[282])^(a[181] & b[283])^(a[180] & b[284])^(a[179] & b[285])^(a[178] & b[286])^(a[177] & b[287])^(a[176] & b[288])^(a[175] & b[289])^(a[174] & b[290])^(a[173] & b[291])^(a[172] & b[292])^(a[171] & b[293])^(a[170] & b[294])^(a[169] & b[295])^(a[168] & b[296])^(a[167] & b[297])^(a[166] & b[298])^(a[165] & b[299])^(a[164] & b[300])^(a[163] & b[301])^(a[162] & b[302])^(a[161] & b[303])^(a[160] & b[304])^(a[159] & b[305])^(a[158] & b[306])^(a[157] & b[307])^(a[156] & b[308])^(a[155] & b[309])^(a[154] & b[310])^(a[153] & b[311])^(a[152] & b[312])^(a[151] & b[313])^(a[150] & b[314])^(a[149] & b[315])^(a[148] & b[316])^(a[147] & b[317])^(a[146] & b[318])^(a[145] & b[319])^(a[144] & b[320])^(a[143] & b[321])^(a[142] & b[322])^(a[141] & b[323])^(a[140] & b[324])^(a[139] & b[325])^(a[138] & b[326])^(a[137] & b[327])^(a[136] & b[328])^(a[135] & b[329])^(a[134] & b[330])^(a[133] & b[331])^(a[132] & b[332])^(a[131] & b[333])^(a[130] & b[334])^(a[129] & b[335])^(a[128] & b[336])^(a[127] & b[337])^(a[126] & b[338])^(a[125] & b[339])^(a[124] & b[340])^(a[123] & b[341])^(a[122] & b[342])^(a[121] & b[343])^(a[120] & b[344])^(a[119] & b[345])^(a[118] & b[346])^(a[117] & b[347])^(a[116] & b[348])^(a[115] & b[349])^(a[114] & b[350])^(a[113] & b[351])^(a[112] & b[352])^(a[111] & b[353])^(a[110] & b[354])^(a[109] & b[355])^(a[108] & b[356])^(a[107] & b[357])^(a[106] & b[358])^(a[105] & b[359])^(a[104] & b[360])^(a[103] & b[361])^(a[102] & b[362])^(a[101] & b[363])^(a[100] & b[364])^(a[99] & b[365])^(a[98] & b[366])^(a[97] & b[367])^(a[96] & b[368])^(a[95] & b[369])^(a[94] & b[370])^(a[93] & b[371])^(a[92] & b[372])^(a[91] & b[373])^(a[90] & b[374])^(a[89] & b[375])^(a[88] & b[376])^(a[87] & b[377])^(a[86] & b[378])^(a[85] & b[379])^(a[84] & b[380])^(a[83] & b[381])^(a[82] & b[382])^(a[81] & b[383])^(a[80] & b[384])^(a[79] & b[385])^(a[78] & b[386])^(a[77] & b[387])^(a[76] & b[388])^(a[75] & b[389])^(a[74] & b[390])^(a[73] & b[391])^(a[72] & b[392])^(a[71] & b[393])^(a[70] & b[394])^(a[69] & b[395])^(a[68] & b[396])^(a[67] & b[397])^(a[66] & b[398])^(a[65] & b[399])^(a[64] & b[400])^(a[63] & b[401])^(a[62] & b[402])^(a[61] & b[403])^(a[60] & b[404])^(a[59] & b[405])^(a[58] & b[406])^(a[57] & b[407])^(a[56] & b[408]);
assign y[465] = (a[408] & b[57])^(a[407] & b[58])^(a[406] & b[59])^(a[405] & b[60])^(a[404] & b[61])^(a[403] & b[62])^(a[402] & b[63])^(a[401] & b[64])^(a[400] & b[65])^(a[399] & b[66])^(a[398] & b[67])^(a[397] & b[68])^(a[396] & b[69])^(a[395] & b[70])^(a[394] & b[71])^(a[393] & b[72])^(a[392] & b[73])^(a[391] & b[74])^(a[390] & b[75])^(a[389] & b[76])^(a[388] & b[77])^(a[387] & b[78])^(a[386] & b[79])^(a[385] & b[80])^(a[384] & b[81])^(a[383] & b[82])^(a[382] & b[83])^(a[381] & b[84])^(a[380] & b[85])^(a[379] & b[86])^(a[378] & b[87])^(a[377] & b[88])^(a[376] & b[89])^(a[375] & b[90])^(a[374] & b[91])^(a[373] & b[92])^(a[372] & b[93])^(a[371] & b[94])^(a[370] & b[95])^(a[369] & b[96])^(a[368] & b[97])^(a[367] & b[98])^(a[366] & b[99])^(a[365] & b[100])^(a[364] & b[101])^(a[363] & b[102])^(a[362] & b[103])^(a[361] & b[104])^(a[360] & b[105])^(a[359] & b[106])^(a[358] & b[107])^(a[357] & b[108])^(a[356] & b[109])^(a[355] & b[110])^(a[354] & b[111])^(a[353] & b[112])^(a[352] & b[113])^(a[351] & b[114])^(a[350] & b[115])^(a[349] & b[116])^(a[348] & b[117])^(a[347] & b[118])^(a[346] & b[119])^(a[345] & b[120])^(a[344] & b[121])^(a[343] & b[122])^(a[342] & b[123])^(a[341] & b[124])^(a[340] & b[125])^(a[339] & b[126])^(a[338] & b[127])^(a[337] & b[128])^(a[336] & b[129])^(a[335] & b[130])^(a[334] & b[131])^(a[333] & b[132])^(a[332] & b[133])^(a[331] & b[134])^(a[330] & b[135])^(a[329] & b[136])^(a[328] & b[137])^(a[327] & b[138])^(a[326] & b[139])^(a[325] & b[140])^(a[324] & b[141])^(a[323] & b[142])^(a[322] & b[143])^(a[321] & b[144])^(a[320] & b[145])^(a[319] & b[146])^(a[318] & b[147])^(a[317] & b[148])^(a[316] & b[149])^(a[315] & b[150])^(a[314] & b[151])^(a[313] & b[152])^(a[312] & b[153])^(a[311] & b[154])^(a[310] & b[155])^(a[309] & b[156])^(a[308] & b[157])^(a[307] & b[158])^(a[306] & b[159])^(a[305] & b[160])^(a[304] & b[161])^(a[303] & b[162])^(a[302] & b[163])^(a[301] & b[164])^(a[300] & b[165])^(a[299] & b[166])^(a[298] & b[167])^(a[297] & b[168])^(a[296] & b[169])^(a[295] & b[170])^(a[294] & b[171])^(a[293] & b[172])^(a[292] & b[173])^(a[291] & b[174])^(a[290] & b[175])^(a[289] & b[176])^(a[288] & b[177])^(a[287] & b[178])^(a[286] & b[179])^(a[285] & b[180])^(a[284] & b[181])^(a[283] & b[182])^(a[282] & b[183])^(a[281] & b[184])^(a[280] & b[185])^(a[279] & b[186])^(a[278] & b[187])^(a[277] & b[188])^(a[276] & b[189])^(a[275] & b[190])^(a[274] & b[191])^(a[273] & b[192])^(a[272] & b[193])^(a[271] & b[194])^(a[270] & b[195])^(a[269] & b[196])^(a[268] & b[197])^(a[267] & b[198])^(a[266] & b[199])^(a[265] & b[200])^(a[264] & b[201])^(a[263] & b[202])^(a[262] & b[203])^(a[261] & b[204])^(a[260] & b[205])^(a[259] & b[206])^(a[258] & b[207])^(a[257] & b[208])^(a[256] & b[209])^(a[255] & b[210])^(a[254] & b[211])^(a[253] & b[212])^(a[252] & b[213])^(a[251] & b[214])^(a[250] & b[215])^(a[249] & b[216])^(a[248] & b[217])^(a[247] & b[218])^(a[246] & b[219])^(a[245] & b[220])^(a[244] & b[221])^(a[243] & b[222])^(a[242] & b[223])^(a[241] & b[224])^(a[240] & b[225])^(a[239] & b[226])^(a[238] & b[227])^(a[237] & b[228])^(a[236] & b[229])^(a[235] & b[230])^(a[234] & b[231])^(a[233] & b[232])^(a[232] & b[233])^(a[231] & b[234])^(a[230] & b[235])^(a[229] & b[236])^(a[228] & b[237])^(a[227] & b[238])^(a[226] & b[239])^(a[225] & b[240])^(a[224] & b[241])^(a[223] & b[242])^(a[222] & b[243])^(a[221] & b[244])^(a[220] & b[245])^(a[219] & b[246])^(a[218] & b[247])^(a[217] & b[248])^(a[216] & b[249])^(a[215] & b[250])^(a[214] & b[251])^(a[213] & b[252])^(a[212] & b[253])^(a[211] & b[254])^(a[210] & b[255])^(a[209] & b[256])^(a[208] & b[257])^(a[207] & b[258])^(a[206] & b[259])^(a[205] & b[260])^(a[204] & b[261])^(a[203] & b[262])^(a[202] & b[263])^(a[201] & b[264])^(a[200] & b[265])^(a[199] & b[266])^(a[198] & b[267])^(a[197] & b[268])^(a[196] & b[269])^(a[195] & b[270])^(a[194] & b[271])^(a[193] & b[272])^(a[192] & b[273])^(a[191] & b[274])^(a[190] & b[275])^(a[189] & b[276])^(a[188] & b[277])^(a[187] & b[278])^(a[186] & b[279])^(a[185] & b[280])^(a[184] & b[281])^(a[183] & b[282])^(a[182] & b[283])^(a[181] & b[284])^(a[180] & b[285])^(a[179] & b[286])^(a[178] & b[287])^(a[177] & b[288])^(a[176] & b[289])^(a[175] & b[290])^(a[174] & b[291])^(a[173] & b[292])^(a[172] & b[293])^(a[171] & b[294])^(a[170] & b[295])^(a[169] & b[296])^(a[168] & b[297])^(a[167] & b[298])^(a[166] & b[299])^(a[165] & b[300])^(a[164] & b[301])^(a[163] & b[302])^(a[162] & b[303])^(a[161] & b[304])^(a[160] & b[305])^(a[159] & b[306])^(a[158] & b[307])^(a[157] & b[308])^(a[156] & b[309])^(a[155] & b[310])^(a[154] & b[311])^(a[153] & b[312])^(a[152] & b[313])^(a[151] & b[314])^(a[150] & b[315])^(a[149] & b[316])^(a[148] & b[317])^(a[147] & b[318])^(a[146] & b[319])^(a[145] & b[320])^(a[144] & b[321])^(a[143] & b[322])^(a[142] & b[323])^(a[141] & b[324])^(a[140] & b[325])^(a[139] & b[326])^(a[138] & b[327])^(a[137] & b[328])^(a[136] & b[329])^(a[135] & b[330])^(a[134] & b[331])^(a[133] & b[332])^(a[132] & b[333])^(a[131] & b[334])^(a[130] & b[335])^(a[129] & b[336])^(a[128] & b[337])^(a[127] & b[338])^(a[126] & b[339])^(a[125] & b[340])^(a[124] & b[341])^(a[123] & b[342])^(a[122] & b[343])^(a[121] & b[344])^(a[120] & b[345])^(a[119] & b[346])^(a[118] & b[347])^(a[117] & b[348])^(a[116] & b[349])^(a[115] & b[350])^(a[114] & b[351])^(a[113] & b[352])^(a[112] & b[353])^(a[111] & b[354])^(a[110] & b[355])^(a[109] & b[356])^(a[108] & b[357])^(a[107] & b[358])^(a[106] & b[359])^(a[105] & b[360])^(a[104] & b[361])^(a[103] & b[362])^(a[102] & b[363])^(a[101] & b[364])^(a[100] & b[365])^(a[99] & b[366])^(a[98] & b[367])^(a[97] & b[368])^(a[96] & b[369])^(a[95] & b[370])^(a[94] & b[371])^(a[93] & b[372])^(a[92] & b[373])^(a[91] & b[374])^(a[90] & b[375])^(a[89] & b[376])^(a[88] & b[377])^(a[87] & b[378])^(a[86] & b[379])^(a[85] & b[380])^(a[84] & b[381])^(a[83] & b[382])^(a[82] & b[383])^(a[81] & b[384])^(a[80] & b[385])^(a[79] & b[386])^(a[78] & b[387])^(a[77] & b[388])^(a[76] & b[389])^(a[75] & b[390])^(a[74] & b[391])^(a[73] & b[392])^(a[72] & b[393])^(a[71] & b[394])^(a[70] & b[395])^(a[69] & b[396])^(a[68] & b[397])^(a[67] & b[398])^(a[66] & b[399])^(a[65] & b[400])^(a[64] & b[401])^(a[63] & b[402])^(a[62] & b[403])^(a[61] & b[404])^(a[60] & b[405])^(a[59] & b[406])^(a[58] & b[407])^(a[57] & b[408]);
assign y[466] = (a[408] & b[58])^(a[407] & b[59])^(a[406] & b[60])^(a[405] & b[61])^(a[404] & b[62])^(a[403] & b[63])^(a[402] & b[64])^(a[401] & b[65])^(a[400] & b[66])^(a[399] & b[67])^(a[398] & b[68])^(a[397] & b[69])^(a[396] & b[70])^(a[395] & b[71])^(a[394] & b[72])^(a[393] & b[73])^(a[392] & b[74])^(a[391] & b[75])^(a[390] & b[76])^(a[389] & b[77])^(a[388] & b[78])^(a[387] & b[79])^(a[386] & b[80])^(a[385] & b[81])^(a[384] & b[82])^(a[383] & b[83])^(a[382] & b[84])^(a[381] & b[85])^(a[380] & b[86])^(a[379] & b[87])^(a[378] & b[88])^(a[377] & b[89])^(a[376] & b[90])^(a[375] & b[91])^(a[374] & b[92])^(a[373] & b[93])^(a[372] & b[94])^(a[371] & b[95])^(a[370] & b[96])^(a[369] & b[97])^(a[368] & b[98])^(a[367] & b[99])^(a[366] & b[100])^(a[365] & b[101])^(a[364] & b[102])^(a[363] & b[103])^(a[362] & b[104])^(a[361] & b[105])^(a[360] & b[106])^(a[359] & b[107])^(a[358] & b[108])^(a[357] & b[109])^(a[356] & b[110])^(a[355] & b[111])^(a[354] & b[112])^(a[353] & b[113])^(a[352] & b[114])^(a[351] & b[115])^(a[350] & b[116])^(a[349] & b[117])^(a[348] & b[118])^(a[347] & b[119])^(a[346] & b[120])^(a[345] & b[121])^(a[344] & b[122])^(a[343] & b[123])^(a[342] & b[124])^(a[341] & b[125])^(a[340] & b[126])^(a[339] & b[127])^(a[338] & b[128])^(a[337] & b[129])^(a[336] & b[130])^(a[335] & b[131])^(a[334] & b[132])^(a[333] & b[133])^(a[332] & b[134])^(a[331] & b[135])^(a[330] & b[136])^(a[329] & b[137])^(a[328] & b[138])^(a[327] & b[139])^(a[326] & b[140])^(a[325] & b[141])^(a[324] & b[142])^(a[323] & b[143])^(a[322] & b[144])^(a[321] & b[145])^(a[320] & b[146])^(a[319] & b[147])^(a[318] & b[148])^(a[317] & b[149])^(a[316] & b[150])^(a[315] & b[151])^(a[314] & b[152])^(a[313] & b[153])^(a[312] & b[154])^(a[311] & b[155])^(a[310] & b[156])^(a[309] & b[157])^(a[308] & b[158])^(a[307] & b[159])^(a[306] & b[160])^(a[305] & b[161])^(a[304] & b[162])^(a[303] & b[163])^(a[302] & b[164])^(a[301] & b[165])^(a[300] & b[166])^(a[299] & b[167])^(a[298] & b[168])^(a[297] & b[169])^(a[296] & b[170])^(a[295] & b[171])^(a[294] & b[172])^(a[293] & b[173])^(a[292] & b[174])^(a[291] & b[175])^(a[290] & b[176])^(a[289] & b[177])^(a[288] & b[178])^(a[287] & b[179])^(a[286] & b[180])^(a[285] & b[181])^(a[284] & b[182])^(a[283] & b[183])^(a[282] & b[184])^(a[281] & b[185])^(a[280] & b[186])^(a[279] & b[187])^(a[278] & b[188])^(a[277] & b[189])^(a[276] & b[190])^(a[275] & b[191])^(a[274] & b[192])^(a[273] & b[193])^(a[272] & b[194])^(a[271] & b[195])^(a[270] & b[196])^(a[269] & b[197])^(a[268] & b[198])^(a[267] & b[199])^(a[266] & b[200])^(a[265] & b[201])^(a[264] & b[202])^(a[263] & b[203])^(a[262] & b[204])^(a[261] & b[205])^(a[260] & b[206])^(a[259] & b[207])^(a[258] & b[208])^(a[257] & b[209])^(a[256] & b[210])^(a[255] & b[211])^(a[254] & b[212])^(a[253] & b[213])^(a[252] & b[214])^(a[251] & b[215])^(a[250] & b[216])^(a[249] & b[217])^(a[248] & b[218])^(a[247] & b[219])^(a[246] & b[220])^(a[245] & b[221])^(a[244] & b[222])^(a[243] & b[223])^(a[242] & b[224])^(a[241] & b[225])^(a[240] & b[226])^(a[239] & b[227])^(a[238] & b[228])^(a[237] & b[229])^(a[236] & b[230])^(a[235] & b[231])^(a[234] & b[232])^(a[233] & b[233])^(a[232] & b[234])^(a[231] & b[235])^(a[230] & b[236])^(a[229] & b[237])^(a[228] & b[238])^(a[227] & b[239])^(a[226] & b[240])^(a[225] & b[241])^(a[224] & b[242])^(a[223] & b[243])^(a[222] & b[244])^(a[221] & b[245])^(a[220] & b[246])^(a[219] & b[247])^(a[218] & b[248])^(a[217] & b[249])^(a[216] & b[250])^(a[215] & b[251])^(a[214] & b[252])^(a[213] & b[253])^(a[212] & b[254])^(a[211] & b[255])^(a[210] & b[256])^(a[209] & b[257])^(a[208] & b[258])^(a[207] & b[259])^(a[206] & b[260])^(a[205] & b[261])^(a[204] & b[262])^(a[203] & b[263])^(a[202] & b[264])^(a[201] & b[265])^(a[200] & b[266])^(a[199] & b[267])^(a[198] & b[268])^(a[197] & b[269])^(a[196] & b[270])^(a[195] & b[271])^(a[194] & b[272])^(a[193] & b[273])^(a[192] & b[274])^(a[191] & b[275])^(a[190] & b[276])^(a[189] & b[277])^(a[188] & b[278])^(a[187] & b[279])^(a[186] & b[280])^(a[185] & b[281])^(a[184] & b[282])^(a[183] & b[283])^(a[182] & b[284])^(a[181] & b[285])^(a[180] & b[286])^(a[179] & b[287])^(a[178] & b[288])^(a[177] & b[289])^(a[176] & b[290])^(a[175] & b[291])^(a[174] & b[292])^(a[173] & b[293])^(a[172] & b[294])^(a[171] & b[295])^(a[170] & b[296])^(a[169] & b[297])^(a[168] & b[298])^(a[167] & b[299])^(a[166] & b[300])^(a[165] & b[301])^(a[164] & b[302])^(a[163] & b[303])^(a[162] & b[304])^(a[161] & b[305])^(a[160] & b[306])^(a[159] & b[307])^(a[158] & b[308])^(a[157] & b[309])^(a[156] & b[310])^(a[155] & b[311])^(a[154] & b[312])^(a[153] & b[313])^(a[152] & b[314])^(a[151] & b[315])^(a[150] & b[316])^(a[149] & b[317])^(a[148] & b[318])^(a[147] & b[319])^(a[146] & b[320])^(a[145] & b[321])^(a[144] & b[322])^(a[143] & b[323])^(a[142] & b[324])^(a[141] & b[325])^(a[140] & b[326])^(a[139] & b[327])^(a[138] & b[328])^(a[137] & b[329])^(a[136] & b[330])^(a[135] & b[331])^(a[134] & b[332])^(a[133] & b[333])^(a[132] & b[334])^(a[131] & b[335])^(a[130] & b[336])^(a[129] & b[337])^(a[128] & b[338])^(a[127] & b[339])^(a[126] & b[340])^(a[125] & b[341])^(a[124] & b[342])^(a[123] & b[343])^(a[122] & b[344])^(a[121] & b[345])^(a[120] & b[346])^(a[119] & b[347])^(a[118] & b[348])^(a[117] & b[349])^(a[116] & b[350])^(a[115] & b[351])^(a[114] & b[352])^(a[113] & b[353])^(a[112] & b[354])^(a[111] & b[355])^(a[110] & b[356])^(a[109] & b[357])^(a[108] & b[358])^(a[107] & b[359])^(a[106] & b[360])^(a[105] & b[361])^(a[104] & b[362])^(a[103] & b[363])^(a[102] & b[364])^(a[101] & b[365])^(a[100] & b[366])^(a[99] & b[367])^(a[98] & b[368])^(a[97] & b[369])^(a[96] & b[370])^(a[95] & b[371])^(a[94] & b[372])^(a[93] & b[373])^(a[92] & b[374])^(a[91] & b[375])^(a[90] & b[376])^(a[89] & b[377])^(a[88] & b[378])^(a[87] & b[379])^(a[86] & b[380])^(a[85] & b[381])^(a[84] & b[382])^(a[83] & b[383])^(a[82] & b[384])^(a[81] & b[385])^(a[80] & b[386])^(a[79] & b[387])^(a[78] & b[388])^(a[77] & b[389])^(a[76] & b[390])^(a[75] & b[391])^(a[74] & b[392])^(a[73] & b[393])^(a[72] & b[394])^(a[71] & b[395])^(a[70] & b[396])^(a[69] & b[397])^(a[68] & b[398])^(a[67] & b[399])^(a[66] & b[400])^(a[65] & b[401])^(a[64] & b[402])^(a[63] & b[403])^(a[62] & b[404])^(a[61] & b[405])^(a[60] & b[406])^(a[59] & b[407])^(a[58] & b[408]);
assign y[467] = (a[408] & b[59])^(a[407] & b[60])^(a[406] & b[61])^(a[405] & b[62])^(a[404] & b[63])^(a[403] & b[64])^(a[402] & b[65])^(a[401] & b[66])^(a[400] & b[67])^(a[399] & b[68])^(a[398] & b[69])^(a[397] & b[70])^(a[396] & b[71])^(a[395] & b[72])^(a[394] & b[73])^(a[393] & b[74])^(a[392] & b[75])^(a[391] & b[76])^(a[390] & b[77])^(a[389] & b[78])^(a[388] & b[79])^(a[387] & b[80])^(a[386] & b[81])^(a[385] & b[82])^(a[384] & b[83])^(a[383] & b[84])^(a[382] & b[85])^(a[381] & b[86])^(a[380] & b[87])^(a[379] & b[88])^(a[378] & b[89])^(a[377] & b[90])^(a[376] & b[91])^(a[375] & b[92])^(a[374] & b[93])^(a[373] & b[94])^(a[372] & b[95])^(a[371] & b[96])^(a[370] & b[97])^(a[369] & b[98])^(a[368] & b[99])^(a[367] & b[100])^(a[366] & b[101])^(a[365] & b[102])^(a[364] & b[103])^(a[363] & b[104])^(a[362] & b[105])^(a[361] & b[106])^(a[360] & b[107])^(a[359] & b[108])^(a[358] & b[109])^(a[357] & b[110])^(a[356] & b[111])^(a[355] & b[112])^(a[354] & b[113])^(a[353] & b[114])^(a[352] & b[115])^(a[351] & b[116])^(a[350] & b[117])^(a[349] & b[118])^(a[348] & b[119])^(a[347] & b[120])^(a[346] & b[121])^(a[345] & b[122])^(a[344] & b[123])^(a[343] & b[124])^(a[342] & b[125])^(a[341] & b[126])^(a[340] & b[127])^(a[339] & b[128])^(a[338] & b[129])^(a[337] & b[130])^(a[336] & b[131])^(a[335] & b[132])^(a[334] & b[133])^(a[333] & b[134])^(a[332] & b[135])^(a[331] & b[136])^(a[330] & b[137])^(a[329] & b[138])^(a[328] & b[139])^(a[327] & b[140])^(a[326] & b[141])^(a[325] & b[142])^(a[324] & b[143])^(a[323] & b[144])^(a[322] & b[145])^(a[321] & b[146])^(a[320] & b[147])^(a[319] & b[148])^(a[318] & b[149])^(a[317] & b[150])^(a[316] & b[151])^(a[315] & b[152])^(a[314] & b[153])^(a[313] & b[154])^(a[312] & b[155])^(a[311] & b[156])^(a[310] & b[157])^(a[309] & b[158])^(a[308] & b[159])^(a[307] & b[160])^(a[306] & b[161])^(a[305] & b[162])^(a[304] & b[163])^(a[303] & b[164])^(a[302] & b[165])^(a[301] & b[166])^(a[300] & b[167])^(a[299] & b[168])^(a[298] & b[169])^(a[297] & b[170])^(a[296] & b[171])^(a[295] & b[172])^(a[294] & b[173])^(a[293] & b[174])^(a[292] & b[175])^(a[291] & b[176])^(a[290] & b[177])^(a[289] & b[178])^(a[288] & b[179])^(a[287] & b[180])^(a[286] & b[181])^(a[285] & b[182])^(a[284] & b[183])^(a[283] & b[184])^(a[282] & b[185])^(a[281] & b[186])^(a[280] & b[187])^(a[279] & b[188])^(a[278] & b[189])^(a[277] & b[190])^(a[276] & b[191])^(a[275] & b[192])^(a[274] & b[193])^(a[273] & b[194])^(a[272] & b[195])^(a[271] & b[196])^(a[270] & b[197])^(a[269] & b[198])^(a[268] & b[199])^(a[267] & b[200])^(a[266] & b[201])^(a[265] & b[202])^(a[264] & b[203])^(a[263] & b[204])^(a[262] & b[205])^(a[261] & b[206])^(a[260] & b[207])^(a[259] & b[208])^(a[258] & b[209])^(a[257] & b[210])^(a[256] & b[211])^(a[255] & b[212])^(a[254] & b[213])^(a[253] & b[214])^(a[252] & b[215])^(a[251] & b[216])^(a[250] & b[217])^(a[249] & b[218])^(a[248] & b[219])^(a[247] & b[220])^(a[246] & b[221])^(a[245] & b[222])^(a[244] & b[223])^(a[243] & b[224])^(a[242] & b[225])^(a[241] & b[226])^(a[240] & b[227])^(a[239] & b[228])^(a[238] & b[229])^(a[237] & b[230])^(a[236] & b[231])^(a[235] & b[232])^(a[234] & b[233])^(a[233] & b[234])^(a[232] & b[235])^(a[231] & b[236])^(a[230] & b[237])^(a[229] & b[238])^(a[228] & b[239])^(a[227] & b[240])^(a[226] & b[241])^(a[225] & b[242])^(a[224] & b[243])^(a[223] & b[244])^(a[222] & b[245])^(a[221] & b[246])^(a[220] & b[247])^(a[219] & b[248])^(a[218] & b[249])^(a[217] & b[250])^(a[216] & b[251])^(a[215] & b[252])^(a[214] & b[253])^(a[213] & b[254])^(a[212] & b[255])^(a[211] & b[256])^(a[210] & b[257])^(a[209] & b[258])^(a[208] & b[259])^(a[207] & b[260])^(a[206] & b[261])^(a[205] & b[262])^(a[204] & b[263])^(a[203] & b[264])^(a[202] & b[265])^(a[201] & b[266])^(a[200] & b[267])^(a[199] & b[268])^(a[198] & b[269])^(a[197] & b[270])^(a[196] & b[271])^(a[195] & b[272])^(a[194] & b[273])^(a[193] & b[274])^(a[192] & b[275])^(a[191] & b[276])^(a[190] & b[277])^(a[189] & b[278])^(a[188] & b[279])^(a[187] & b[280])^(a[186] & b[281])^(a[185] & b[282])^(a[184] & b[283])^(a[183] & b[284])^(a[182] & b[285])^(a[181] & b[286])^(a[180] & b[287])^(a[179] & b[288])^(a[178] & b[289])^(a[177] & b[290])^(a[176] & b[291])^(a[175] & b[292])^(a[174] & b[293])^(a[173] & b[294])^(a[172] & b[295])^(a[171] & b[296])^(a[170] & b[297])^(a[169] & b[298])^(a[168] & b[299])^(a[167] & b[300])^(a[166] & b[301])^(a[165] & b[302])^(a[164] & b[303])^(a[163] & b[304])^(a[162] & b[305])^(a[161] & b[306])^(a[160] & b[307])^(a[159] & b[308])^(a[158] & b[309])^(a[157] & b[310])^(a[156] & b[311])^(a[155] & b[312])^(a[154] & b[313])^(a[153] & b[314])^(a[152] & b[315])^(a[151] & b[316])^(a[150] & b[317])^(a[149] & b[318])^(a[148] & b[319])^(a[147] & b[320])^(a[146] & b[321])^(a[145] & b[322])^(a[144] & b[323])^(a[143] & b[324])^(a[142] & b[325])^(a[141] & b[326])^(a[140] & b[327])^(a[139] & b[328])^(a[138] & b[329])^(a[137] & b[330])^(a[136] & b[331])^(a[135] & b[332])^(a[134] & b[333])^(a[133] & b[334])^(a[132] & b[335])^(a[131] & b[336])^(a[130] & b[337])^(a[129] & b[338])^(a[128] & b[339])^(a[127] & b[340])^(a[126] & b[341])^(a[125] & b[342])^(a[124] & b[343])^(a[123] & b[344])^(a[122] & b[345])^(a[121] & b[346])^(a[120] & b[347])^(a[119] & b[348])^(a[118] & b[349])^(a[117] & b[350])^(a[116] & b[351])^(a[115] & b[352])^(a[114] & b[353])^(a[113] & b[354])^(a[112] & b[355])^(a[111] & b[356])^(a[110] & b[357])^(a[109] & b[358])^(a[108] & b[359])^(a[107] & b[360])^(a[106] & b[361])^(a[105] & b[362])^(a[104] & b[363])^(a[103] & b[364])^(a[102] & b[365])^(a[101] & b[366])^(a[100] & b[367])^(a[99] & b[368])^(a[98] & b[369])^(a[97] & b[370])^(a[96] & b[371])^(a[95] & b[372])^(a[94] & b[373])^(a[93] & b[374])^(a[92] & b[375])^(a[91] & b[376])^(a[90] & b[377])^(a[89] & b[378])^(a[88] & b[379])^(a[87] & b[380])^(a[86] & b[381])^(a[85] & b[382])^(a[84] & b[383])^(a[83] & b[384])^(a[82] & b[385])^(a[81] & b[386])^(a[80] & b[387])^(a[79] & b[388])^(a[78] & b[389])^(a[77] & b[390])^(a[76] & b[391])^(a[75] & b[392])^(a[74] & b[393])^(a[73] & b[394])^(a[72] & b[395])^(a[71] & b[396])^(a[70] & b[397])^(a[69] & b[398])^(a[68] & b[399])^(a[67] & b[400])^(a[66] & b[401])^(a[65] & b[402])^(a[64] & b[403])^(a[63] & b[404])^(a[62] & b[405])^(a[61] & b[406])^(a[60] & b[407])^(a[59] & b[408]);
assign y[468] = (a[408] & b[60])^(a[407] & b[61])^(a[406] & b[62])^(a[405] & b[63])^(a[404] & b[64])^(a[403] & b[65])^(a[402] & b[66])^(a[401] & b[67])^(a[400] & b[68])^(a[399] & b[69])^(a[398] & b[70])^(a[397] & b[71])^(a[396] & b[72])^(a[395] & b[73])^(a[394] & b[74])^(a[393] & b[75])^(a[392] & b[76])^(a[391] & b[77])^(a[390] & b[78])^(a[389] & b[79])^(a[388] & b[80])^(a[387] & b[81])^(a[386] & b[82])^(a[385] & b[83])^(a[384] & b[84])^(a[383] & b[85])^(a[382] & b[86])^(a[381] & b[87])^(a[380] & b[88])^(a[379] & b[89])^(a[378] & b[90])^(a[377] & b[91])^(a[376] & b[92])^(a[375] & b[93])^(a[374] & b[94])^(a[373] & b[95])^(a[372] & b[96])^(a[371] & b[97])^(a[370] & b[98])^(a[369] & b[99])^(a[368] & b[100])^(a[367] & b[101])^(a[366] & b[102])^(a[365] & b[103])^(a[364] & b[104])^(a[363] & b[105])^(a[362] & b[106])^(a[361] & b[107])^(a[360] & b[108])^(a[359] & b[109])^(a[358] & b[110])^(a[357] & b[111])^(a[356] & b[112])^(a[355] & b[113])^(a[354] & b[114])^(a[353] & b[115])^(a[352] & b[116])^(a[351] & b[117])^(a[350] & b[118])^(a[349] & b[119])^(a[348] & b[120])^(a[347] & b[121])^(a[346] & b[122])^(a[345] & b[123])^(a[344] & b[124])^(a[343] & b[125])^(a[342] & b[126])^(a[341] & b[127])^(a[340] & b[128])^(a[339] & b[129])^(a[338] & b[130])^(a[337] & b[131])^(a[336] & b[132])^(a[335] & b[133])^(a[334] & b[134])^(a[333] & b[135])^(a[332] & b[136])^(a[331] & b[137])^(a[330] & b[138])^(a[329] & b[139])^(a[328] & b[140])^(a[327] & b[141])^(a[326] & b[142])^(a[325] & b[143])^(a[324] & b[144])^(a[323] & b[145])^(a[322] & b[146])^(a[321] & b[147])^(a[320] & b[148])^(a[319] & b[149])^(a[318] & b[150])^(a[317] & b[151])^(a[316] & b[152])^(a[315] & b[153])^(a[314] & b[154])^(a[313] & b[155])^(a[312] & b[156])^(a[311] & b[157])^(a[310] & b[158])^(a[309] & b[159])^(a[308] & b[160])^(a[307] & b[161])^(a[306] & b[162])^(a[305] & b[163])^(a[304] & b[164])^(a[303] & b[165])^(a[302] & b[166])^(a[301] & b[167])^(a[300] & b[168])^(a[299] & b[169])^(a[298] & b[170])^(a[297] & b[171])^(a[296] & b[172])^(a[295] & b[173])^(a[294] & b[174])^(a[293] & b[175])^(a[292] & b[176])^(a[291] & b[177])^(a[290] & b[178])^(a[289] & b[179])^(a[288] & b[180])^(a[287] & b[181])^(a[286] & b[182])^(a[285] & b[183])^(a[284] & b[184])^(a[283] & b[185])^(a[282] & b[186])^(a[281] & b[187])^(a[280] & b[188])^(a[279] & b[189])^(a[278] & b[190])^(a[277] & b[191])^(a[276] & b[192])^(a[275] & b[193])^(a[274] & b[194])^(a[273] & b[195])^(a[272] & b[196])^(a[271] & b[197])^(a[270] & b[198])^(a[269] & b[199])^(a[268] & b[200])^(a[267] & b[201])^(a[266] & b[202])^(a[265] & b[203])^(a[264] & b[204])^(a[263] & b[205])^(a[262] & b[206])^(a[261] & b[207])^(a[260] & b[208])^(a[259] & b[209])^(a[258] & b[210])^(a[257] & b[211])^(a[256] & b[212])^(a[255] & b[213])^(a[254] & b[214])^(a[253] & b[215])^(a[252] & b[216])^(a[251] & b[217])^(a[250] & b[218])^(a[249] & b[219])^(a[248] & b[220])^(a[247] & b[221])^(a[246] & b[222])^(a[245] & b[223])^(a[244] & b[224])^(a[243] & b[225])^(a[242] & b[226])^(a[241] & b[227])^(a[240] & b[228])^(a[239] & b[229])^(a[238] & b[230])^(a[237] & b[231])^(a[236] & b[232])^(a[235] & b[233])^(a[234] & b[234])^(a[233] & b[235])^(a[232] & b[236])^(a[231] & b[237])^(a[230] & b[238])^(a[229] & b[239])^(a[228] & b[240])^(a[227] & b[241])^(a[226] & b[242])^(a[225] & b[243])^(a[224] & b[244])^(a[223] & b[245])^(a[222] & b[246])^(a[221] & b[247])^(a[220] & b[248])^(a[219] & b[249])^(a[218] & b[250])^(a[217] & b[251])^(a[216] & b[252])^(a[215] & b[253])^(a[214] & b[254])^(a[213] & b[255])^(a[212] & b[256])^(a[211] & b[257])^(a[210] & b[258])^(a[209] & b[259])^(a[208] & b[260])^(a[207] & b[261])^(a[206] & b[262])^(a[205] & b[263])^(a[204] & b[264])^(a[203] & b[265])^(a[202] & b[266])^(a[201] & b[267])^(a[200] & b[268])^(a[199] & b[269])^(a[198] & b[270])^(a[197] & b[271])^(a[196] & b[272])^(a[195] & b[273])^(a[194] & b[274])^(a[193] & b[275])^(a[192] & b[276])^(a[191] & b[277])^(a[190] & b[278])^(a[189] & b[279])^(a[188] & b[280])^(a[187] & b[281])^(a[186] & b[282])^(a[185] & b[283])^(a[184] & b[284])^(a[183] & b[285])^(a[182] & b[286])^(a[181] & b[287])^(a[180] & b[288])^(a[179] & b[289])^(a[178] & b[290])^(a[177] & b[291])^(a[176] & b[292])^(a[175] & b[293])^(a[174] & b[294])^(a[173] & b[295])^(a[172] & b[296])^(a[171] & b[297])^(a[170] & b[298])^(a[169] & b[299])^(a[168] & b[300])^(a[167] & b[301])^(a[166] & b[302])^(a[165] & b[303])^(a[164] & b[304])^(a[163] & b[305])^(a[162] & b[306])^(a[161] & b[307])^(a[160] & b[308])^(a[159] & b[309])^(a[158] & b[310])^(a[157] & b[311])^(a[156] & b[312])^(a[155] & b[313])^(a[154] & b[314])^(a[153] & b[315])^(a[152] & b[316])^(a[151] & b[317])^(a[150] & b[318])^(a[149] & b[319])^(a[148] & b[320])^(a[147] & b[321])^(a[146] & b[322])^(a[145] & b[323])^(a[144] & b[324])^(a[143] & b[325])^(a[142] & b[326])^(a[141] & b[327])^(a[140] & b[328])^(a[139] & b[329])^(a[138] & b[330])^(a[137] & b[331])^(a[136] & b[332])^(a[135] & b[333])^(a[134] & b[334])^(a[133] & b[335])^(a[132] & b[336])^(a[131] & b[337])^(a[130] & b[338])^(a[129] & b[339])^(a[128] & b[340])^(a[127] & b[341])^(a[126] & b[342])^(a[125] & b[343])^(a[124] & b[344])^(a[123] & b[345])^(a[122] & b[346])^(a[121] & b[347])^(a[120] & b[348])^(a[119] & b[349])^(a[118] & b[350])^(a[117] & b[351])^(a[116] & b[352])^(a[115] & b[353])^(a[114] & b[354])^(a[113] & b[355])^(a[112] & b[356])^(a[111] & b[357])^(a[110] & b[358])^(a[109] & b[359])^(a[108] & b[360])^(a[107] & b[361])^(a[106] & b[362])^(a[105] & b[363])^(a[104] & b[364])^(a[103] & b[365])^(a[102] & b[366])^(a[101] & b[367])^(a[100] & b[368])^(a[99] & b[369])^(a[98] & b[370])^(a[97] & b[371])^(a[96] & b[372])^(a[95] & b[373])^(a[94] & b[374])^(a[93] & b[375])^(a[92] & b[376])^(a[91] & b[377])^(a[90] & b[378])^(a[89] & b[379])^(a[88] & b[380])^(a[87] & b[381])^(a[86] & b[382])^(a[85] & b[383])^(a[84] & b[384])^(a[83] & b[385])^(a[82] & b[386])^(a[81] & b[387])^(a[80] & b[388])^(a[79] & b[389])^(a[78] & b[390])^(a[77] & b[391])^(a[76] & b[392])^(a[75] & b[393])^(a[74] & b[394])^(a[73] & b[395])^(a[72] & b[396])^(a[71] & b[397])^(a[70] & b[398])^(a[69] & b[399])^(a[68] & b[400])^(a[67] & b[401])^(a[66] & b[402])^(a[65] & b[403])^(a[64] & b[404])^(a[63] & b[405])^(a[62] & b[406])^(a[61] & b[407])^(a[60] & b[408]);
assign y[469] = (a[408] & b[61])^(a[407] & b[62])^(a[406] & b[63])^(a[405] & b[64])^(a[404] & b[65])^(a[403] & b[66])^(a[402] & b[67])^(a[401] & b[68])^(a[400] & b[69])^(a[399] & b[70])^(a[398] & b[71])^(a[397] & b[72])^(a[396] & b[73])^(a[395] & b[74])^(a[394] & b[75])^(a[393] & b[76])^(a[392] & b[77])^(a[391] & b[78])^(a[390] & b[79])^(a[389] & b[80])^(a[388] & b[81])^(a[387] & b[82])^(a[386] & b[83])^(a[385] & b[84])^(a[384] & b[85])^(a[383] & b[86])^(a[382] & b[87])^(a[381] & b[88])^(a[380] & b[89])^(a[379] & b[90])^(a[378] & b[91])^(a[377] & b[92])^(a[376] & b[93])^(a[375] & b[94])^(a[374] & b[95])^(a[373] & b[96])^(a[372] & b[97])^(a[371] & b[98])^(a[370] & b[99])^(a[369] & b[100])^(a[368] & b[101])^(a[367] & b[102])^(a[366] & b[103])^(a[365] & b[104])^(a[364] & b[105])^(a[363] & b[106])^(a[362] & b[107])^(a[361] & b[108])^(a[360] & b[109])^(a[359] & b[110])^(a[358] & b[111])^(a[357] & b[112])^(a[356] & b[113])^(a[355] & b[114])^(a[354] & b[115])^(a[353] & b[116])^(a[352] & b[117])^(a[351] & b[118])^(a[350] & b[119])^(a[349] & b[120])^(a[348] & b[121])^(a[347] & b[122])^(a[346] & b[123])^(a[345] & b[124])^(a[344] & b[125])^(a[343] & b[126])^(a[342] & b[127])^(a[341] & b[128])^(a[340] & b[129])^(a[339] & b[130])^(a[338] & b[131])^(a[337] & b[132])^(a[336] & b[133])^(a[335] & b[134])^(a[334] & b[135])^(a[333] & b[136])^(a[332] & b[137])^(a[331] & b[138])^(a[330] & b[139])^(a[329] & b[140])^(a[328] & b[141])^(a[327] & b[142])^(a[326] & b[143])^(a[325] & b[144])^(a[324] & b[145])^(a[323] & b[146])^(a[322] & b[147])^(a[321] & b[148])^(a[320] & b[149])^(a[319] & b[150])^(a[318] & b[151])^(a[317] & b[152])^(a[316] & b[153])^(a[315] & b[154])^(a[314] & b[155])^(a[313] & b[156])^(a[312] & b[157])^(a[311] & b[158])^(a[310] & b[159])^(a[309] & b[160])^(a[308] & b[161])^(a[307] & b[162])^(a[306] & b[163])^(a[305] & b[164])^(a[304] & b[165])^(a[303] & b[166])^(a[302] & b[167])^(a[301] & b[168])^(a[300] & b[169])^(a[299] & b[170])^(a[298] & b[171])^(a[297] & b[172])^(a[296] & b[173])^(a[295] & b[174])^(a[294] & b[175])^(a[293] & b[176])^(a[292] & b[177])^(a[291] & b[178])^(a[290] & b[179])^(a[289] & b[180])^(a[288] & b[181])^(a[287] & b[182])^(a[286] & b[183])^(a[285] & b[184])^(a[284] & b[185])^(a[283] & b[186])^(a[282] & b[187])^(a[281] & b[188])^(a[280] & b[189])^(a[279] & b[190])^(a[278] & b[191])^(a[277] & b[192])^(a[276] & b[193])^(a[275] & b[194])^(a[274] & b[195])^(a[273] & b[196])^(a[272] & b[197])^(a[271] & b[198])^(a[270] & b[199])^(a[269] & b[200])^(a[268] & b[201])^(a[267] & b[202])^(a[266] & b[203])^(a[265] & b[204])^(a[264] & b[205])^(a[263] & b[206])^(a[262] & b[207])^(a[261] & b[208])^(a[260] & b[209])^(a[259] & b[210])^(a[258] & b[211])^(a[257] & b[212])^(a[256] & b[213])^(a[255] & b[214])^(a[254] & b[215])^(a[253] & b[216])^(a[252] & b[217])^(a[251] & b[218])^(a[250] & b[219])^(a[249] & b[220])^(a[248] & b[221])^(a[247] & b[222])^(a[246] & b[223])^(a[245] & b[224])^(a[244] & b[225])^(a[243] & b[226])^(a[242] & b[227])^(a[241] & b[228])^(a[240] & b[229])^(a[239] & b[230])^(a[238] & b[231])^(a[237] & b[232])^(a[236] & b[233])^(a[235] & b[234])^(a[234] & b[235])^(a[233] & b[236])^(a[232] & b[237])^(a[231] & b[238])^(a[230] & b[239])^(a[229] & b[240])^(a[228] & b[241])^(a[227] & b[242])^(a[226] & b[243])^(a[225] & b[244])^(a[224] & b[245])^(a[223] & b[246])^(a[222] & b[247])^(a[221] & b[248])^(a[220] & b[249])^(a[219] & b[250])^(a[218] & b[251])^(a[217] & b[252])^(a[216] & b[253])^(a[215] & b[254])^(a[214] & b[255])^(a[213] & b[256])^(a[212] & b[257])^(a[211] & b[258])^(a[210] & b[259])^(a[209] & b[260])^(a[208] & b[261])^(a[207] & b[262])^(a[206] & b[263])^(a[205] & b[264])^(a[204] & b[265])^(a[203] & b[266])^(a[202] & b[267])^(a[201] & b[268])^(a[200] & b[269])^(a[199] & b[270])^(a[198] & b[271])^(a[197] & b[272])^(a[196] & b[273])^(a[195] & b[274])^(a[194] & b[275])^(a[193] & b[276])^(a[192] & b[277])^(a[191] & b[278])^(a[190] & b[279])^(a[189] & b[280])^(a[188] & b[281])^(a[187] & b[282])^(a[186] & b[283])^(a[185] & b[284])^(a[184] & b[285])^(a[183] & b[286])^(a[182] & b[287])^(a[181] & b[288])^(a[180] & b[289])^(a[179] & b[290])^(a[178] & b[291])^(a[177] & b[292])^(a[176] & b[293])^(a[175] & b[294])^(a[174] & b[295])^(a[173] & b[296])^(a[172] & b[297])^(a[171] & b[298])^(a[170] & b[299])^(a[169] & b[300])^(a[168] & b[301])^(a[167] & b[302])^(a[166] & b[303])^(a[165] & b[304])^(a[164] & b[305])^(a[163] & b[306])^(a[162] & b[307])^(a[161] & b[308])^(a[160] & b[309])^(a[159] & b[310])^(a[158] & b[311])^(a[157] & b[312])^(a[156] & b[313])^(a[155] & b[314])^(a[154] & b[315])^(a[153] & b[316])^(a[152] & b[317])^(a[151] & b[318])^(a[150] & b[319])^(a[149] & b[320])^(a[148] & b[321])^(a[147] & b[322])^(a[146] & b[323])^(a[145] & b[324])^(a[144] & b[325])^(a[143] & b[326])^(a[142] & b[327])^(a[141] & b[328])^(a[140] & b[329])^(a[139] & b[330])^(a[138] & b[331])^(a[137] & b[332])^(a[136] & b[333])^(a[135] & b[334])^(a[134] & b[335])^(a[133] & b[336])^(a[132] & b[337])^(a[131] & b[338])^(a[130] & b[339])^(a[129] & b[340])^(a[128] & b[341])^(a[127] & b[342])^(a[126] & b[343])^(a[125] & b[344])^(a[124] & b[345])^(a[123] & b[346])^(a[122] & b[347])^(a[121] & b[348])^(a[120] & b[349])^(a[119] & b[350])^(a[118] & b[351])^(a[117] & b[352])^(a[116] & b[353])^(a[115] & b[354])^(a[114] & b[355])^(a[113] & b[356])^(a[112] & b[357])^(a[111] & b[358])^(a[110] & b[359])^(a[109] & b[360])^(a[108] & b[361])^(a[107] & b[362])^(a[106] & b[363])^(a[105] & b[364])^(a[104] & b[365])^(a[103] & b[366])^(a[102] & b[367])^(a[101] & b[368])^(a[100] & b[369])^(a[99] & b[370])^(a[98] & b[371])^(a[97] & b[372])^(a[96] & b[373])^(a[95] & b[374])^(a[94] & b[375])^(a[93] & b[376])^(a[92] & b[377])^(a[91] & b[378])^(a[90] & b[379])^(a[89] & b[380])^(a[88] & b[381])^(a[87] & b[382])^(a[86] & b[383])^(a[85] & b[384])^(a[84] & b[385])^(a[83] & b[386])^(a[82] & b[387])^(a[81] & b[388])^(a[80] & b[389])^(a[79] & b[390])^(a[78] & b[391])^(a[77] & b[392])^(a[76] & b[393])^(a[75] & b[394])^(a[74] & b[395])^(a[73] & b[396])^(a[72] & b[397])^(a[71] & b[398])^(a[70] & b[399])^(a[69] & b[400])^(a[68] & b[401])^(a[67] & b[402])^(a[66] & b[403])^(a[65] & b[404])^(a[64] & b[405])^(a[63] & b[406])^(a[62] & b[407])^(a[61] & b[408]);
assign y[470] = (a[408] & b[62])^(a[407] & b[63])^(a[406] & b[64])^(a[405] & b[65])^(a[404] & b[66])^(a[403] & b[67])^(a[402] & b[68])^(a[401] & b[69])^(a[400] & b[70])^(a[399] & b[71])^(a[398] & b[72])^(a[397] & b[73])^(a[396] & b[74])^(a[395] & b[75])^(a[394] & b[76])^(a[393] & b[77])^(a[392] & b[78])^(a[391] & b[79])^(a[390] & b[80])^(a[389] & b[81])^(a[388] & b[82])^(a[387] & b[83])^(a[386] & b[84])^(a[385] & b[85])^(a[384] & b[86])^(a[383] & b[87])^(a[382] & b[88])^(a[381] & b[89])^(a[380] & b[90])^(a[379] & b[91])^(a[378] & b[92])^(a[377] & b[93])^(a[376] & b[94])^(a[375] & b[95])^(a[374] & b[96])^(a[373] & b[97])^(a[372] & b[98])^(a[371] & b[99])^(a[370] & b[100])^(a[369] & b[101])^(a[368] & b[102])^(a[367] & b[103])^(a[366] & b[104])^(a[365] & b[105])^(a[364] & b[106])^(a[363] & b[107])^(a[362] & b[108])^(a[361] & b[109])^(a[360] & b[110])^(a[359] & b[111])^(a[358] & b[112])^(a[357] & b[113])^(a[356] & b[114])^(a[355] & b[115])^(a[354] & b[116])^(a[353] & b[117])^(a[352] & b[118])^(a[351] & b[119])^(a[350] & b[120])^(a[349] & b[121])^(a[348] & b[122])^(a[347] & b[123])^(a[346] & b[124])^(a[345] & b[125])^(a[344] & b[126])^(a[343] & b[127])^(a[342] & b[128])^(a[341] & b[129])^(a[340] & b[130])^(a[339] & b[131])^(a[338] & b[132])^(a[337] & b[133])^(a[336] & b[134])^(a[335] & b[135])^(a[334] & b[136])^(a[333] & b[137])^(a[332] & b[138])^(a[331] & b[139])^(a[330] & b[140])^(a[329] & b[141])^(a[328] & b[142])^(a[327] & b[143])^(a[326] & b[144])^(a[325] & b[145])^(a[324] & b[146])^(a[323] & b[147])^(a[322] & b[148])^(a[321] & b[149])^(a[320] & b[150])^(a[319] & b[151])^(a[318] & b[152])^(a[317] & b[153])^(a[316] & b[154])^(a[315] & b[155])^(a[314] & b[156])^(a[313] & b[157])^(a[312] & b[158])^(a[311] & b[159])^(a[310] & b[160])^(a[309] & b[161])^(a[308] & b[162])^(a[307] & b[163])^(a[306] & b[164])^(a[305] & b[165])^(a[304] & b[166])^(a[303] & b[167])^(a[302] & b[168])^(a[301] & b[169])^(a[300] & b[170])^(a[299] & b[171])^(a[298] & b[172])^(a[297] & b[173])^(a[296] & b[174])^(a[295] & b[175])^(a[294] & b[176])^(a[293] & b[177])^(a[292] & b[178])^(a[291] & b[179])^(a[290] & b[180])^(a[289] & b[181])^(a[288] & b[182])^(a[287] & b[183])^(a[286] & b[184])^(a[285] & b[185])^(a[284] & b[186])^(a[283] & b[187])^(a[282] & b[188])^(a[281] & b[189])^(a[280] & b[190])^(a[279] & b[191])^(a[278] & b[192])^(a[277] & b[193])^(a[276] & b[194])^(a[275] & b[195])^(a[274] & b[196])^(a[273] & b[197])^(a[272] & b[198])^(a[271] & b[199])^(a[270] & b[200])^(a[269] & b[201])^(a[268] & b[202])^(a[267] & b[203])^(a[266] & b[204])^(a[265] & b[205])^(a[264] & b[206])^(a[263] & b[207])^(a[262] & b[208])^(a[261] & b[209])^(a[260] & b[210])^(a[259] & b[211])^(a[258] & b[212])^(a[257] & b[213])^(a[256] & b[214])^(a[255] & b[215])^(a[254] & b[216])^(a[253] & b[217])^(a[252] & b[218])^(a[251] & b[219])^(a[250] & b[220])^(a[249] & b[221])^(a[248] & b[222])^(a[247] & b[223])^(a[246] & b[224])^(a[245] & b[225])^(a[244] & b[226])^(a[243] & b[227])^(a[242] & b[228])^(a[241] & b[229])^(a[240] & b[230])^(a[239] & b[231])^(a[238] & b[232])^(a[237] & b[233])^(a[236] & b[234])^(a[235] & b[235])^(a[234] & b[236])^(a[233] & b[237])^(a[232] & b[238])^(a[231] & b[239])^(a[230] & b[240])^(a[229] & b[241])^(a[228] & b[242])^(a[227] & b[243])^(a[226] & b[244])^(a[225] & b[245])^(a[224] & b[246])^(a[223] & b[247])^(a[222] & b[248])^(a[221] & b[249])^(a[220] & b[250])^(a[219] & b[251])^(a[218] & b[252])^(a[217] & b[253])^(a[216] & b[254])^(a[215] & b[255])^(a[214] & b[256])^(a[213] & b[257])^(a[212] & b[258])^(a[211] & b[259])^(a[210] & b[260])^(a[209] & b[261])^(a[208] & b[262])^(a[207] & b[263])^(a[206] & b[264])^(a[205] & b[265])^(a[204] & b[266])^(a[203] & b[267])^(a[202] & b[268])^(a[201] & b[269])^(a[200] & b[270])^(a[199] & b[271])^(a[198] & b[272])^(a[197] & b[273])^(a[196] & b[274])^(a[195] & b[275])^(a[194] & b[276])^(a[193] & b[277])^(a[192] & b[278])^(a[191] & b[279])^(a[190] & b[280])^(a[189] & b[281])^(a[188] & b[282])^(a[187] & b[283])^(a[186] & b[284])^(a[185] & b[285])^(a[184] & b[286])^(a[183] & b[287])^(a[182] & b[288])^(a[181] & b[289])^(a[180] & b[290])^(a[179] & b[291])^(a[178] & b[292])^(a[177] & b[293])^(a[176] & b[294])^(a[175] & b[295])^(a[174] & b[296])^(a[173] & b[297])^(a[172] & b[298])^(a[171] & b[299])^(a[170] & b[300])^(a[169] & b[301])^(a[168] & b[302])^(a[167] & b[303])^(a[166] & b[304])^(a[165] & b[305])^(a[164] & b[306])^(a[163] & b[307])^(a[162] & b[308])^(a[161] & b[309])^(a[160] & b[310])^(a[159] & b[311])^(a[158] & b[312])^(a[157] & b[313])^(a[156] & b[314])^(a[155] & b[315])^(a[154] & b[316])^(a[153] & b[317])^(a[152] & b[318])^(a[151] & b[319])^(a[150] & b[320])^(a[149] & b[321])^(a[148] & b[322])^(a[147] & b[323])^(a[146] & b[324])^(a[145] & b[325])^(a[144] & b[326])^(a[143] & b[327])^(a[142] & b[328])^(a[141] & b[329])^(a[140] & b[330])^(a[139] & b[331])^(a[138] & b[332])^(a[137] & b[333])^(a[136] & b[334])^(a[135] & b[335])^(a[134] & b[336])^(a[133] & b[337])^(a[132] & b[338])^(a[131] & b[339])^(a[130] & b[340])^(a[129] & b[341])^(a[128] & b[342])^(a[127] & b[343])^(a[126] & b[344])^(a[125] & b[345])^(a[124] & b[346])^(a[123] & b[347])^(a[122] & b[348])^(a[121] & b[349])^(a[120] & b[350])^(a[119] & b[351])^(a[118] & b[352])^(a[117] & b[353])^(a[116] & b[354])^(a[115] & b[355])^(a[114] & b[356])^(a[113] & b[357])^(a[112] & b[358])^(a[111] & b[359])^(a[110] & b[360])^(a[109] & b[361])^(a[108] & b[362])^(a[107] & b[363])^(a[106] & b[364])^(a[105] & b[365])^(a[104] & b[366])^(a[103] & b[367])^(a[102] & b[368])^(a[101] & b[369])^(a[100] & b[370])^(a[99] & b[371])^(a[98] & b[372])^(a[97] & b[373])^(a[96] & b[374])^(a[95] & b[375])^(a[94] & b[376])^(a[93] & b[377])^(a[92] & b[378])^(a[91] & b[379])^(a[90] & b[380])^(a[89] & b[381])^(a[88] & b[382])^(a[87] & b[383])^(a[86] & b[384])^(a[85] & b[385])^(a[84] & b[386])^(a[83] & b[387])^(a[82] & b[388])^(a[81] & b[389])^(a[80] & b[390])^(a[79] & b[391])^(a[78] & b[392])^(a[77] & b[393])^(a[76] & b[394])^(a[75] & b[395])^(a[74] & b[396])^(a[73] & b[397])^(a[72] & b[398])^(a[71] & b[399])^(a[70] & b[400])^(a[69] & b[401])^(a[68] & b[402])^(a[67] & b[403])^(a[66] & b[404])^(a[65] & b[405])^(a[64] & b[406])^(a[63] & b[407])^(a[62] & b[408]);
assign y[471] = (a[408] & b[63])^(a[407] & b[64])^(a[406] & b[65])^(a[405] & b[66])^(a[404] & b[67])^(a[403] & b[68])^(a[402] & b[69])^(a[401] & b[70])^(a[400] & b[71])^(a[399] & b[72])^(a[398] & b[73])^(a[397] & b[74])^(a[396] & b[75])^(a[395] & b[76])^(a[394] & b[77])^(a[393] & b[78])^(a[392] & b[79])^(a[391] & b[80])^(a[390] & b[81])^(a[389] & b[82])^(a[388] & b[83])^(a[387] & b[84])^(a[386] & b[85])^(a[385] & b[86])^(a[384] & b[87])^(a[383] & b[88])^(a[382] & b[89])^(a[381] & b[90])^(a[380] & b[91])^(a[379] & b[92])^(a[378] & b[93])^(a[377] & b[94])^(a[376] & b[95])^(a[375] & b[96])^(a[374] & b[97])^(a[373] & b[98])^(a[372] & b[99])^(a[371] & b[100])^(a[370] & b[101])^(a[369] & b[102])^(a[368] & b[103])^(a[367] & b[104])^(a[366] & b[105])^(a[365] & b[106])^(a[364] & b[107])^(a[363] & b[108])^(a[362] & b[109])^(a[361] & b[110])^(a[360] & b[111])^(a[359] & b[112])^(a[358] & b[113])^(a[357] & b[114])^(a[356] & b[115])^(a[355] & b[116])^(a[354] & b[117])^(a[353] & b[118])^(a[352] & b[119])^(a[351] & b[120])^(a[350] & b[121])^(a[349] & b[122])^(a[348] & b[123])^(a[347] & b[124])^(a[346] & b[125])^(a[345] & b[126])^(a[344] & b[127])^(a[343] & b[128])^(a[342] & b[129])^(a[341] & b[130])^(a[340] & b[131])^(a[339] & b[132])^(a[338] & b[133])^(a[337] & b[134])^(a[336] & b[135])^(a[335] & b[136])^(a[334] & b[137])^(a[333] & b[138])^(a[332] & b[139])^(a[331] & b[140])^(a[330] & b[141])^(a[329] & b[142])^(a[328] & b[143])^(a[327] & b[144])^(a[326] & b[145])^(a[325] & b[146])^(a[324] & b[147])^(a[323] & b[148])^(a[322] & b[149])^(a[321] & b[150])^(a[320] & b[151])^(a[319] & b[152])^(a[318] & b[153])^(a[317] & b[154])^(a[316] & b[155])^(a[315] & b[156])^(a[314] & b[157])^(a[313] & b[158])^(a[312] & b[159])^(a[311] & b[160])^(a[310] & b[161])^(a[309] & b[162])^(a[308] & b[163])^(a[307] & b[164])^(a[306] & b[165])^(a[305] & b[166])^(a[304] & b[167])^(a[303] & b[168])^(a[302] & b[169])^(a[301] & b[170])^(a[300] & b[171])^(a[299] & b[172])^(a[298] & b[173])^(a[297] & b[174])^(a[296] & b[175])^(a[295] & b[176])^(a[294] & b[177])^(a[293] & b[178])^(a[292] & b[179])^(a[291] & b[180])^(a[290] & b[181])^(a[289] & b[182])^(a[288] & b[183])^(a[287] & b[184])^(a[286] & b[185])^(a[285] & b[186])^(a[284] & b[187])^(a[283] & b[188])^(a[282] & b[189])^(a[281] & b[190])^(a[280] & b[191])^(a[279] & b[192])^(a[278] & b[193])^(a[277] & b[194])^(a[276] & b[195])^(a[275] & b[196])^(a[274] & b[197])^(a[273] & b[198])^(a[272] & b[199])^(a[271] & b[200])^(a[270] & b[201])^(a[269] & b[202])^(a[268] & b[203])^(a[267] & b[204])^(a[266] & b[205])^(a[265] & b[206])^(a[264] & b[207])^(a[263] & b[208])^(a[262] & b[209])^(a[261] & b[210])^(a[260] & b[211])^(a[259] & b[212])^(a[258] & b[213])^(a[257] & b[214])^(a[256] & b[215])^(a[255] & b[216])^(a[254] & b[217])^(a[253] & b[218])^(a[252] & b[219])^(a[251] & b[220])^(a[250] & b[221])^(a[249] & b[222])^(a[248] & b[223])^(a[247] & b[224])^(a[246] & b[225])^(a[245] & b[226])^(a[244] & b[227])^(a[243] & b[228])^(a[242] & b[229])^(a[241] & b[230])^(a[240] & b[231])^(a[239] & b[232])^(a[238] & b[233])^(a[237] & b[234])^(a[236] & b[235])^(a[235] & b[236])^(a[234] & b[237])^(a[233] & b[238])^(a[232] & b[239])^(a[231] & b[240])^(a[230] & b[241])^(a[229] & b[242])^(a[228] & b[243])^(a[227] & b[244])^(a[226] & b[245])^(a[225] & b[246])^(a[224] & b[247])^(a[223] & b[248])^(a[222] & b[249])^(a[221] & b[250])^(a[220] & b[251])^(a[219] & b[252])^(a[218] & b[253])^(a[217] & b[254])^(a[216] & b[255])^(a[215] & b[256])^(a[214] & b[257])^(a[213] & b[258])^(a[212] & b[259])^(a[211] & b[260])^(a[210] & b[261])^(a[209] & b[262])^(a[208] & b[263])^(a[207] & b[264])^(a[206] & b[265])^(a[205] & b[266])^(a[204] & b[267])^(a[203] & b[268])^(a[202] & b[269])^(a[201] & b[270])^(a[200] & b[271])^(a[199] & b[272])^(a[198] & b[273])^(a[197] & b[274])^(a[196] & b[275])^(a[195] & b[276])^(a[194] & b[277])^(a[193] & b[278])^(a[192] & b[279])^(a[191] & b[280])^(a[190] & b[281])^(a[189] & b[282])^(a[188] & b[283])^(a[187] & b[284])^(a[186] & b[285])^(a[185] & b[286])^(a[184] & b[287])^(a[183] & b[288])^(a[182] & b[289])^(a[181] & b[290])^(a[180] & b[291])^(a[179] & b[292])^(a[178] & b[293])^(a[177] & b[294])^(a[176] & b[295])^(a[175] & b[296])^(a[174] & b[297])^(a[173] & b[298])^(a[172] & b[299])^(a[171] & b[300])^(a[170] & b[301])^(a[169] & b[302])^(a[168] & b[303])^(a[167] & b[304])^(a[166] & b[305])^(a[165] & b[306])^(a[164] & b[307])^(a[163] & b[308])^(a[162] & b[309])^(a[161] & b[310])^(a[160] & b[311])^(a[159] & b[312])^(a[158] & b[313])^(a[157] & b[314])^(a[156] & b[315])^(a[155] & b[316])^(a[154] & b[317])^(a[153] & b[318])^(a[152] & b[319])^(a[151] & b[320])^(a[150] & b[321])^(a[149] & b[322])^(a[148] & b[323])^(a[147] & b[324])^(a[146] & b[325])^(a[145] & b[326])^(a[144] & b[327])^(a[143] & b[328])^(a[142] & b[329])^(a[141] & b[330])^(a[140] & b[331])^(a[139] & b[332])^(a[138] & b[333])^(a[137] & b[334])^(a[136] & b[335])^(a[135] & b[336])^(a[134] & b[337])^(a[133] & b[338])^(a[132] & b[339])^(a[131] & b[340])^(a[130] & b[341])^(a[129] & b[342])^(a[128] & b[343])^(a[127] & b[344])^(a[126] & b[345])^(a[125] & b[346])^(a[124] & b[347])^(a[123] & b[348])^(a[122] & b[349])^(a[121] & b[350])^(a[120] & b[351])^(a[119] & b[352])^(a[118] & b[353])^(a[117] & b[354])^(a[116] & b[355])^(a[115] & b[356])^(a[114] & b[357])^(a[113] & b[358])^(a[112] & b[359])^(a[111] & b[360])^(a[110] & b[361])^(a[109] & b[362])^(a[108] & b[363])^(a[107] & b[364])^(a[106] & b[365])^(a[105] & b[366])^(a[104] & b[367])^(a[103] & b[368])^(a[102] & b[369])^(a[101] & b[370])^(a[100] & b[371])^(a[99] & b[372])^(a[98] & b[373])^(a[97] & b[374])^(a[96] & b[375])^(a[95] & b[376])^(a[94] & b[377])^(a[93] & b[378])^(a[92] & b[379])^(a[91] & b[380])^(a[90] & b[381])^(a[89] & b[382])^(a[88] & b[383])^(a[87] & b[384])^(a[86] & b[385])^(a[85] & b[386])^(a[84] & b[387])^(a[83] & b[388])^(a[82] & b[389])^(a[81] & b[390])^(a[80] & b[391])^(a[79] & b[392])^(a[78] & b[393])^(a[77] & b[394])^(a[76] & b[395])^(a[75] & b[396])^(a[74] & b[397])^(a[73] & b[398])^(a[72] & b[399])^(a[71] & b[400])^(a[70] & b[401])^(a[69] & b[402])^(a[68] & b[403])^(a[67] & b[404])^(a[66] & b[405])^(a[65] & b[406])^(a[64] & b[407])^(a[63] & b[408]);
assign y[472] = (a[408] & b[64])^(a[407] & b[65])^(a[406] & b[66])^(a[405] & b[67])^(a[404] & b[68])^(a[403] & b[69])^(a[402] & b[70])^(a[401] & b[71])^(a[400] & b[72])^(a[399] & b[73])^(a[398] & b[74])^(a[397] & b[75])^(a[396] & b[76])^(a[395] & b[77])^(a[394] & b[78])^(a[393] & b[79])^(a[392] & b[80])^(a[391] & b[81])^(a[390] & b[82])^(a[389] & b[83])^(a[388] & b[84])^(a[387] & b[85])^(a[386] & b[86])^(a[385] & b[87])^(a[384] & b[88])^(a[383] & b[89])^(a[382] & b[90])^(a[381] & b[91])^(a[380] & b[92])^(a[379] & b[93])^(a[378] & b[94])^(a[377] & b[95])^(a[376] & b[96])^(a[375] & b[97])^(a[374] & b[98])^(a[373] & b[99])^(a[372] & b[100])^(a[371] & b[101])^(a[370] & b[102])^(a[369] & b[103])^(a[368] & b[104])^(a[367] & b[105])^(a[366] & b[106])^(a[365] & b[107])^(a[364] & b[108])^(a[363] & b[109])^(a[362] & b[110])^(a[361] & b[111])^(a[360] & b[112])^(a[359] & b[113])^(a[358] & b[114])^(a[357] & b[115])^(a[356] & b[116])^(a[355] & b[117])^(a[354] & b[118])^(a[353] & b[119])^(a[352] & b[120])^(a[351] & b[121])^(a[350] & b[122])^(a[349] & b[123])^(a[348] & b[124])^(a[347] & b[125])^(a[346] & b[126])^(a[345] & b[127])^(a[344] & b[128])^(a[343] & b[129])^(a[342] & b[130])^(a[341] & b[131])^(a[340] & b[132])^(a[339] & b[133])^(a[338] & b[134])^(a[337] & b[135])^(a[336] & b[136])^(a[335] & b[137])^(a[334] & b[138])^(a[333] & b[139])^(a[332] & b[140])^(a[331] & b[141])^(a[330] & b[142])^(a[329] & b[143])^(a[328] & b[144])^(a[327] & b[145])^(a[326] & b[146])^(a[325] & b[147])^(a[324] & b[148])^(a[323] & b[149])^(a[322] & b[150])^(a[321] & b[151])^(a[320] & b[152])^(a[319] & b[153])^(a[318] & b[154])^(a[317] & b[155])^(a[316] & b[156])^(a[315] & b[157])^(a[314] & b[158])^(a[313] & b[159])^(a[312] & b[160])^(a[311] & b[161])^(a[310] & b[162])^(a[309] & b[163])^(a[308] & b[164])^(a[307] & b[165])^(a[306] & b[166])^(a[305] & b[167])^(a[304] & b[168])^(a[303] & b[169])^(a[302] & b[170])^(a[301] & b[171])^(a[300] & b[172])^(a[299] & b[173])^(a[298] & b[174])^(a[297] & b[175])^(a[296] & b[176])^(a[295] & b[177])^(a[294] & b[178])^(a[293] & b[179])^(a[292] & b[180])^(a[291] & b[181])^(a[290] & b[182])^(a[289] & b[183])^(a[288] & b[184])^(a[287] & b[185])^(a[286] & b[186])^(a[285] & b[187])^(a[284] & b[188])^(a[283] & b[189])^(a[282] & b[190])^(a[281] & b[191])^(a[280] & b[192])^(a[279] & b[193])^(a[278] & b[194])^(a[277] & b[195])^(a[276] & b[196])^(a[275] & b[197])^(a[274] & b[198])^(a[273] & b[199])^(a[272] & b[200])^(a[271] & b[201])^(a[270] & b[202])^(a[269] & b[203])^(a[268] & b[204])^(a[267] & b[205])^(a[266] & b[206])^(a[265] & b[207])^(a[264] & b[208])^(a[263] & b[209])^(a[262] & b[210])^(a[261] & b[211])^(a[260] & b[212])^(a[259] & b[213])^(a[258] & b[214])^(a[257] & b[215])^(a[256] & b[216])^(a[255] & b[217])^(a[254] & b[218])^(a[253] & b[219])^(a[252] & b[220])^(a[251] & b[221])^(a[250] & b[222])^(a[249] & b[223])^(a[248] & b[224])^(a[247] & b[225])^(a[246] & b[226])^(a[245] & b[227])^(a[244] & b[228])^(a[243] & b[229])^(a[242] & b[230])^(a[241] & b[231])^(a[240] & b[232])^(a[239] & b[233])^(a[238] & b[234])^(a[237] & b[235])^(a[236] & b[236])^(a[235] & b[237])^(a[234] & b[238])^(a[233] & b[239])^(a[232] & b[240])^(a[231] & b[241])^(a[230] & b[242])^(a[229] & b[243])^(a[228] & b[244])^(a[227] & b[245])^(a[226] & b[246])^(a[225] & b[247])^(a[224] & b[248])^(a[223] & b[249])^(a[222] & b[250])^(a[221] & b[251])^(a[220] & b[252])^(a[219] & b[253])^(a[218] & b[254])^(a[217] & b[255])^(a[216] & b[256])^(a[215] & b[257])^(a[214] & b[258])^(a[213] & b[259])^(a[212] & b[260])^(a[211] & b[261])^(a[210] & b[262])^(a[209] & b[263])^(a[208] & b[264])^(a[207] & b[265])^(a[206] & b[266])^(a[205] & b[267])^(a[204] & b[268])^(a[203] & b[269])^(a[202] & b[270])^(a[201] & b[271])^(a[200] & b[272])^(a[199] & b[273])^(a[198] & b[274])^(a[197] & b[275])^(a[196] & b[276])^(a[195] & b[277])^(a[194] & b[278])^(a[193] & b[279])^(a[192] & b[280])^(a[191] & b[281])^(a[190] & b[282])^(a[189] & b[283])^(a[188] & b[284])^(a[187] & b[285])^(a[186] & b[286])^(a[185] & b[287])^(a[184] & b[288])^(a[183] & b[289])^(a[182] & b[290])^(a[181] & b[291])^(a[180] & b[292])^(a[179] & b[293])^(a[178] & b[294])^(a[177] & b[295])^(a[176] & b[296])^(a[175] & b[297])^(a[174] & b[298])^(a[173] & b[299])^(a[172] & b[300])^(a[171] & b[301])^(a[170] & b[302])^(a[169] & b[303])^(a[168] & b[304])^(a[167] & b[305])^(a[166] & b[306])^(a[165] & b[307])^(a[164] & b[308])^(a[163] & b[309])^(a[162] & b[310])^(a[161] & b[311])^(a[160] & b[312])^(a[159] & b[313])^(a[158] & b[314])^(a[157] & b[315])^(a[156] & b[316])^(a[155] & b[317])^(a[154] & b[318])^(a[153] & b[319])^(a[152] & b[320])^(a[151] & b[321])^(a[150] & b[322])^(a[149] & b[323])^(a[148] & b[324])^(a[147] & b[325])^(a[146] & b[326])^(a[145] & b[327])^(a[144] & b[328])^(a[143] & b[329])^(a[142] & b[330])^(a[141] & b[331])^(a[140] & b[332])^(a[139] & b[333])^(a[138] & b[334])^(a[137] & b[335])^(a[136] & b[336])^(a[135] & b[337])^(a[134] & b[338])^(a[133] & b[339])^(a[132] & b[340])^(a[131] & b[341])^(a[130] & b[342])^(a[129] & b[343])^(a[128] & b[344])^(a[127] & b[345])^(a[126] & b[346])^(a[125] & b[347])^(a[124] & b[348])^(a[123] & b[349])^(a[122] & b[350])^(a[121] & b[351])^(a[120] & b[352])^(a[119] & b[353])^(a[118] & b[354])^(a[117] & b[355])^(a[116] & b[356])^(a[115] & b[357])^(a[114] & b[358])^(a[113] & b[359])^(a[112] & b[360])^(a[111] & b[361])^(a[110] & b[362])^(a[109] & b[363])^(a[108] & b[364])^(a[107] & b[365])^(a[106] & b[366])^(a[105] & b[367])^(a[104] & b[368])^(a[103] & b[369])^(a[102] & b[370])^(a[101] & b[371])^(a[100] & b[372])^(a[99] & b[373])^(a[98] & b[374])^(a[97] & b[375])^(a[96] & b[376])^(a[95] & b[377])^(a[94] & b[378])^(a[93] & b[379])^(a[92] & b[380])^(a[91] & b[381])^(a[90] & b[382])^(a[89] & b[383])^(a[88] & b[384])^(a[87] & b[385])^(a[86] & b[386])^(a[85] & b[387])^(a[84] & b[388])^(a[83] & b[389])^(a[82] & b[390])^(a[81] & b[391])^(a[80] & b[392])^(a[79] & b[393])^(a[78] & b[394])^(a[77] & b[395])^(a[76] & b[396])^(a[75] & b[397])^(a[74] & b[398])^(a[73] & b[399])^(a[72] & b[400])^(a[71] & b[401])^(a[70] & b[402])^(a[69] & b[403])^(a[68] & b[404])^(a[67] & b[405])^(a[66] & b[406])^(a[65] & b[407])^(a[64] & b[408]);
assign y[473] = (a[408] & b[65])^(a[407] & b[66])^(a[406] & b[67])^(a[405] & b[68])^(a[404] & b[69])^(a[403] & b[70])^(a[402] & b[71])^(a[401] & b[72])^(a[400] & b[73])^(a[399] & b[74])^(a[398] & b[75])^(a[397] & b[76])^(a[396] & b[77])^(a[395] & b[78])^(a[394] & b[79])^(a[393] & b[80])^(a[392] & b[81])^(a[391] & b[82])^(a[390] & b[83])^(a[389] & b[84])^(a[388] & b[85])^(a[387] & b[86])^(a[386] & b[87])^(a[385] & b[88])^(a[384] & b[89])^(a[383] & b[90])^(a[382] & b[91])^(a[381] & b[92])^(a[380] & b[93])^(a[379] & b[94])^(a[378] & b[95])^(a[377] & b[96])^(a[376] & b[97])^(a[375] & b[98])^(a[374] & b[99])^(a[373] & b[100])^(a[372] & b[101])^(a[371] & b[102])^(a[370] & b[103])^(a[369] & b[104])^(a[368] & b[105])^(a[367] & b[106])^(a[366] & b[107])^(a[365] & b[108])^(a[364] & b[109])^(a[363] & b[110])^(a[362] & b[111])^(a[361] & b[112])^(a[360] & b[113])^(a[359] & b[114])^(a[358] & b[115])^(a[357] & b[116])^(a[356] & b[117])^(a[355] & b[118])^(a[354] & b[119])^(a[353] & b[120])^(a[352] & b[121])^(a[351] & b[122])^(a[350] & b[123])^(a[349] & b[124])^(a[348] & b[125])^(a[347] & b[126])^(a[346] & b[127])^(a[345] & b[128])^(a[344] & b[129])^(a[343] & b[130])^(a[342] & b[131])^(a[341] & b[132])^(a[340] & b[133])^(a[339] & b[134])^(a[338] & b[135])^(a[337] & b[136])^(a[336] & b[137])^(a[335] & b[138])^(a[334] & b[139])^(a[333] & b[140])^(a[332] & b[141])^(a[331] & b[142])^(a[330] & b[143])^(a[329] & b[144])^(a[328] & b[145])^(a[327] & b[146])^(a[326] & b[147])^(a[325] & b[148])^(a[324] & b[149])^(a[323] & b[150])^(a[322] & b[151])^(a[321] & b[152])^(a[320] & b[153])^(a[319] & b[154])^(a[318] & b[155])^(a[317] & b[156])^(a[316] & b[157])^(a[315] & b[158])^(a[314] & b[159])^(a[313] & b[160])^(a[312] & b[161])^(a[311] & b[162])^(a[310] & b[163])^(a[309] & b[164])^(a[308] & b[165])^(a[307] & b[166])^(a[306] & b[167])^(a[305] & b[168])^(a[304] & b[169])^(a[303] & b[170])^(a[302] & b[171])^(a[301] & b[172])^(a[300] & b[173])^(a[299] & b[174])^(a[298] & b[175])^(a[297] & b[176])^(a[296] & b[177])^(a[295] & b[178])^(a[294] & b[179])^(a[293] & b[180])^(a[292] & b[181])^(a[291] & b[182])^(a[290] & b[183])^(a[289] & b[184])^(a[288] & b[185])^(a[287] & b[186])^(a[286] & b[187])^(a[285] & b[188])^(a[284] & b[189])^(a[283] & b[190])^(a[282] & b[191])^(a[281] & b[192])^(a[280] & b[193])^(a[279] & b[194])^(a[278] & b[195])^(a[277] & b[196])^(a[276] & b[197])^(a[275] & b[198])^(a[274] & b[199])^(a[273] & b[200])^(a[272] & b[201])^(a[271] & b[202])^(a[270] & b[203])^(a[269] & b[204])^(a[268] & b[205])^(a[267] & b[206])^(a[266] & b[207])^(a[265] & b[208])^(a[264] & b[209])^(a[263] & b[210])^(a[262] & b[211])^(a[261] & b[212])^(a[260] & b[213])^(a[259] & b[214])^(a[258] & b[215])^(a[257] & b[216])^(a[256] & b[217])^(a[255] & b[218])^(a[254] & b[219])^(a[253] & b[220])^(a[252] & b[221])^(a[251] & b[222])^(a[250] & b[223])^(a[249] & b[224])^(a[248] & b[225])^(a[247] & b[226])^(a[246] & b[227])^(a[245] & b[228])^(a[244] & b[229])^(a[243] & b[230])^(a[242] & b[231])^(a[241] & b[232])^(a[240] & b[233])^(a[239] & b[234])^(a[238] & b[235])^(a[237] & b[236])^(a[236] & b[237])^(a[235] & b[238])^(a[234] & b[239])^(a[233] & b[240])^(a[232] & b[241])^(a[231] & b[242])^(a[230] & b[243])^(a[229] & b[244])^(a[228] & b[245])^(a[227] & b[246])^(a[226] & b[247])^(a[225] & b[248])^(a[224] & b[249])^(a[223] & b[250])^(a[222] & b[251])^(a[221] & b[252])^(a[220] & b[253])^(a[219] & b[254])^(a[218] & b[255])^(a[217] & b[256])^(a[216] & b[257])^(a[215] & b[258])^(a[214] & b[259])^(a[213] & b[260])^(a[212] & b[261])^(a[211] & b[262])^(a[210] & b[263])^(a[209] & b[264])^(a[208] & b[265])^(a[207] & b[266])^(a[206] & b[267])^(a[205] & b[268])^(a[204] & b[269])^(a[203] & b[270])^(a[202] & b[271])^(a[201] & b[272])^(a[200] & b[273])^(a[199] & b[274])^(a[198] & b[275])^(a[197] & b[276])^(a[196] & b[277])^(a[195] & b[278])^(a[194] & b[279])^(a[193] & b[280])^(a[192] & b[281])^(a[191] & b[282])^(a[190] & b[283])^(a[189] & b[284])^(a[188] & b[285])^(a[187] & b[286])^(a[186] & b[287])^(a[185] & b[288])^(a[184] & b[289])^(a[183] & b[290])^(a[182] & b[291])^(a[181] & b[292])^(a[180] & b[293])^(a[179] & b[294])^(a[178] & b[295])^(a[177] & b[296])^(a[176] & b[297])^(a[175] & b[298])^(a[174] & b[299])^(a[173] & b[300])^(a[172] & b[301])^(a[171] & b[302])^(a[170] & b[303])^(a[169] & b[304])^(a[168] & b[305])^(a[167] & b[306])^(a[166] & b[307])^(a[165] & b[308])^(a[164] & b[309])^(a[163] & b[310])^(a[162] & b[311])^(a[161] & b[312])^(a[160] & b[313])^(a[159] & b[314])^(a[158] & b[315])^(a[157] & b[316])^(a[156] & b[317])^(a[155] & b[318])^(a[154] & b[319])^(a[153] & b[320])^(a[152] & b[321])^(a[151] & b[322])^(a[150] & b[323])^(a[149] & b[324])^(a[148] & b[325])^(a[147] & b[326])^(a[146] & b[327])^(a[145] & b[328])^(a[144] & b[329])^(a[143] & b[330])^(a[142] & b[331])^(a[141] & b[332])^(a[140] & b[333])^(a[139] & b[334])^(a[138] & b[335])^(a[137] & b[336])^(a[136] & b[337])^(a[135] & b[338])^(a[134] & b[339])^(a[133] & b[340])^(a[132] & b[341])^(a[131] & b[342])^(a[130] & b[343])^(a[129] & b[344])^(a[128] & b[345])^(a[127] & b[346])^(a[126] & b[347])^(a[125] & b[348])^(a[124] & b[349])^(a[123] & b[350])^(a[122] & b[351])^(a[121] & b[352])^(a[120] & b[353])^(a[119] & b[354])^(a[118] & b[355])^(a[117] & b[356])^(a[116] & b[357])^(a[115] & b[358])^(a[114] & b[359])^(a[113] & b[360])^(a[112] & b[361])^(a[111] & b[362])^(a[110] & b[363])^(a[109] & b[364])^(a[108] & b[365])^(a[107] & b[366])^(a[106] & b[367])^(a[105] & b[368])^(a[104] & b[369])^(a[103] & b[370])^(a[102] & b[371])^(a[101] & b[372])^(a[100] & b[373])^(a[99] & b[374])^(a[98] & b[375])^(a[97] & b[376])^(a[96] & b[377])^(a[95] & b[378])^(a[94] & b[379])^(a[93] & b[380])^(a[92] & b[381])^(a[91] & b[382])^(a[90] & b[383])^(a[89] & b[384])^(a[88] & b[385])^(a[87] & b[386])^(a[86] & b[387])^(a[85] & b[388])^(a[84] & b[389])^(a[83] & b[390])^(a[82] & b[391])^(a[81] & b[392])^(a[80] & b[393])^(a[79] & b[394])^(a[78] & b[395])^(a[77] & b[396])^(a[76] & b[397])^(a[75] & b[398])^(a[74] & b[399])^(a[73] & b[400])^(a[72] & b[401])^(a[71] & b[402])^(a[70] & b[403])^(a[69] & b[404])^(a[68] & b[405])^(a[67] & b[406])^(a[66] & b[407])^(a[65] & b[408]);
assign y[474] = (a[408] & b[66])^(a[407] & b[67])^(a[406] & b[68])^(a[405] & b[69])^(a[404] & b[70])^(a[403] & b[71])^(a[402] & b[72])^(a[401] & b[73])^(a[400] & b[74])^(a[399] & b[75])^(a[398] & b[76])^(a[397] & b[77])^(a[396] & b[78])^(a[395] & b[79])^(a[394] & b[80])^(a[393] & b[81])^(a[392] & b[82])^(a[391] & b[83])^(a[390] & b[84])^(a[389] & b[85])^(a[388] & b[86])^(a[387] & b[87])^(a[386] & b[88])^(a[385] & b[89])^(a[384] & b[90])^(a[383] & b[91])^(a[382] & b[92])^(a[381] & b[93])^(a[380] & b[94])^(a[379] & b[95])^(a[378] & b[96])^(a[377] & b[97])^(a[376] & b[98])^(a[375] & b[99])^(a[374] & b[100])^(a[373] & b[101])^(a[372] & b[102])^(a[371] & b[103])^(a[370] & b[104])^(a[369] & b[105])^(a[368] & b[106])^(a[367] & b[107])^(a[366] & b[108])^(a[365] & b[109])^(a[364] & b[110])^(a[363] & b[111])^(a[362] & b[112])^(a[361] & b[113])^(a[360] & b[114])^(a[359] & b[115])^(a[358] & b[116])^(a[357] & b[117])^(a[356] & b[118])^(a[355] & b[119])^(a[354] & b[120])^(a[353] & b[121])^(a[352] & b[122])^(a[351] & b[123])^(a[350] & b[124])^(a[349] & b[125])^(a[348] & b[126])^(a[347] & b[127])^(a[346] & b[128])^(a[345] & b[129])^(a[344] & b[130])^(a[343] & b[131])^(a[342] & b[132])^(a[341] & b[133])^(a[340] & b[134])^(a[339] & b[135])^(a[338] & b[136])^(a[337] & b[137])^(a[336] & b[138])^(a[335] & b[139])^(a[334] & b[140])^(a[333] & b[141])^(a[332] & b[142])^(a[331] & b[143])^(a[330] & b[144])^(a[329] & b[145])^(a[328] & b[146])^(a[327] & b[147])^(a[326] & b[148])^(a[325] & b[149])^(a[324] & b[150])^(a[323] & b[151])^(a[322] & b[152])^(a[321] & b[153])^(a[320] & b[154])^(a[319] & b[155])^(a[318] & b[156])^(a[317] & b[157])^(a[316] & b[158])^(a[315] & b[159])^(a[314] & b[160])^(a[313] & b[161])^(a[312] & b[162])^(a[311] & b[163])^(a[310] & b[164])^(a[309] & b[165])^(a[308] & b[166])^(a[307] & b[167])^(a[306] & b[168])^(a[305] & b[169])^(a[304] & b[170])^(a[303] & b[171])^(a[302] & b[172])^(a[301] & b[173])^(a[300] & b[174])^(a[299] & b[175])^(a[298] & b[176])^(a[297] & b[177])^(a[296] & b[178])^(a[295] & b[179])^(a[294] & b[180])^(a[293] & b[181])^(a[292] & b[182])^(a[291] & b[183])^(a[290] & b[184])^(a[289] & b[185])^(a[288] & b[186])^(a[287] & b[187])^(a[286] & b[188])^(a[285] & b[189])^(a[284] & b[190])^(a[283] & b[191])^(a[282] & b[192])^(a[281] & b[193])^(a[280] & b[194])^(a[279] & b[195])^(a[278] & b[196])^(a[277] & b[197])^(a[276] & b[198])^(a[275] & b[199])^(a[274] & b[200])^(a[273] & b[201])^(a[272] & b[202])^(a[271] & b[203])^(a[270] & b[204])^(a[269] & b[205])^(a[268] & b[206])^(a[267] & b[207])^(a[266] & b[208])^(a[265] & b[209])^(a[264] & b[210])^(a[263] & b[211])^(a[262] & b[212])^(a[261] & b[213])^(a[260] & b[214])^(a[259] & b[215])^(a[258] & b[216])^(a[257] & b[217])^(a[256] & b[218])^(a[255] & b[219])^(a[254] & b[220])^(a[253] & b[221])^(a[252] & b[222])^(a[251] & b[223])^(a[250] & b[224])^(a[249] & b[225])^(a[248] & b[226])^(a[247] & b[227])^(a[246] & b[228])^(a[245] & b[229])^(a[244] & b[230])^(a[243] & b[231])^(a[242] & b[232])^(a[241] & b[233])^(a[240] & b[234])^(a[239] & b[235])^(a[238] & b[236])^(a[237] & b[237])^(a[236] & b[238])^(a[235] & b[239])^(a[234] & b[240])^(a[233] & b[241])^(a[232] & b[242])^(a[231] & b[243])^(a[230] & b[244])^(a[229] & b[245])^(a[228] & b[246])^(a[227] & b[247])^(a[226] & b[248])^(a[225] & b[249])^(a[224] & b[250])^(a[223] & b[251])^(a[222] & b[252])^(a[221] & b[253])^(a[220] & b[254])^(a[219] & b[255])^(a[218] & b[256])^(a[217] & b[257])^(a[216] & b[258])^(a[215] & b[259])^(a[214] & b[260])^(a[213] & b[261])^(a[212] & b[262])^(a[211] & b[263])^(a[210] & b[264])^(a[209] & b[265])^(a[208] & b[266])^(a[207] & b[267])^(a[206] & b[268])^(a[205] & b[269])^(a[204] & b[270])^(a[203] & b[271])^(a[202] & b[272])^(a[201] & b[273])^(a[200] & b[274])^(a[199] & b[275])^(a[198] & b[276])^(a[197] & b[277])^(a[196] & b[278])^(a[195] & b[279])^(a[194] & b[280])^(a[193] & b[281])^(a[192] & b[282])^(a[191] & b[283])^(a[190] & b[284])^(a[189] & b[285])^(a[188] & b[286])^(a[187] & b[287])^(a[186] & b[288])^(a[185] & b[289])^(a[184] & b[290])^(a[183] & b[291])^(a[182] & b[292])^(a[181] & b[293])^(a[180] & b[294])^(a[179] & b[295])^(a[178] & b[296])^(a[177] & b[297])^(a[176] & b[298])^(a[175] & b[299])^(a[174] & b[300])^(a[173] & b[301])^(a[172] & b[302])^(a[171] & b[303])^(a[170] & b[304])^(a[169] & b[305])^(a[168] & b[306])^(a[167] & b[307])^(a[166] & b[308])^(a[165] & b[309])^(a[164] & b[310])^(a[163] & b[311])^(a[162] & b[312])^(a[161] & b[313])^(a[160] & b[314])^(a[159] & b[315])^(a[158] & b[316])^(a[157] & b[317])^(a[156] & b[318])^(a[155] & b[319])^(a[154] & b[320])^(a[153] & b[321])^(a[152] & b[322])^(a[151] & b[323])^(a[150] & b[324])^(a[149] & b[325])^(a[148] & b[326])^(a[147] & b[327])^(a[146] & b[328])^(a[145] & b[329])^(a[144] & b[330])^(a[143] & b[331])^(a[142] & b[332])^(a[141] & b[333])^(a[140] & b[334])^(a[139] & b[335])^(a[138] & b[336])^(a[137] & b[337])^(a[136] & b[338])^(a[135] & b[339])^(a[134] & b[340])^(a[133] & b[341])^(a[132] & b[342])^(a[131] & b[343])^(a[130] & b[344])^(a[129] & b[345])^(a[128] & b[346])^(a[127] & b[347])^(a[126] & b[348])^(a[125] & b[349])^(a[124] & b[350])^(a[123] & b[351])^(a[122] & b[352])^(a[121] & b[353])^(a[120] & b[354])^(a[119] & b[355])^(a[118] & b[356])^(a[117] & b[357])^(a[116] & b[358])^(a[115] & b[359])^(a[114] & b[360])^(a[113] & b[361])^(a[112] & b[362])^(a[111] & b[363])^(a[110] & b[364])^(a[109] & b[365])^(a[108] & b[366])^(a[107] & b[367])^(a[106] & b[368])^(a[105] & b[369])^(a[104] & b[370])^(a[103] & b[371])^(a[102] & b[372])^(a[101] & b[373])^(a[100] & b[374])^(a[99] & b[375])^(a[98] & b[376])^(a[97] & b[377])^(a[96] & b[378])^(a[95] & b[379])^(a[94] & b[380])^(a[93] & b[381])^(a[92] & b[382])^(a[91] & b[383])^(a[90] & b[384])^(a[89] & b[385])^(a[88] & b[386])^(a[87] & b[387])^(a[86] & b[388])^(a[85] & b[389])^(a[84] & b[390])^(a[83] & b[391])^(a[82] & b[392])^(a[81] & b[393])^(a[80] & b[394])^(a[79] & b[395])^(a[78] & b[396])^(a[77] & b[397])^(a[76] & b[398])^(a[75] & b[399])^(a[74] & b[400])^(a[73] & b[401])^(a[72] & b[402])^(a[71] & b[403])^(a[70] & b[404])^(a[69] & b[405])^(a[68] & b[406])^(a[67] & b[407])^(a[66] & b[408]);
assign y[475] = (a[408] & b[67])^(a[407] & b[68])^(a[406] & b[69])^(a[405] & b[70])^(a[404] & b[71])^(a[403] & b[72])^(a[402] & b[73])^(a[401] & b[74])^(a[400] & b[75])^(a[399] & b[76])^(a[398] & b[77])^(a[397] & b[78])^(a[396] & b[79])^(a[395] & b[80])^(a[394] & b[81])^(a[393] & b[82])^(a[392] & b[83])^(a[391] & b[84])^(a[390] & b[85])^(a[389] & b[86])^(a[388] & b[87])^(a[387] & b[88])^(a[386] & b[89])^(a[385] & b[90])^(a[384] & b[91])^(a[383] & b[92])^(a[382] & b[93])^(a[381] & b[94])^(a[380] & b[95])^(a[379] & b[96])^(a[378] & b[97])^(a[377] & b[98])^(a[376] & b[99])^(a[375] & b[100])^(a[374] & b[101])^(a[373] & b[102])^(a[372] & b[103])^(a[371] & b[104])^(a[370] & b[105])^(a[369] & b[106])^(a[368] & b[107])^(a[367] & b[108])^(a[366] & b[109])^(a[365] & b[110])^(a[364] & b[111])^(a[363] & b[112])^(a[362] & b[113])^(a[361] & b[114])^(a[360] & b[115])^(a[359] & b[116])^(a[358] & b[117])^(a[357] & b[118])^(a[356] & b[119])^(a[355] & b[120])^(a[354] & b[121])^(a[353] & b[122])^(a[352] & b[123])^(a[351] & b[124])^(a[350] & b[125])^(a[349] & b[126])^(a[348] & b[127])^(a[347] & b[128])^(a[346] & b[129])^(a[345] & b[130])^(a[344] & b[131])^(a[343] & b[132])^(a[342] & b[133])^(a[341] & b[134])^(a[340] & b[135])^(a[339] & b[136])^(a[338] & b[137])^(a[337] & b[138])^(a[336] & b[139])^(a[335] & b[140])^(a[334] & b[141])^(a[333] & b[142])^(a[332] & b[143])^(a[331] & b[144])^(a[330] & b[145])^(a[329] & b[146])^(a[328] & b[147])^(a[327] & b[148])^(a[326] & b[149])^(a[325] & b[150])^(a[324] & b[151])^(a[323] & b[152])^(a[322] & b[153])^(a[321] & b[154])^(a[320] & b[155])^(a[319] & b[156])^(a[318] & b[157])^(a[317] & b[158])^(a[316] & b[159])^(a[315] & b[160])^(a[314] & b[161])^(a[313] & b[162])^(a[312] & b[163])^(a[311] & b[164])^(a[310] & b[165])^(a[309] & b[166])^(a[308] & b[167])^(a[307] & b[168])^(a[306] & b[169])^(a[305] & b[170])^(a[304] & b[171])^(a[303] & b[172])^(a[302] & b[173])^(a[301] & b[174])^(a[300] & b[175])^(a[299] & b[176])^(a[298] & b[177])^(a[297] & b[178])^(a[296] & b[179])^(a[295] & b[180])^(a[294] & b[181])^(a[293] & b[182])^(a[292] & b[183])^(a[291] & b[184])^(a[290] & b[185])^(a[289] & b[186])^(a[288] & b[187])^(a[287] & b[188])^(a[286] & b[189])^(a[285] & b[190])^(a[284] & b[191])^(a[283] & b[192])^(a[282] & b[193])^(a[281] & b[194])^(a[280] & b[195])^(a[279] & b[196])^(a[278] & b[197])^(a[277] & b[198])^(a[276] & b[199])^(a[275] & b[200])^(a[274] & b[201])^(a[273] & b[202])^(a[272] & b[203])^(a[271] & b[204])^(a[270] & b[205])^(a[269] & b[206])^(a[268] & b[207])^(a[267] & b[208])^(a[266] & b[209])^(a[265] & b[210])^(a[264] & b[211])^(a[263] & b[212])^(a[262] & b[213])^(a[261] & b[214])^(a[260] & b[215])^(a[259] & b[216])^(a[258] & b[217])^(a[257] & b[218])^(a[256] & b[219])^(a[255] & b[220])^(a[254] & b[221])^(a[253] & b[222])^(a[252] & b[223])^(a[251] & b[224])^(a[250] & b[225])^(a[249] & b[226])^(a[248] & b[227])^(a[247] & b[228])^(a[246] & b[229])^(a[245] & b[230])^(a[244] & b[231])^(a[243] & b[232])^(a[242] & b[233])^(a[241] & b[234])^(a[240] & b[235])^(a[239] & b[236])^(a[238] & b[237])^(a[237] & b[238])^(a[236] & b[239])^(a[235] & b[240])^(a[234] & b[241])^(a[233] & b[242])^(a[232] & b[243])^(a[231] & b[244])^(a[230] & b[245])^(a[229] & b[246])^(a[228] & b[247])^(a[227] & b[248])^(a[226] & b[249])^(a[225] & b[250])^(a[224] & b[251])^(a[223] & b[252])^(a[222] & b[253])^(a[221] & b[254])^(a[220] & b[255])^(a[219] & b[256])^(a[218] & b[257])^(a[217] & b[258])^(a[216] & b[259])^(a[215] & b[260])^(a[214] & b[261])^(a[213] & b[262])^(a[212] & b[263])^(a[211] & b[264])^(a[210] & b[265])^(a[209] & b[266])^(a[208] & b[267])^(a[207] & b[268])^(a[206] & b[269])^(a[205] & b[270])^(a[204] & b[271])^(a[203] & b[272])^(a[202] & b[273])^(a[201] & b[274])^(a[200] & b[275])^(a[199] & b[276])^(a[198] & b[277])^(a[197] & b[278])^(a[196] & b[279])^(a[195] & b[280])^(a[194] & b[281])^(a[193] & b[282])^(a[192] & b[283])^(a[191] & b[284])^(a[190] & b[285])^(a[189] & b[286])^(a[188] & b[287])^(a[187] & b[288])^(a[186] & b[289])^(a[185] & b[290])^(a[184] & b[291])^(a[183] & b[292])^(a[182] & b[293])^(a[181] & b[294])^(a[180] & b[295])^(a[179] & b[296])^(a[178] & b[297])^(a[177] & b[298])^(a[176] & b[299])^(a[175] & b[300])^(a[174] & b[301])^(a[173] & b[302])^(a[172] & b[303])^(a[171] & b[304])^(a[170] & b[305])^(a[169] & b[306])^(a[168] & b[307])^(a[167] & b[308])^(a[166] & b[309])^(a[165] & b[310])^(a[164] & b[311])^(a[163] & b[312])^(a[162] & b[313])^(a[161] & b[314])^(a[160] & b[315])^(a[159] & b[316])^(a[158] & b[317])^(a[157] & b[318])^(a[156] & b[319])^(a[155] & b[320])^(a[154] & b[321])^(a[153] & b[322])^(a[152] & b[323])^(a[151] & b[324])^(a[150] & b[325])^(a[149] & b[326])^(a[148] & b[327])^(a[147] & b[328])^(a[146] & b[329])^(a[145] & b[330])^(a[144] & b[331])^(a[143] & b[332])^(a[142] & b[333])^(a[141] & b[334])^(a[140] & b[335])^(a[139] & b[336])^(a[138] & b[337])^(a[137] & b[338])^(a[136] & b[339])^(a[135] & b[340])^(a[134] & b[341])^(a[133] & b[342])^(a[132] & b[343])^(a[131] & b[344])^(a[130] & b[345])^(a[129] & b[346])^(a[128] & b[347])^(a[127] & b[348])^(a[126] & b[349])^(a[125] & b[350])^(a[124] & b[351])^(a[123] & b[352])^(a[122] & b[353])^(a[121] & b[354])^(a[120] & b[355])^(a[119] & b[356])^(a[118] & b[357])^(a[117] & b[358])^(a[116] & b[359])^(a[115] & b[360])^(a[114] & b[361])^(a[113] & b[362])^(a[112] & b[363])^(a[111] & b[364])^(a[110] & b[365])^(a[109] & b[366])^(a[108] & b[367])^(a[107] & b[368])^(a[106] & b[369])^(a[105] & b[370])^(a[104] & b[371])^(a[103] & b[372])^(a[102] & b[373])^(a[101] & b[374])^(a[100] & b[375])^(a[99] & b[376])^(a[98] & b[377])^(a[97] & b[378])^(a[96] & b[379])^(a[95] & b[380])^(a[94] & b[381])^(a[93] & b[382])^(a[92] & b[383])^(a[91] & b[384])^(a[90] & b[385])^(a[89] & b[386])^(a[88] & b[387])^(a[87] & b[388])^(a[86] & b[389])^(a[85] & b[390])^(a[84] & b[391])^(a[83] & b[392])^(a[82] & b[393])^(a[81] & b[394])^(a[80] & b[395])^(a[79] & b[396])^(a[78] & b[397])^(a[77] & b[398])^(a[76] & b[399])^(a[75] & b[400])^(a[74] & b[401])^(a[73] & b[402])^(a[72] & b[403])^(a[71] & b[404])^(a[70] & b[405])^(a[69] & b[406])^(a[68] & b[407])^(a[67] & b[408]);
assign y[476] = (a[408] & b[68])^(a[407] & b[69])^(a[406] & b[70])^(a[405] & b[71])^(a[404] & b[72])^(a[403] & b[73])^(a[402] & b[74])^(a[401] & b[75])^(a[400] & b[76])^(a[399] & b[77])^(a[398] & b[78])^(a[397] & b[79])^(a[396] & b[80])^(a[395] & b[81])^(a[394] & b[82])^(a[393] & b[83])^(a[392] & b[84])^(a[391] & b[85])^(a[390] & b[86])^(a[389] & b[87])^(a[388] & b[88])^(a[387] & b[89])^(a[386] & b[90])^(a[385] & b[91])^(a[384] & b[92])^(a[383] & b[93])^(a[382] & b[94])^(a[381] & b[95])^(a[380] & b[96])^(a[379] & b[97])^(a[378] & b[98])^(a[377] & b[99])^(a[376] & b[100])^(a[375] & b[101])^(a[374] & b[102])^(a[373] & b[103])^(a[372] & b[104])^(a[371] & b[105])^(a[370] & b[106])^(a[369] & b[107])^(a[368] & b[108])^(a[367] & b[109])^(a[366] & b[110])^(a[365] & b[111])^(a[364] & b[112])^(a[363] & b[113])^(a[362] & b[114])^(a[361] & b[115])^(a[360] & b[116])^(a[359] & b[117])^(a[358] & b[118])^(a[357] & b[119])^(a[356] & b[120])^(a[355] & b[121])^(a[354] & b[122])^(a[353] & b[123])^(a[352] & b[124])^(a[351] & b[125])^(a[350] & b[126])^(a[349] & b[127])^(a[348] & b[128])^(a[347] & b[129])^(a[346] & b[130])^(a[345] & b[131])^(a[344] & b[132])^(a[343] & b[133])^(a[342] & b[134])^(a[341] & b[135])^(a[340] & b[136])^(a[339] & b[137])^(a[338] & b[138])^(a[337] & b[139])^(a[336] & b[140])^(a[335] & b[141])^(a[334] & b[142])^(a[333] & b[143])^(a[332] & b[144])^(a[331] & b[145])^(a[330] & b[146])^(a[329] & b[147])^(a[328] & b[148])^(a[327] & b[149])^(a[326] & b[150])^(a[325] & b[151])^(a[324] & b[152])^(a[323] & b[153])^(a[322] & b[154])^(a[321] & b[155])^(a[320] & b[156])^(a[319] & b[157])^(a[318] & b[158])^(a[317] & b[159])^(a[316] & b[160])^(a[315] & b[161])^(a[314] & b[162])^(a[313] & b[163])^(a[312] & b[164])^(a[311] & b[165])^(a[310] & b[166])^(a[309] & b[167])^(a[308] & b[168])^(a[307] & b[169])^(a[306] & b[170])^(a[305] & b[171])^(a[304] & b[172])^(a[303] & b[173])^(a[302] & b[174])^(a[301] & b[175])^(a[300] & b[176])^(a[299] & b[177])^(a[298] & b[178])^(a[297] & b[179])^(a[296] & b[180])^(a[295] & b[181])^(a[294] & b[182])^(a[293] & b[183])^(a[292] & b[184])^(a[291] & b[185])^(a[290] & b[186])^(a[289] & b[187])^(a[288] & b[188])^(a[287] & b[189])^(a[286] & b[190])^(a[285] & b[191])^(a[284] & b[192])^(a[283] & b[193])^(a[282] & b[194])^(a[281] & b[195])^(a[280] & b[196])^(a[279] & b[197])^(a[278] & b[198])^(a[277] & b[199])^(a[276] & b[200])^(a[275] & b[201])^(a[274] & b[202])^(a[273] & b[203])^(a[272] & b[204])^(a[271] & b[205])^(a[270] & b[206])^(a[269] & b[207])^(a[268] & b[208])^(a[267] & b[209])^(a[266] & b[210])^(a[265] & b[211])^(a[264] & b[212])^(a[263] & b[213])^(a[262] & b[214])^(a[261] & b[215])^(a[260] & b[216])^(a[259] & b[217])^(a[258] & b[218])^(a[257] & b[219])^(a[256] & b[220])^(a[255] & b[221])^(a[254] & b[222])^(a[253] & b[223])^(a[252] & b[224])^(a[251] & b[225])^(a[250] & b[226])^(a[249] & b[227])^(a[248] & b[228])^(a[247] & b[229])^(a[246] & b[230])^(a[245] & b[231])^(a[244] & b[232])^(a[243] & b[233])^(a[242] & b[234])^(a[241] & b[235])^(a[240] & b[236])^(a[239] & b[237])^(a[238] & b[238])^(a[237] & b[239])^(a[236] & b[240])^(a[235] & b[241])^(a[234] & b[242])^(a[233] & b[243])^(a[232] & b[244])^(a[231] & b[245])^(a[230] & b[246])^(a[229] & b[247])^(a[228] & b[248])^(a[227] & b[249])^(a[226] & b[250])^(a[225] & b[251])^(a[224] & b[252])^(a[223] & b[253])^(a[222] & b[254])^(a[221] & b[255])^(a[220] & b[256])^(a[219] & b[257])^(a[218] & b[258])^(a[217] & b[259])^(a[216] & b[260])^(a[215] & b[261])^(a[214] & b[262])^(a[213] & b[263])^(a[212] & b[264])^(a[211] & b[265])^(a[210] & b[266])^(a[209] & b[267])^(a[208] & b[268])^(a[207] & b[269])^(a[206] & b[270])^(a[205] & b[271])^(a[204] & b[272])^(a[203] & b[273])^(a[202] & b[274])^(a[201] & b[275])^(a[200] & b[276])^(a[199] & b[277])^(a[198] & b[278])^(a[197] & b[279])^(a[196] & b[280])^(a[195] & b[281])^(a[194] & b[282])^(a[193] & b[283])^(a[192] & b[284])^(a[191] & b[285])^(a[190] & b[286])^(a[189] & b[287])^(a[188] & b[288])^(a[187] & b[289])^(a[186] & b[290])^(a[185] & b[291])^(a[184] & b[292])^(a[183] & b[293])^(a[182] & b[294])^(a[181] & b[295])^(a[180] & b[296])^(a[179] & b[297])^(a[178] & b[298])^(a[177] & b[299])^(a[176] & b[300])^(a[175] & b[301])^(a[174] & b[302])^(a[173] & b[303])^(a[172] & b[304])^(a[171] & b[305])^(a[170] & b[306])^(a[169] & b[307])^(a[168] & b[308])^(a[167] & b[309])^(a[166] & b[310])^(a[165] & b[311])^(a[164] & b[312])^(a[163] & b[313])^(a[162] & b[314])^(a[161] & b[315])^(a[160] & b[316])^(a[159] & b[317])^(a[158] & b[318])^(a[157] & b[319])^(a[156] & b[320])^(a[155] & b[321])^(a[154] & b[322])^(a[153] & b[323])^(a[152] & b[324])^(a[151] & b[325])^(a[150] & b[326])^(a[149] & b[327])^(a[148] & b[328])^(a[147] & b[329])^(a[146] & b[330])^(a[145] & b[331])^(a[144] & b[332])^(a[143] & b[333])^(a[142] & b[334])^(a[141] & b[335])^(a[140] & b[336])^(a[139] & b[337])^(a[138] & b[338])^(a[137] & b[339])^(a[136] & b[340])^(a[135] & b[341])^(a[134] & b[342])^(a[133] & b[343])^(a[132] & b[344])^(a[131] & b[345])^(a[130] & b[346])^(a[129] & b[347])^(a[128] & b[348])^(a[127] & b[349])^(a[126] & b[350])^(a[125] & b[351])^(a[124] & b[352])^(a[123] & b[353])^(a[122] & b[354])^(a[121] & b[355])^(a[120] & b[356])^(a[119] & b[357])^(a[118] & b[358])^(a[117] & b[359])^(a[116] & b[360])^(a[115] & b[361])^(a[114] & b[362])^(a[113] & b[363])^(a[112] & b[364])^(a[111] & b[365])^(a[110] & b[366])^(a[109] & b[367])^(a[108] & b[368])^(a[107] & b[369])^(a[106] & b[370])^(a[105] & b[371])^(a[104] & b[372])^(a[103] & b[373])^(a[102] & b[374])^(a[101] & b[375])^(a[100] & b[376])^(a[99] & b[377])^(a[98] & b[378])^(a[97] & b[379])^(a[96] & b[380])^(a[95] & b[381])^(a[94] & b[382])^(a[93] & b[383])^(a[92] & b[384])^(a[91] & b[385])^(a[90] & b[386])^(a[89] & b[387])^(a[88] & b[388])^(a[87] & b[389])^(a[86] & b[390])^(a[85] & b[391])^(a[84] & b[392])^(a[83] & b[393])^(a[82] & b[394])^(a[81] & b[395])^(a[80] & b[396])^(a[79] & b[397])^(a[78] & b[398])^(a[77] & b[399])^(a[76] & b[400])^(a[75] & b[401])^(a[74] & b[402])^(a[73] & b[403])^(a[72] & b[404])^(a[71] & b[405])^(a[70] & b[406])^(a[69] & b[407])^(a[68] & b[408]);
assign y[477] = (a[408] & b[69])^(a[407] & b[70])^(a[406] & b[71])^(a[405] & b[72])^(a[404] & b[73])^(a[403] & b[74])^(a[402] & b[75])^(a[401] & b[76])^(a[400] & b[77])^(a[399] & b[78])^(a[398] & b[79])^(a[397] & b[80])^(a[396] & b[81])^(a[395] & b[82])^(a[394] & b[83])^(a[393] & b[84])^(a[392] & b[85])^(a[391] & b[86])^(a[390] & b[87])^(a[389] & b[88])^(a[388] & b[89])^(a[387] & b[90])^(a[386] & b[91])^(a[385] & b[92])^(a[384] & b[93])^(a[383] & b[94])^(a[382] & b[95])^(a[381] & b[96])^(a[380] & b[97])^(a[379] & b[98])^(a[378] & b[99])^(a[377] & b[100])^(a[376] & b[101])^(a[375] & b[102])^(a[374] & b[103])^(a[373] & b[104])^(a[372] & b[105])^(a[371] & b[106])^(a[370] & b[107])^(a[369] & b[108])^(a[368] & b[109])^(a[367] & b[110])^(a[366] & b[111])^(a[365] & b[112])^(a[364] & b[113])^(a[363] & b[114])^(a[362] & b[115])^(a[361] & b[116])^(a[360] & b[117])^(a[359] & b[118])^(a[358] & b[119])^(a[357] & b[120])^(a[356] & b[121])^(a[355] & b[122])^(a[354] & b[123])^(a[353] & b[124])^(a[352] & b[125])^(a[351] & b[126])^(a[350] & b[127])^(a[349] & b[128])^(a[348] & b[129])^(a[347] & b[130])^(a[346] & b[131])^(a[345] & b[132])^(a[344] & b[133])^(a[343] & b[134])^(a[342] & b[135])^(a[341] & b[136])^(a[340] & b[137])^(a[339] & b[138])^(a[338] & b[139])^(a[337] & b[140])^(a[336] & b[141])^(a[335] & b[142])^(a[334] & b[143])^(a[333] & b[144])^(a[332] & b[145])^(a[331] & b[146])^(a[330] & b[147])^(a[329] & b[148])^(a[328] & b[149])^(a[327] & b[150])^(a[326] & b[151])^(a[325] & b[152])^(a[324] & b[153])^(a[323] & b[154])^(a[322] & b[155])^(a[321] & b[156])^(a[320] & b[157])^(a[319] & b[158])^(a[318] & b[159])^(a[317] & b[160])^(a[316] & b[161])^(a[315] & b[162])^(a[314] & b[163])^(a[313] & b[164])^(a[312] & b[165])^(a[311] & b[166])^(a[310] & b[167])^(a[309] & b[168])^(a[308] & b[169])^(a[307] & b[170])^(a[306] & b[171])^(a[305] & b[172])^(a[304] & b[173])^(a[303] & b[174])^(a[302] & b[175])^(a[301] & b[176])^(a[300] & b[177])^(a[299] & b[178])^(a[298] & b[179])^(a[297] & b[180])^(a[296] & b[181])^(a[295] & b[182])^(a[294] & b[183])^(a[293] & b[184])^(a[292] & b[185])^(a[291] & b[186])^(a[290] & b[187])^(a[289] & b[188])^(a[288] & b[189])^(a[287] & b[190])^(a[286] & b[191])^(a[285] & b[192])^(a[284] & b[193])^(a[283] & b[194])^(a[282] & b[195])^(a[281] & b[196])^(a[280] & b[197])^(a[279] & b[198])^(a[278] & b[199])^(a[277] & b[200])^(a[276] & b[201])^(a[275] & b[202])^(a[274] & b[203])^(a[273] & b[204])^(a[272] & b[205])^(a[271] & b[206])^(a[270] & b[207])^(a[269] & b[208])^(a[268] & b[209])^(a[267] & b[210])^(a[266] & b[211])^(a[265] & b[212])^(a[264] & b[213])^(a[263] & b[214])^(a[262] & b[215])^(a[261] & b[216])^(a[260] & b[217])^(a[259] & b[218])^(a[258] & b[219])^(a[257] & b[220])^(a[256] & b[221])^(a[255] & b[222])^(a[254] & b[223])^(a[253] & b[224])^(a[252] & b[225])^(a[251] & b[226])^(a[250] & b[227])^(a[249] & b[228])^(a[248] & b[229])^(a[247] & b[230])^(a[246] & b[231])^(a[245] & b[232])^(a[244] & b[233])^(a[243] & b[234])^(a[242] & b[235])^(a[241] & b[236])^(a[240] & b[237])^(a[239] & b[238])^(a[238] & b[239])^(a[237] & b[240])^(a[236] & b[241])^(a[235] & b[242])^(a[234] & b[243])^(a[233] & b[244])^(a[232] & b[245])^(a[231] & b[246])^(a[230] & b[247])^(a[229] & b[248])^(a[228] & b[249])^(a[227] & b[250])^(a[226] & b[251])^(a[225] & b[252])^(a[224] & b[253])^(a[223] & b[254])^(a[222] & b[255])^(a[221] & b[256])^(a[220] & b[257])^(a[219] & b[258])^(a[218] & b[259])^(a[217] & b[260])^(a[216] & b[261])^(a[215] & b[262])^(a[214] & b[263])^(a[213] & b[264])^(a[212] & b[265])^(a[211] & b[266])^(a[210] & b[267])^(a[209] & b[268])^(a[208] & b[269])^(a[207] & b[270])^(a[206] & b[271])^(a[205] & b[272])^(a[204] & b[273])^(a[203] & b[274])^(a[202] & b[275])^(a[201] & b[276])^(a[200] & b[277])^(a[199] & b[278])^(a[198] & b[279])^(a[197] & b[280])^(a[196] & b[281])^(a[195] & b[282])^(a[194] & b[283])^(a[193] & b[284])^(a[192] & b[285])^(a[191] & b[286])^(a[190] & b[287])^(a[189] & b[288])^(a[188] & b[289])^(a[187] & b[290])^(a[186] & b[291])^(a[185] & b[292])^(a[184] & b[293])^(a[183] & b[294])^(a[182] & b[295])^(a[181] & b[296])^(a[180] & b[297])^(a[179] & b[298])^(a[178] & b[299])^(a[177] & b[300])^(a[176] & b[301])^(a[175] & b[302])^(a[174] & b[303])^(a[173] & b[304])^(a[172] & b[305])^(a[171] & b[306])^(a[170] & b[307])^(a[169] & b[308])^(a[168] & b[309])^(a[167] & b[310])^(a[166] & b[311])^(a[165] & b[312])^(a[164] & b[313])^(a[163] & b[314])^(a[162] & b[315])^(a[161] & b[316])^(a[160] & b[317])^(a[159] & b[318])^(a[158] & b[319])^(a[157] & b[320])^(a[156] & b[321])^(a[155] & b[322])^(a[154] & b[323])^(a[153] & b[324])^(a[152] & b[325])^(a[151] & b[326])^(a[150] & b[327])^(a[149] & b[328])^(a[148] & b[329])^(a[147] & b[330])^(a[146] & b[331])^(a[145] & b[332])^(a[144] & b[333])^(a[143] & b[334])^(a[142] & b[335])^(a[141] & b[336])^(a[140] & b[337])^(a[139] & b[338])^(a[138] & b[339])^(a[137] & b[340])^(a[136] & b[341])^(a[135] & b[342])^(a[134] & b[343])^(a[133] & b[344])^(a[132] & b[345])^(a[131] & b[346])^(a[130] & b[347])^(a[129] & b[348])^(a[128] & b[349])^(a[127] & b[350])^(a[126] & b[351])^(a[125] & b[352])^(a[124] & b[353])^(a[123] & b[354])^(a[122] & b[355])^(a[121] & b[356])^(a[120] & b[357])^(a[119] & b[358])^(a[118] & b[359])^(a[117] & b[360])^(a[116] & b[361])^(a[115] & b[362])^(a[114] & b[363])^(a[113] & b[364])^(a[112] & b[365])^(a[111] & b[366])^(a[110] & b[367])^(a[109] & b[368])^(a[108] & b[369])^(a[107] & b[370])^(a[106] & b[371])^(a[105] & b[372])^(a[104] & b[373])^(a[103] & b[374])^(a[102] & b[375])^(a[101] & b[376])^(a[100] & b[377])^(a[99] & b[378])^(a[98] & b[379])^(a[97] & b[380])^(a[96] & b[381])^(a[95] & b[382])^(a[94] & b[383])^(a[93] & b[384])^(a[92] & b[385])^(a[91] & b[386])^(a[90] & b[387])^(a[89] & b[388])^(a[88] & b[389])^(a[87] & b[390])^(a[86] & b[391])^(a[85] & b[392])^(a[84] & b[393])^(a[83] & b[394])^(a[82] & b[395])^(a[81] & b[396])^(a[80] & b[397])^(a[79] & b[398])^(a[78] & b[399])^(a[77] & b[400])^(a[76] & b[401])^(a[75] & b[402])^(a[74] & b[403])^(a[73] & b[404])^(a[72] & b[405])^(a[71] & b[406])^(a[70] & b[407])^(a[69] & b[408]);
assign y[478] = (a[408] & b[70])^(a[407] & b[71])^(a[406] & b[72])^(a[405] & b[73])^(a[404] & b[74])^(a[403] & b[75])^(a[402] & b[76])^(a[401] & b[77])^(a[400] & b[78])^(a[399] & b[79])^(a[398] & b[80])^(a[397] & b[81])^(a[396] & b[82])^(a[395] & b[83])^(a[394] & b[84])^(a[393] & b[85])^(a[392] & b[86])^(a[391] & b[87])^(a[390] & b[88])^(a[389] & b[89])^(a[388] & b[90])^(a[387] & b[91])^(a[386] & b[92])^(a[385] & b[93])^(a[384] & b[94])^(a[383] & b[95])^(a[382] & b[96])^(a[381] & b[97])^(a[380] & b[98])^(a[379] & b[99])^(a[378] & b[100])^(a[377] & b[101])^(a[376] & b[102])^(a[375] & b[103])^(a[374] & b[104])^(a[373] & b[105])^(a[372] & b[106])^(a[371] & b[107])^(a[370] & b[108])^(a[369] & b[109])^(a[368] & b[110])^(a[367] & b[111])^(a[366] & b[112])^(a[365] & b[113])^(a[364] & b[114])^(a[363] & b[115])^(a[362] & b[116])^(a[361] & b[117])^(a[360] & b[118])^(a[359] & b[119])^(a[358] & b[120])^(a[357] & b[121])^(a[356] & b[122])^(a[355] & b[123])^(a[354] & b[124])^(a[353] & b[125])^(a[352] & b[126])^(a[351] & b[127])^(a[350] & b[128])^(a[349] & b[129])^(a[348] & b[130])^(a[347] & b[131])^(a[346] & b[132])^(a[345] & b[133])^(a[344] & b[134])^(a[343] & b[135])^(a[342] & b[136])^(a[341] & b[137])^(a[340] & b[138])^(a[339] & b[139])^(a[338] & b[140])^(a[337] & b[141])^(a[336] & b[142])^(a[335] & b[143])^(a[334] & b[144])^(a[333] & b[145])^(a[332] & b[146])^(a[331] & b[147])^(a[330] & b[148])^(a[329] & b[149])^(a[328] & b[150])^(a[327] & b[151])^(a[326] & b[152])^(a[325] & b[153])^(a[324] & b[154])^(a[323] & b[155])^(a[322] & b[156])^(a[321] & b[157])^(a[320] & b[158])^(a[319] & b[159])^(a[318] & b[160])^(a[317] & b[161])^(a[316] & b[162])^(a[315] & b[163])^(a[314] & b[164])^(a[313] & b[165])^(a[312] & b[166])^(a[311] & b[167])^(a[310] & b[168])^(a[309] & b[169])^(a[308] & b[170])^(a[307] & b[171])^(a[306] & b[172])^(a[305] & b[173])^(a[304] & b[174])^(a[303] & b[175])^(a[302] & b[176])^(a[301] & b[177])^(a[300] & b[178])^(a[299] & b[179])^(a[298] & b[180])^(a[297] & b[181])^(a[296] & b[182])^(a[295] & b[183])^(a[294] & b[184])^(a[293] & b[185])^(a[292] & b[186])^(a[291] & b[187])^(a[290] & b[188])^(a[289] & b[189])^(a[288] & b[190])^(a[287] & b[191])^(a[286] & b[192])^(a[285] & b[193])^(a[284] & b[194])^(a[283] & b[195])^(a[282] & b[196])^(a[281] & b[197])^(a[280] & b[198])^(a[279] & b[199])^(a[278] & b[200])^(a[277] & b[201])^(a[276] & b[202])^(a[275] & b[203])^(a[274] & b[204])^(a[273] & b[205])^(a[272] & b[206])^(a[271] & b[207])^(a[270] & b[208])^(a[269] & b[209])^(a[268] & b[210])^(a[267] & b[211])^(a[266] & b[212])^(a[265] & b[213])^(a[264] & b[214])^(a[263] & b[215])^(a[262] & b[216])^(a[261] & b[217])^(a[260] & b[218])^(a[259] & b[219])^(a[258] & b[220])^(a[257] & b[221])^(a[256] & b[222])^(a[255] & b[223])^(a[254] & b[224])^(a[253] & b[225])^(a[252] & b[226])^(a[251] & b[227])^(a[250] & b[228])^(a[249] & b[229])^(a[248] & b[230])^(a[247] & b[231])^(a[246] & b[232])^(a[245] & b[233])^(a[244] & b[234])^(a[243] & b[235])^(a[242] & b[236])^(a[241] & b[237])^(a[240] & b[238])^(a[239] & b[239])^(a[238] & b[240])^(a[237] & b[241])^(a[236] & b[242])^(a[235] & b[243])^(a[234] & b[244])^(a[233] & b[245])^(a[232] & b[246])^(a[231] & b[247])^(a[230] & b[248])^(a[229] & b[249])^(a[228] & b[250])^(a[227] & b[251])^(a[226] & b[252])^(a[225] & b[253])^(a[224] & b[254])^(a[223] & b[255])^(a[222] & b[256])^(a[221] & b[257])^(a[220] & b[258])^(a[219] & b[259])^(a[218] & b[260])^(a[217] & b[261])^(a[216] & b[262])^(a[215] & b[263])^(a[214] & b[264])^(a[213] & b[265])^(a[212] & b[266])^(a[211] & b[267])^(a[210] & b[268])^(a[209] & b[269])^(a[208] & b[270])^(a[207] & b[271])^(a[206] & b[272])^(a[205] & b[273])^(a[204] & b[274])^(a[203] & b[275])^(a[202] & b[276])^(a[201] & b[277])^(a[200] & b[278])^(a[199] & b[279])^(a[198] & b[280])^(a[197] & b[281])^(a[196] & b[282])^(a[195] & b[283])^(a[194] & b[284])^(a[193] & b[285])^(a[192] & b[286])^(a[191] & b[287])^(a[190] & b[288])^(a[189] & b[289])^(a[188] & b[290])^(a[187] & b[291])^(a[186] & b[292])^(a[185] & b[293])^(a[184] & b[294])^(a[183] & b[295])^(a[182] & b[296])^(a[181] & b[297])^(a[180] & b[298])^(a[179] & b[299])^(a[178] & b[300])^(a[177] & b[301])^(a[176] & b[302])^(a[175] & b[303])^(a[174] & b[304])^(a[173] & b[305])^(a[172] & b[306])^(a[171] & b[307])^(a[170] & b[308])^(a[169] & b[309])^(a[168] & b[310])^(a[167] & b[311])^(a[166] & b[312])^(a[165] & b[313])^(a[164] & b[314])^(a[163] & b[315])^(a[162] & b[316])^(a[161] & b[317])^(a[160] & b[318])^(a[159] & b[319])^(a[158] & b[320])^(a[157] & b[321])^(a[156] & b[322])^(a[155] & b[323])^(a[154] & b[324])^(a[153] & b[325])^(a[152] & b[326])^(a[151] & b[327])^(a[150] & b[328])^(a[149] & b[329])^(a[148] & b[330])^(a[147] & b[331])^(a[146] & b[332])^(a[145] & b[333])^(a[144] & b[334])^(a[143] & b[335])^(a[142] & b[336])^(a[141] & b[337])^(a[140] & b[338])^(a[139] & b[339])^(a[138] & b[340])^(a[137] & b[341])^(a[136] & b[342])^(a[135] & b[343])^(a[134] & b[344])^(a[133] & b[345])^(a[132] & b[346])^(a[131] & b[347])^(a[130] & b[348])^(a[129] & b[349])^(a[128] & b[350])^(a[127] & b[351])^(a[126] & b[352])^(a[125] & b[353])^(a[124] & b[354])^(a[123] & b[355])^(a[122] & b[356])^(a[121] & b[357])^(a[120] & b[358])^(a[119] & b[359])^(a[118] & b[360])^(a[117] & b[361])^(a[116] & b[362])^(a[115] & b[363])^(a[114] & b[364])^(a[113] & b[365])^(a[112] & b[366])^(a[111] & b[367])^(a[110] & b[368])^(a[109] & b[369])^(a[108] & b[370])^(a[107] & b[371])^(a[106] & b[372])^(a[105] & b[373])^(a[104] & b[374])^(a[103] & b[375])^(a[102] & b[376])^(a[101] & b[377])^(a[100] & b[378])^(a[99] & b[379])^(a[98] & b[380])^(a[97] & b[381])^(a[96] & b[382])^(a[95] & b[383])^(a[94] & b[384])^(a[93] & b[385])^(a[92] & b[386])^(a[91] & b[387])^(a[90] & b[388])^(a[89] & b[389])^(a[88] & b[390])^(a[87] & b[391])^(a[86] & b[392])^(a[85] & b[393])^(a[84] & b[394])^(a[83] & b[395])^(a[82] & b[396])^(a[81] & b[397])^(a[80] & b[398])^(a[79] & b[399])^(a[78] & b[400])^(a[77] & b[401])^(a[76] & b[402])^(a[75] & b[403])^(a[74] & b[404])^(a[73] & b[405])^(a[72] & b[406])^(a[71] & b[407])^(a[70] & b[408]);
assign y[479] = (a[408] & b[71])^(a[407] & b[72])^(a[406] & b[73])^(a[405] & b[74])^(a[404] & b[75])^(a[403] & b[76])^(a[402] & b[77])^(a[401] & b[78])^(a[400] & b[79])^(a[399] & b[80])^(a[398] & b[81])^(a[397] & b[82])^(a[396] & b[83])^(a[395] & b[84])^(a[394] & b[85])^(a[393] & b[86])^(a[392] & b[87])^(a[391] & b[88])^(a[390] & b[89])^(a[389] & b[90])^(a[388] & b[91])^(a[387] & b[92])^(a[386] & b[93])^(a[385] & b[94])^(a[384] & b[95])^(a[383] & b[96])^(a[382] & b[97])^(a[381] & b[98])^(a[380] & b[99])^(a[379] & b[100])^(a[378] & b[101])^(a[377] & b[102])^(a[376] & b[103])^(a[375] & b[104])^(a[374] & b[105])^(a[373] & b[106])^(a[372] & b[107])^(a[371] & b[108])^(a[370] & b[109])^(a[369] & b[110])^(a[368] & b[111])^(a[367] & b[112])^(a[366] & b[113])^(a[365] & b[114])^(a[364] & b[115])^(a[363] & b[116])^(a[362] & b[117])^(a[361] & b[118])^(a[360] & b[119])^(a[359] & b[120])^(a[358] & b[121])^(a[357] & b[122])^(a[356] & b[123])^(a[355] & b[124])^(a[354] & b[125])^(a[353] & b[126])^(a[352] & b[127])^(a[351] & b[128])^(a[350] & b[129])^(a[349] & b[130])^(a[348] & b[131])^(a[347] & b[132])^(a[346] & b[133])^(a[345] & b[134])^(a[344] & b[135])^(a[343] & b[136])^(a[342] & b[137])^(a[341] & b[138])^(a[340] & b[139])^(a[339] & b[140])^(a[338] & b[141])^(a[337] & b[142])^(a[336] & b[143])^(a[335] & b[144])^(a[334] & b[145])^(a[333] & b[146])^(a[332] & b[147])^(a[331] & b[148])^(a[330] & b[149])^(a[329] & b[150])^(a[328] & b[151])^(a[327] & b[152])^(a[326] & b[153])^(a[325] & b[154])^(a[324] & b[155])^(a[323] & b[156])^(a[322] & b[157])^(a[321] & b[158])^(a[320] & b[159])^(a[319] & b[160])^(a[318] & b[161])^(a[317] & b[162])^(a[316] & b[163])^(a[315] & b[164])^(a[314] & b[165])^(a[313] & b[166])^(a[312] & b[167])^(a[311] & b[168])^(a[310] & b[169])^(a[309] & b[170])^(a[308] & b[171])^(a[307] & b[172])^(a[306] & b[173])^(a[305] & b[174])^(a[304] & b[175])^(a[303] & b[176])^(a[302] & b[177])^(a[301] & b[178])^(a[300] & b[179])^(a[299] & b[180])^(a[298] & b[181])^(a[297] & b[182])^(a[296] & b[183])^(a[295] & b[184])^(a[294] & b[185])^(a[293] & b[186])^(a[292] & b[187])^(a[291] & b[188])^(a[290] & b[189])^(a[289] & b[190])^(a[288] & b[191])^(a[287] & b[192])^(a[286] & b[193])^(a[285] & b[194])^(a[284] & b[195])^(a[283] & b[196])^(a[282] & b[197])^(a[281] & b[198])^(a[280] & b[199])^(a[279] & b[200])^(a[278] & b[201])^(a[277] & b[202])^(a[276] & b[203])^(a[275] & b[204])^(a[274] & b[205])^(a[273] & b[206])^(a[272] & b[207])^(a[271] & b[208])^(a[270] & b[209])^(a[269] & b[210])^(a[268] & b[211])^(a[267] & b[212])^(a[266] & b[213])^(a[265] & b[214])^(a[264] & b[215])^(a[263] & b[216])^(a[262] & b[217])^(a[261] & b[218])^(a[260] & b[219])^(a[259] & b[220])^(a[258] & b[221])^(a[257] & b[222])^(a[256] & b[223])^(a[255] & b[224])^(a[254] & b[225])^(a[253] & b[226])^(a[252] & b[227])^(a[251] & b[228])^(a[250] & b[229])^(a[249] & b[230])^(a[248] & b[231])^(a[247] & b[232])^(a[246] & b[233])^(a[245] & b[234])^(a[244] & b[235])^(a[243] & b[236])^(a[242] & b[237])^(a[241] & b[238])^(a[240] & b[239])^(a[239] & b[240])^(a[238] & b[241])^(a[237] & b[242])^(a[236] & b[243])^(a[235] & b[244])^(a[234] & b[245])^(a[233] & b[246])^(a[232] & b[247])^(a[231] & b[248])^(a[230] & b[249])^(a[229] & b[250])^(a[228] & b[251])^(a[227] & b[252])^(a[226] & b[253])^(a[225] & b[254])^(a[224] & b[255])^(a[223] & b[256])^(a[222] & b[257])^(a[221] & b[258])^(a[220] & b[259])^(a[219] & b[260])^(a[218] & b[261])^(a[217] & b[262])^(a[216] & b[263])^(a[215] & b[264])^(a[214] & b[265])^(a[213] & b[266])^(a[212] & b[267])^(a[211] & b[268])^(a[210] & b[269])^(a[209] & b[270])^(a[208] & b[271])^(a[207] & b[272])^(a[206] & b[273])^(a[205] & b[274])^(a[204] & b[275])^(a[203] & b[276])^(a[202] & b[277])^(a[201] & b[278])^(a[200] & b[279])^(a[199] & b[280])^(a[198] & b[281])^(a[197] & b[282])^(a[196] & b[283])^(a[195] & b[284])^(a[194] & b[285])^(a[193] & b[286])^(a[192] & b[287])^(a[191] & b[288])^(a[190] & b[289])^(a[189] & b[290])^(a[188] & b[291])^(a[187] & b[292])^(a[186] & b[293])^(a[185] & b[294])^(a[184] & b[295])^(a[183] & b[296])^(a[182] & b[297])^(a[181] & b[298])^(a[180] & b[299])^(a[179] & b[300])^(a[178] & b[301])^(a[177] & b[302])^(a[176] & b[303])^(a[175] & b[304])^(a[174] & b[305])^(a[173] & b[306])^(a[172] & b[307])^(a[171] & b[308])^(a[170] & b[309])^(a[169] & b[310])^(a[168] & b[311])^(a[167] & b[312])^(a[166] & b[313])^(a[165] & b[314])^(a[164] & b[315])^(a[163] & b[316])^(a[162] & b[317])^(a[161] & b[318])^(a[160] & b[319])^(a[159] & b[320])^(a[158] & b[321])^(a[157] & b[322])^(a[156] & b[323])^(a[155] & b[324])^(a[154] & b[325])^(a[153] & b[326])^(a[152] & b[327])^(a[151] & b[328])^(a[150] & b[329])^(a[149] & b[330])^(a[148] & b[331])^(a[147] & b[332])^(a[146] & b[333])^(a[145] & b[334])^(a[144] & b[335])^(a[143] & b[336])^(a[142] & b[337])^(a[141] & b[338])^(a[140] & b[339])^(a[139] & b[340])^(a[138] & b[341])^(a[137] & b[342])^(a[136] & b[343])^(a[135] & b[344])^(a[134] & b[345])^(a[133] & b[346])^(a[132] & b[347])^(a[131] & b[348])^(a[130] & b[349])^(a[129] & b[350])^(a[128] & b[351])^(a[127] & b[352])^(a[126] & b[353])^(a[125] & b[354])^(a[124] & b[355])^(a[123] & b[356])^(a[122] & b[357])^(a[121] & b[358])^(a[120] & b[359])^(a[119] & b[360])^(a[118] & b[361])^(a[117] & b[362])^(a[116] & b[363])^(a[115] & b[364])^(a[114] & b[365])^(a[113] & b[366])^(a[112] & b[367])^(a[111] & b[368])^(a[110] & b[369])^(a[109] & b[370])^(a[108] & b[371])^(a[107] & b[372])^(a[106] & b[373])^(a[105] & b[374])^(a[104] & b[375])^(a[103] & b[376])^(a[102] & b[377])^(a[101] & b[378])^(a[100] & b[379])^(a[99] & b[380])^(a[98] & b[381])^(a[97] & b[382])^(a[96] & b[383])^(a[95] & b[384])^(a[94] & b[385])^(a[93] & b[386])^(a[92] & b[387])^(a[91] & b[388])^(a[90] & b[389])^(a[89] & b[390])^(a[88] & b[391])^(a[87] & b[392])^(a[86] & b[393])^(a[85] & b[394])^(a[84] & b[395])^(a[83] & b[396])^(a[82] & b[397])^(a[81] & b[398])^(a[80] & b[399])^(a[79] & b[400])^(a[78] & b[401])^(a[77] & b[402])^(a[76] & b[403])^(a[75] & b[404])^(a[74] & b[405])^(a[73] & b[406])^(a[72] & b[407])^(a[71] & b[408]);
assign y[480] = (a[408] & b[72])^(a[407] & b[73])^(a[406] & b[74])^(a[405] & b[75])^(a[404] & b[76])^(a[403] & b[77])^(a[402] & b[78])^(a[401] & b[79])^(a[400] & b[80])^(a[399] & b[81])^(a[398] & b[82])^(a[397] & b[83])^(a[396] & b[84])^(a[395] & b[85])^(a[394] & b[86])^(a[393] & b[87])^(a[392] & b[88])^(a[391] & b[89])^(a[390] & b[90])^(a[389] & b[91])^(a[388] & b[92])^(a[387] & b[93])^(a[386] & b[94])^(a[385] & b[95])^(a[384] & b[96])^(a[383] & b[97])^(a[382] & b[98])^(a[381] & b[99])^(a[380] & b[100])^(a[379] & b[101])^(a[378] & b[102])^(a[377] & b[103])^(a[376] & b[104])^(a[375] & b[105])^(a[374] & b[106])^(a[373] & b[107])^(a[372] & b[108])^(a[371] & b[109])^(a[370] & b[110])^(a[369] & b[111])^(a[368] & b[112])^(a[367] & b[113])^(a[366] & b[114])^(a[365] & b[115])^(a[364] & b[116])^(a[363] & b[117])^(a[362] & b[118])^(a[361] & b[119])^(a[360] & b[120])^(a[359] & b[121])^(a[358] & b[122])^(a[357] & b[123])^(a[356] & b[124])^(a[355] & b[125])^(a[354] & b[126])^(a[353] & b[127])^(a[352] & b[128])^(a[351] & b[129])^(a[350] & b[130])^(a[349] & b[131])^(a[348] & b[132])^(a[347] & b[133])^(a[346] & b[134])^(a[345] & b[135])^(a[344] & b[136])^(a[343] & b[137])^(a[342] & b[138])^(a[341] & b[139])^(a[340] & b[140])^(a[339] & b[141])^(a[338] & b[142])^(a[337] & b[143])^(a[336] & b[144])^(a[335] & b[145])^(a[334] & b[146])^(a[333] & b[147])^(a[332] & b[148])^(a[331] & b[149])^(a[330] & b[150])^(a[329] & b[151])^(a[328] & b[152])^(a[327] & b[153])^(a[326] & b[154])^(a[325] & b[155])^(a[324] & b[156])^(a[323] & b[157])^(a[322] & b[158])^(a[321] & b[159])^(a[320] & b[160])^(a[319] & b[161])^(a[318] & b[162])^(a[317] & b[163])^(a[316] & b[164])^(a[315] & b[165])^(a[314] & b[166])^(a[313] & b[167])^(a[312] & b[168])^(a[311] & b[169])^(a[310] & b[170])^(a[309] & b[171])^(a[308] & b[172])^(a[307] & b[173])^(a[306] & b[174])^(a[305] & b[175])^(a[304] & b[176])^(a[303] & b[177])^(a[302] & b[178])^(a[301] & b[179])^(a[300] & b[180])^(a[299] & b[181])^(a[298] & b[182])^(a[297] & b[183])^(a[296] & b[184])^(a[295] & b[185])^(a[294] & b[186])^(a[293] & b[187])^(a[292] & b[188])^(a[291] & b[189])^(a[290] & b[190])^(a[289] & b[191])^(a[288] & b[192])^(a[287] & b[193])^(a[286] & b[194])^(a[285] & b[195])^(a[284] & b[196])^(a[283] & b[197])^(a[282] & b[198])^(a[281] & b[199])^(a[280] & b[200])^(a[279] & b[201])^(a[278] & b[202])^(a[277] & b[203])^(a[276] & b[204])^(a[275] & b[205])^(a[274] & b[206])^(a[273] & b[207])^(a[272] & b[208])^(a[271] & b[209])^(a[270] & b[210])^(a[269] & b[211])^(a[268] & b[212])^(a[267] & b[213])^(a[266] & b[214])^(a[265] & b[215])^(a[264] & b[216])^(a[263] & b[217])^(a[262] & b[218])^(a[261] & b[219])^(a[260] & b[220])^(a[259] & b[221])^(a[258] & b[222])^(a[257] & b[223])^(a[256] & b[224])^(a[255] & b[225])^(a[254] & b[226])^(a[253] & b[227])^(a[252] & b[228])^(a[251] & b[229])^(a[250] & b[230])^(a[249] & b[231])^(a[248] & b[232])^(a[247] & b[233])^(a[246] & b[234])^(a[245] & b[235])^(a[244] & b[236])^(a[243] & b[237])^(a[242] & b[238])^(a[241] & b[239])^(a[240] & b[240])^(a[239] & b[241])^(a[238] & b[242])^(a[237] & b[243])^(a[236] & b[244])^(a[235] & b[245])^(a[234] & b[246])^(a[233] & b[247])^(a[232] & b[248])^(a[231] & b[249])^(a[230] & b[250])^(a[229] & b[251])^(a[228] & b[252])^(a[227] & b[253])^(a[226] & b[254])^(a[225] & b[255])^(a[224] & b[256])^(a[223] & b[257])^(a[222] & b[258])^(a[221] & b[259])^(a[220] & b[260])^(a[219] & b[261])^(a[218] & b[262])^(a[217] & b[263])^(a[216] & b[264])^(a[215] & b[265])^(a[214] & b[266])^(a[213] & b[267])^(a[212] & b[268])^(a[211] & b[269])^(a[210] & b[270])^(a[209] & b[271])^(a[208] & b[272])^(a[207] & b[273])^(a[206] & b[274])^(a[205] & b[275])^(a[204] & b[276])^(a[203] & b[277])^(a[202] & b[278])^(a[201] & b[279])^(a[200] & b[280])^(a[199] & b[281])^(a[198] & b[282])^(a[197] & b[283])^(a[196] & b[284])^(a[195] & b[285])^(a[194] & b[286])^(a[193] & b[287])^(a[192] & b[288])^(a[191] & b[289])^(a[190] & b[290])^(a[189] & b[291])^(a[188] & b[292])^(a[187] & b[293])^(a[186] & b[294])^(a[185] & b[295])^(a[184] & b[296])^(a[183] & b[297])^(a[182] & b[298])^(a[181] & b[299])^(a[180] & b[300])^(a[179] & b[301])^(a[178] & b[302])^(a[177] & b[303])^(a[176] & b[304])^(a[175] & b[305])^(a[174] & b[306])^(a[173] & b[307])^(a[172] & b[308])^(a[171] & b[309])^(a[170] & b[310])^(a[169] & b[311])^(a[168] & b[312])^(a[167] & b[313])^(a[166] & b[314])^(a[165] & b[315])^(a[164] & b[316])^(a[163] & b[317])^(a[162] & b[318])^(a[161] & b[319])^(a[160] & b[320])^(a[159] & b[321])^(a[158] & b[322])^(a[157] & b[323])^(a[156] & b[324])^(a[155] & b[325])^(a[154] & b[326])^(a[153] & b[327])^(a[152] & b[328])^(a[151] & b[329])^(a[150] & b[330])^(a[149] & b[331])^(a[148] & b[332])^(a[147] & b[333])^(a[146] & b[334])^(a[145] & b[335])^(a[144] & b[336])^(a[143] & b[337])^(a[142] & b[338])^(a[141] & b[339])^(a[140] & b[340])^(a[139] & b[341])^(a[138] & b[342])^(a[137] & b[343])^(a[136] & b[344])^(a[135] & b[345])^(a[134] & b[346])^(a[133] & b[347])^(a[132] & b[348])^(a[131] & b[349])^(a[130] & b[350])^(a[129] & b[351])^(a[128] & b[352])^(a[127] & b[353])^(a[126] & b[354])^(a[125] & b[355])^(a[124] & b[356])^(a[123] & b[357])^(a[122] & b[358])^(a[121] & b[359])^(a[120] & b[360])^(a[119] & b[361])^(a[118] & b[362])^(a[117] & b[363])^(a[116] & b[364])^(a[115] & b[365])^(a[114] & b[366])^(a[113] & b[367])^(a[112] & b[368])^(a[111] & b[369])^(a[110] & b[370])^(a[109] & b[371])^(a[108] & b[372])^(a[107] & b[373])^(a[106] & b[374])^(a[105] & b[375])^(a[104] & b[376])^(a[103] & b[377])^(a[102] & b[378])^(a[101] & b[379])^(a[100] & b[380])^(a[99] & b[381])^(a[98] & b[382])^(a[97] & b[383])^(a[96] & b[384])^(a[95] & b[385])^(a[94] & b[386])^(a[93] & b[387])^(a[92] & b[388])^(a[91] & b[389])^(a[90] & b[390])^(a[89] & b[391])^(a[88] & b[392])^(a[87] & b[393])^(a[86] & b[394])^(a[85] & b[395])^(a[84] & b[396])^(a[83] & b[397])^(a[82] & b[398])^(a[81] & b[399])^(a[80] & b[400])^(a[79] & b[401])^(a[78] & b[402])^(a[77] & b[403])^(a[76] & b[404])^(a[75] & b[405])^(a[74] & b[406])^(a[73] & b[407])^(a[72] & b[408]);
assign y[481] = (a[408] & b[73])^(a[407] & b[74])^(a[406] & b[75])^(a[405] & b[76])^(a[404] & b[77])^(a[403] & b[78])^(a[402] & b[79])^(a[401] & b[80])^(a[400] & b[81])^(a[399] & b[82])^(a[398] & b[83])^(a[397] & b[84])^(a[396] & b[85])^(a[395] & b[86])^(a[394] & b[87])^(a[393] & b[88])^(a[392] & b[89])^(a[391] & b[90])^(a[390] & b[91])^(a[389] & b[92])^(a[388] & b[93])^(a[387] & b[94])^(a[386] & b[95])^(a[385] & b[96])^(a[384] & b[97])^(a[383] & b[98])^(a[382] & b[99])^(a[381] & b[100])^(a[380] & b[101])^(a[379] & b[102])^(a[378] & b[103])^(a[377] & b[104])^(a[376] & b[105])^(a[375] & b[106])^(a[374] & b[107])^(a[373] & b[108])^(a[372] & b[109])^(a[371] & b[110])^(a[370] & b[111])^(a[369] & b[112])^(a[368] & b[113])^(a[367] & b[114])^(a[366] & b[115])^(a[365] & b[116])^(a[364] & b[117])^(a[363] & b[118])^(a[362] & b[119])^(a[361] & b[120])^(a[360] & b[121])^(a[359] & b[122])^(a[358] & b[123])^(a[357] & b[124])^(a[356] & b[125])^(a[355] & b[126])^(a[354] & b[127])^(a[353] & b[128])^(a[352] & b[129])^(a[351] & b[130])^(a[350] & b[131])^(a[349] & b[132])^(a[348] & b[133])^(a[347] & b[134])^(a[346] & b[135])^(a[345] & b[136])^(a[344] & b[137])^(a[343] & b[138])^(a[342] & b[139])^(a[341] & b[140])^(a[340] & b[141])^(a[339] & b[142])^(a[338] & b[143])^(a[337] & b[144])^(a[336] & b[145])^(a[335] & b[146])^(a[334] & b[147])^(a[333] & b[148])^(a[332] & b[149])^(a[331] & b[150])^(a[330] & b[151])^(a[329] & b[152])^(a[328] & b[153])^(a[327] & b[154])^(a[326] & b[155])^(a[325] & b[156])^(a[324] & b[157])^(a[323] & b[158])^(a[322] & b[159])^(a[321] & b[160])^(a[320] & b[161])^(a[319] & b[162])^(a[318] & b[163])^(a[317] & b[164])^(a[316] & b[165])^(a[315] & b[166])^(a[314] & b[167])^(a[313] & b[168])^(a[312] & b[169])^(a[311] & b[170])^(a[310] & b[171])^(a[309] & b[172])^(a[308] & b[173])^(a[307] & b[174])^(a[306] & b[175])^(a[305] & b[176])^(a[304] & b[177])^(a[303] & b[178])^(a[302] & b[179])^(a[301] & b[180])^(a[300] & b[181])^(a[299] & b[182])^(a[298] & b[183])^(a[297] & b[184])^(a[296] & b[185])^(a[295] & b[186])^(a[294] & b[187])^(a[293] & b[188])^(a[292] & b[189])^(a[291] & b[190])^(a[290] & b[191])^(a[289] & b[192])^(a[288] & b[193])^(a[287] & b[194])^(a[286] & b[195])^(a[285] & b[196])^(a[284] & b[197])^(a[283] & b[198])^(a[282] & b[199])^(a[281] & b[200])^(a[280] & b[201])^(a[279] & b[202])^(a[278] & b[203])^(a[277] & b[204])^(a[276] & b[205])^(a[275] & b[206])^(a[274] & b[207])^(a[273] & b[208])^(a[272] & b[209])^(a[271] & b[210])^(a[270] & b[211])^(a[269] & b[212])^(a[268] & b[213])^(a[267] & b[214])^(a[266] & b[215])^(a[265] & b[216])^(a[264] & b[217])^(a[263] & b[218])^(a[262] & b[219])^(a[261] & b[220])^(a[260] & b[221])^(a[259] & b[222])^(a[258] & b[223])^(a[257] & b[224])^(a[256] & b[225])^(a[255] & b[226])^(a[254] & b[227])^(a[253] & b[228])^(a[252] & b[229])^(a[251] & b[230])^(a[250] & b[231])^(a[249] & b[232])^(a[248] & b[233])^(a[247] & b[234])^(a[246] & b[235])^(a[245] & b[236])^(a[244] & b[237])^(a[243] & b[238])^(a[242] & b[239])^(a[241] & b[240])^(a[240] & b[241])^(a[239] & b[242])^(a[238] & b[243])^(a[237] & b[244])^(a[236] & b[245])^(a[235] & b[246])^(a[234] & b[247])^(a[233] & b[248])^(a[232] & b[249])^(a[231] & b[250])^(a[230] & b[251])^(a[229] & b[252])^(a[228] & b[253])^(a[227] & b[254])^(a[226] & b[255])^(a[225] & b[256])^(a[224] & b[257])^(a[223] & b[258])^(a[222] & b[259])^(a[221] & b[260])^(a[220] & b[261])^(a[219] & b[262])^(a[218] & b[263])^(a[217] & b[264])^(a[216] & b[265])^(a[215] & b[266])^(a[214] & b[267])^(a[213] & b[268])^(a[212] & b[269])^(a[211] & b[270])^(a[210] & b[271])^(a[209] & b[272])^(a[208] & b[273])^(a[207] & b[274])^(a[206] & b[275])^(a[205] & b[276])^(a[204] & b[277])^(a[203] & b[278])^(a[202] & b[279])^(a[201] & b[280])^(a[200] & b[281])^(a[199] & b[282])^(a[198] & b[283])^(a[197] & b[284])^(a[196] & b[285])^(a[195] & b[286])^(a[194] & b[287])^(a[193] & b[288])^(a[192] & b[289])^(a[191] & b[290])^(a[190] & b[291])^(a[189] & b[292])^(a[188] & b[293])^(a[187] & b[294])^(a[186] & b[295])^(a[185] & b[296])^(a[184] & b[297])^(a[183] & b[298])^(a[182] & b[299])^(a[181] & b[300])^(a[180] & b[301])^(a[179] & b[302])^(a[178] & b[303])^(a[177] & b[304])^(a[176] & b[305])^(a[175] & b[306])^(a[174] & b[307])^(a[173] & b[308])^(a[172] & b[309])^(a[171] & b[310])^(a[170] & b[311])^(a[169] & b[312])^(a[168] & b[313])^(a[167] & b[314])^(a[166] & b[315])^(a[165] & b[316])^(a[164] & b[317])^(a[163] & b[318])^(a[162] & b[319])^(a[161] & b[320])^(a[160] & b[321])^(a[159] & b[322])^(a[158] & b[323])^(a[157] & b[324])^(a[156] & b[325])^(a[155] & b[326])^(a[154] & b[327])^(a[153] & b[328])^(a[152] & b[329])^(a[151] & b[330])^(a[150] & b[331])^(a[149] & b[332])^(a[148] & b[333])^(a[147] & b[334])^(a[146] & b[335])^(a[145] & b[336])^(a[144] & b[337])^(a[143] & b[338])^(a[142] & b[339])^(a[141] & b[340])^(a[140] & b[341])^(a[139] & b[342])^(a[138] & b[343])^(a[137] & b[344])^(a[136] & b[345])^(a[135] & b[346])^(a[134] & b[347])^(a[133] & b[348])^(a[132] & b[349])^(a[131] & b[350])^(a[130] & b[351])^(a[129] & b[352])^(a[128] & b[353])^(a[127] & b[354])^(a[126] & b[355])^(a[125] & b[356])^(a[124] & b[357])^(a[123] & b[358])^(a[122] & b[359])^(a[121] & b[360])^(a[120] & b[361])^(a[119] & b[362])^(a[118] & b[363])^(a[117] & b[364])^(a[116] & b[365])^(a[115] & b[366])^(a[114] & b[367])^(a[113] & b[368])^(a[112] & b[369])^(a[111] & b[370])^(a[110] & b[371])^(a[109] & b[372])^(a[108] & b[373])^(a[107] & b[374])^(a[106] & b[375])^(a[105] & b[376])^(a[104] & b[377])^(a[103] & b[378])^(a[102] & b[379])^(a[101] & b[380])^(a[100] & b[381])^(a[99] & b[382])^(a[98] & b[383])^(a[97] & b[384])^(a[96] & b[385])^(a[95] & b[386])^(a[94] & b[387])^(a[93] & b[388])^(a[92] & b[389])^(a[91] & b[390])^(a[90] & b[391])^(a[89] & b[392])^(a[88] & b[393])^(a[87] & b[394])^(a[86] & b[395])^(a[85] & b[396])^(a[84] & b[397])^(a[83] & b[398])^(a[82] & b[399])^(a[81] & b[400])^(a[80] & b[401])^(a[79] & b[402])^(a[78] & b[403])^(a[77] & b[404])^(a[76] & b[405])^(a[75] & b[406])^(a[74] & b[407])^(a[73] & b[408]);
assign y[482] = (a[408] & b[74])^(a[407] & b[75])^(a[406] & b[76])^(a[405] & b[77])^(a[404] & b[78])^(a[403] & b[79])^(a[402] & b[80])^(a[401] & b[81])^(a[400] & b[82])^(a[399] & b[83])^(a[398] & b[84])^(a[397] & b[85])^(a[396] & b[86])^(a[395] & b[87])^(a[394] & b[88])^(a[393] & b[89])^(a[392] & b[90])^(a[391] & b[91])^(a[390] & b[92])^(a[389] & b[93])^(a[388] & b[94])^(a[387] & b[95])^(a[386] & b[96])^(a[385] & b[97])^(a[384] & b[98])^(a[383] & b[99])^(a[382] & b[100])^(a[381] & b[101])^(a[380] & b[102])^(a[379] & b[103])^(a[378] & b[104])^(a[377] & b[105])^(a[376] & b[106])^(a[375] & b[107])^(a[374] & b[108])^(a[373] & b[109])^(a[372] & b[110])^(a[371] & b[111])^(a[370] & b[112])^(a[369] & b[113])^(a[368] & b[114])^(a[367] & b[115])^(a[366] & b[116])^(a[365] & b[117])^(a[364] & b[118])^(a[363] & b[119])^(a[362] & b[120])^(a[361] & b[121])^(a[360] & b[122])^(a[359] & b[123])^(a[358] & b[124])^(a[357] & b[125])^(a[356] & b[126])^(a[355] & b[127])^(a[354] & b[128])^(a[353] & b[129])^(a[352] & b[130])^(a[351] & b[131])^(a[350] & b[132])^(a[349] & b[133])^(a[348] & b[134])^(a[347] & b[135])^(a[346] & b[136])^(a[345] & b[137])^(a[344] & b[138])^(a[343] & b[139])^(a[342] & b[140])^(a[341] & b[141])^(a[340] & b[142])^(a[339] & b[143])^(a[338] & b[144])^(a[337] & b[145])^(a[336] & b[146])^(a[335] & b[147])^(a[334] & b[148])^(a[333] & b[149])^(a[332] & b[150])^(a[331] & b[151])^(a[330] & b[152])^(a[329] & b[153])^(a[328] & b[154])^(a[327] & b[155])^(a[326] & b[156])^(a[325] & b[157])^(a[324] & b[158])^(a[323] & b[159])^(a[322] & b[160])^(a[321] & b[161])^(a[320] & b[162])^(a[319] & b[163])^(a[318] & b[164])^(a[317] & b[165])^(a[316] & b[166])^(a[315] & b[167])^(a[314] & b[168])^(a[313] & b[169])^(a[312] & b[170])^(a[311] & b[171])^(a[310] & b[172])^(a[309] & b[173])^(a[308] & b[174])^(a[307] & b[175])^(a[306] & b[176])^(a[305] & b[177])^(a[304] & b[178])^(a[303] & b[179])^(a[302] & b[180])^(a[301] & b[181])^(a[300] & b[182])^(a[299] & b[183])^(a[298] & b[184])^(a[297] & b[185])^(a[296] & b[186])^(a[295] & b[187])^(a[294] & b[188])^(a[293] & b[189])^(a[292] & b[190])^(a[291] & b[191])^(a[290] & b[192])^(a[289] & b[193])^(a[288] & b[194])^(a[287] & b[195])^(a[286] & b[196])^(a[285] & b[197])^(a[284] & b[198])^(a[283] & b[199])^(a[282] & b[200])^(a[281] & b[201])^(a[280] & b[202])^(a[279] & b[203])^(a[278] & b[204])^(a[277] & b[205])^(a[276] & b[206])^(a[275] & b[207])^(a[274] & b[208])^(a[273] & b[209])^(a[272] & b[210])^(a[271] & b[211])^(a[270] & b[212])^(a[269] & b[213])^(a[268] & b[214])^(a[267] & b[215])^(a[266] & b[216])^(a[265] & b[217])^(a[264] & b[218])^(a[263] & b[219])^(a[262] & b[220])^(a[261] & b[221])^(a[260] & b[222])^(a[259] & b[223])^(a[258] & b[224])^(a[257] & b[225])^(a[256] & b[226])^(a[255] & b[227])^(a[254] & b[228])^(a[253] & b[229])^(a[252] & b[230])^(a[251] & b[231])^(a[250] & b[232])^(a[249] & b[233])^(a[248] & b[234])^(a[247] & b[235])^(a[246] & b[236])^(a[245] & b[237])^(a[244] & b[238])^(a[243] & b[239])^(a[242] & b[240])^(a[241] & b[241])^(a[240] & b[242])^(a[239] & b[243])^(a[238] & b[244])^(a[237] & b[245])^(a[236] & b[246])^(a[235] & b[247])^(a[234] & b[248])^(a[233] & b[249])^(a[232] & b[250])^(a[231] & b[251])^(a[230] & b[252])^(a[229] & b[253])^(a[228] & b[254])^(a[227] & b[255])^(a[226] & b[256])^(a[225] & b[257])^(a[224] & b[258])^(a[223] & b[259])^(a[222] & b[260])^(a[221] & b[261])^(a[220] & b[262])^(a[219] & b[263])^(a[218] & b[264])^(a[217] & b[265])^(a[216] & b[266])^(a[215] & b[267])^(a[214] & b[268])^(a[213] & b[269])^(a[212] & b[270])^(a[211] & b[271])^(a[210] & b[272])^(a[209] & b[273])^(a[208] & b[274])^(a[207] & b[275])^(a[206] & b[276])^(a[205] & b[277])^(a[204] & b[278])^(a[203] & b[279])^(a[202] & b[280])^(a[201] & b[281])^(a[200] & b[282])^(a[199] & b[283])^(a[198] & b[284])^(a[197] & b[285])^(a[196] & b[286])^(a[195] & b[287])^(a[194] & b[288])^(a[193] & b[289])^(a[192] & b[290])^(a[191] & b[291])^(a[190] & b[292])^(a[189] & b[293])^(a[188] & b[294])^(a[187] & b[295])^(a[186] & b[296])^(a[185] & b[297])^(a[184] & b[298])^(a[183] & b[299])^(a[182] & b[300])^(a[181] & b[301])^(a[180] & b[302])^(a[179] & b[303])^(a[178] & b[304])^(a[177] & b[305])^(a[176] & b[306])^(a[175] & b[307])^(a[174] & b[308])^(a[173] & b[309])^(a[172] & b[310])^(a[171] & b[311])^(a[170] & b[312])^(a[169] & b[313])^(a[168] & b[314])^(a[167] & b[315])^(a[166] & b[316])^(a[165] & b[317])^(a[164] & b[318])^(a[163] & b[319])^(a[162] & b[320])^(a[161] & b[321])^(a[160] & b[322])^(a[159] & b[323])^(a[158] & b[324])^(a[157] & b[325])^(a[156] & b[326])^(a[155] & b[327])^(a[154] & b[328])^(a[153] & b[329])^(a[152] & b[330])^(a[151] & b[331])^(a[150] & b[332])^(a[149] & b[333])^(a[148] & b[334])^(a[147] & b[335])^(a[146] & b[336])^(a[145] & b[337])^(a[144] & b[338])^(a[143] & b[339])^(a[142] & b[340])^(a[141] & b[341])^(a[140] & b[342])^(a[139] & b[343])^(a[138] & b[344])^(a[137] & b[345])^(a[136] & b[346])^(a[135] & b[347])^(a[134] & b[348])^(a[133] & b[349])^(a[132] & b[350])^(a[131] & b[351])^(a[130] & b[352])^(a[129] & b[353])^(a[128] & b[354])^(a[127] & b[355])^(a[126] & b[356])^(a[125] & b[357])^(a[124] & b[358])^(a[123] & b[359])^(a[122] & b[360])^(a[121] & b[361])^(a[120] & b[362])^(a[119] & b[363])^(a[118] & b[364])^(a[117] & b[365])^(a[116] & b[366])^(a[115] & b[367])^(a[114] & b[368])^(a[113] & b[369])^(a[112] & b[370])^(a[111] & b[371])^(a[110] & b[372])^(a[109] & b[373])^(a[108] & b[374])^(a[107] & b[375])^(a[106] & b[376])^(a[105] & b[377])^(a[104] & b[378])^(a[103] & b[379])^(a[102] & b[380])^(a[101] & b[381])^(a[100] & b[382])^(a[99] & b[383])^(a[98] & b[384])^(a[97] & b[385])^(a[96] & b[386])^(a[95] & b[387])^(a[94] & b[388])^(a[93] & b[389])^(a[92] & b[390])^(a[91] & b[391])^(a[90] & b[392])^(a[89] & b[393])^(a[88] & b[394])^(a[87] & b[395])^(a[86] & b[396])^(a[85] & b[397])^(a[84] & b[398])^(a[83] & b[399])^(a[82] & b[400])^(a[81] & b[401])^(a[80] & b[402])^(a[79] & b[403])^(a[78] & b[404])^(a[77] & b[405])^(a[76] & b[406])^(a[75] & b[407])^(a[74] & b[408]);
assign y[483] = (a[408] & b[75])^(a[407] & b[76])^(a[406] & b[77])^(a[405] & b[78])^(a[404] & b[79])^(a[403] & b[80])^(a[402] & b[81])^(a[401] & b[82])^(a[400] & b[83])^(a[399] & b[84])^(a[398] & b[85])^(a[397] & b[86])^(a[396] & b[87])^(a[395] & b[88])^(a[394] & b[89])^(a[393] & b[90])^(a[392] & b[91])^(a[391] & b[92])^(a[390] & b[93])^(a[389] & b[94])^(a[388] & b[95])^(a[387] & b[96])^(a[386] & b[97])^(a[385] & b[98])^(a[384] & b[99])^(a[383] & b[100])^(a[382] & b[101])^(a[381] & b[102])^(a[380] & b[103])^(a[379] & b[104])^(a[378] & b[105])^(a[377] & b[106])^(a[376] & b[107])^(a[375] & b[108])^(a[374] & b[109])^(a[373] & b[110])^(a[372] & b[111])^(a[371] & b[112])^(a[370] & b[113])^(a[369] & b[114])^(a[368] & b[115])^(a[367] & b[116])^(a[366] & b[117])^(a[365] & b[118])^(a[364] & b[119])^(a[363] & b[120])^(a[362] & b[121])^(a[361] & b[122])^(a[360] & b[123])^(a[359] & b[124])^(a[358] & b[125])^(a[357] & b[126])^(a[356] & b[127])^(a[355] & b[128])^(a[354] & b[129])^(a[353] & b[130])^(a[352] & b[131])^(a[351] & b[132])^(a[350] & b[133])^(a[349] & b[134])^(a[348] & b[135])^(a[347] & b[136])^(a[346] & b[137])^(a[345] & b[138])^(a[344] & b[139])^(a[343] & b[140])^(a[342] & b[141])^(a[341] & b[142])^(a[340] & b[143])^(a[339] & b[144])^(a[338] & b[145])^(a[337] & b[146])^(a[336] & b[147])^(a[335] & b[148])^(a[334] & b[149])^(a[333] & b[150])^(a[332] & b[151])^(a[331] & b[152])^(a[330] & b[153])^(a[329] & b[154])^(a[328] & b[155])^(a[327] & b[156])^(a[326] & b[157])^(a[325] & b[158])^(a[324] & b[159])^(a[323] & b[160])^(a[322] & b[161])^(a[321] & b[162])^(a[320] & b[163])^(a[319] & b[164])^(a[318] & b[165])^(a[317] & b[166])^(a[316] & b[167])^(a[315] & b[168])^(a[314] & b[169])^(a[313] & b[170])^(a[312] & b[171])^(a[311] & b[172])^(a[310] & b[173])^(a[309] & b[174])^(a[308] & b[175])^(a[307] & b[176])^(a[306] & b[177])^(a[305] & b[178])^(a[304] & b[179])^(a[303] & b[180])^(a[302] & b[181])^(a[301] & b[182])^(a[300] & b[183])^(a[299] & b[184])^(a[298] & b[185])^(a[297] & b[186])^(a[296] & b[187])^(a[295] & b[188])^(a[294] & b[189])^(a[293] & b[190])^(a[292] & b[191])^(a[291] & b[192])^(a[290] & b[193])^(a[289] & b[194])^(a[288] & b[195])^(a[287] & b[196])^(a[286] & b[197])^(a[285] & b[198])^(a[284] & b[199])^(a[283] & b[200])^(a[282] & b[201])^(a[281] & b[202])^(a[280] & b[203])^(a[279] & b[204])^(a[278] & b[205])^(a[277] & b[206])^(a[276] & b[207])^(a[275] & b[208])^(a[274] & b[209])^(a[273] & b[210])^(a[272] & b[211])^(a[271] & b[212])^(a[270] & b[213])^(a[269] & b[214])^(a[268] & b[215])^(a[267] & b[216])^(a[266] & b[217])^(a[265] & b[218])^(a[264] & b[219])^(a[263] & b[220])^(a[262] & b[221])^(a[261] & b[222])^(a[260] & b[223])^(a[259] & b[224])^(a[258] & b[225])^(a[257] & b[226])^(a[256] & b[227])^(a[255] & b[228])^(a[254] & b[229])^(a[253] & b[230])^(a[252] & b[231])^(a[251] & b[232])^(a[250] & b[233])^(a[249] & b[234])^(a[248] & b[235])^(a[247] & b[236])^(a[246] & b[237])^(a[245] & b[238])^(a[244] & b[239])^(a[243] & b[240])^(a[242] & b[241])^(a[241] & b[242])^(a[240] & b[243])^(a[239] & b[244])^(a[238] & b[245])^(a[237] & b[246])^(a[236] & b[247])^(a[235] & b[248])^(a[234] & b[249])^(a[233] & b[250])^(a[232] & b[251])^(a[231] & b[252])^(a[230] & b[253])^(a[229] & b[254])^(a[228] & b[255])^(a[227] & b[256])^(a[226] & b[257])^(a[225] & b[258])^(a[224] & b[259])^(a[223] & b[260])^(a[222] & b[261])^(a[221] & b[262])^(a[220] & b[263])^(a[219] & b[264])^(a[218] & b[265])^(a[217] & b[266])^(a[216] & b[267])^(a[215] & b[268])^(a[214] & b[269])^(a[213] & b[270])^(a[212] & b[271])^(a[211] & b[272])^(a[210] & b[273])^(a[209] & b[274])^(a[208] & b[275])^(a[207] & b[276])^(a[206] & b[277])^(a[205] & b[278])^(a[204] & b[279])^(a[203] & b[280])^(a[202] & b[281])^(a[201] & b[282])^(a[200] & b[283])^(a[199] & b[284])^(a[198] & b[285])^(a[197] & b[286])^(a[196] & b[287])^(a[195] & b[288])^(a[194] & b[289])^(a[193] & b[290])^(a[192] & b[291])^(a[191] & b[292])^(a[190] & b[293])^(a[189] & b[294])^(a[188] & b[295])^(a[187] & b[296])^(a[186] & b[297])^(a[185] & b[298])^(a[184] & b[299])^(a[183] & b[300])^(a[182] & b[301])^(a[181] & b[302])^(a[180] & b[303])^(a[179] & b[304])^(a[178] & b[305])^(a[177] & b[306])^(a[176] & b[307])^(a[175] & b[308])^(a[174] & b[309])^(a[173] & b[310])^(a[172] & b[311])^(a[171] & b[312])^(a[170] & b[313])^(a[169] & b[314])^(a[168] & b[315])^(a[167] & b[316])^(a[166] & b[317])^(a[165] & b[318])^(a[164] & b[319])^(a[163] & b[320])^(a[162] & b[321])^(a[161] & b[322])^(a[160] & b[323])^(a[159] & b[324])^(a[158] & b[325])^(a[157] & b[326])^(a[156] & b[327])^(a[155] & b[328])^(a[154] & b[329])^(a[153] & b[330])^(a[152] & b[331])^(a[151] & b[332])^(a[150] & b[333])^(a[149] & b[334])^(a[148] & b[335])^(a[147] & b[336])^(a[146] & b[337])^(a[145] & b[338])^(a[144] & b[339])^(a[143] & b[340])^(a[142] & b[341])^(a[141] & b[342])^(a[140] & b[343])^(a[139] & b[344])^(a[138] & b[345])^(a[137] & b[346])^(a[136] & b[347])^(a[135] & b[348])^(a[134] & b[349])^(a[133] & b[350])^(a[132] & b[351])^(a[131] & b[352])^(a[130] & b[353])^(a[129] & b[354])^(a[128] & b[355])^(a[127] & b[356])^(a[126] & b[357])^(a[125] & b[358])^(a[124] & b[359])^(a[123] & b[360])^(a[122] & b[361])^(a[121] & b[362])^(a[120] & b[363])^(a[119] & b[364])^(a[118] & b[365])^(a[117] & b[366])^(a[116] & b[367])^(a[115] & b[368])^(a[114] & b[369])^(a[113] & b[370])^(a[112] & b[371])^(a[111] & b[372])^(a[110] & b[373])^(a[109] & b[374])^(a[108] & b[375])^(a[107] & b[376])^(a[106] & b[377])^(a[105] & b[378])^(a[104] & b[379])^(a[103] & b[380])^(a[102] & b[381])^(a[101] & b[382])^(a[100] & b[383])^(a[99] & b[384])^(a[98] & b[385])^(a[97] & b[386])^(a[96] & b[387])^(a[95] & b[388])^(a[94] & b[389])^(a[93] & b[390])^(a[92] & b[391])^(a[91] & b[392])^(a[90] & b[393])^(a[89] & b[394])^(a[88] & b[395])^(a[87] & b[396])^(a[86] & b[397])^(a[85] & b[398])^(a[84] & b[399])^(a[83] & b[400])^(a[82] & b[401])^(a[81] & b[402])^(a[80] & b[403])^(a[79] & b[404])^(a[78] & b[405])^(a[77] & b[406])^(a[76] & b[407])^(a[75] & b[408]);
assign y[484] = (a[408] & b[76])^(a[407] & b[77])^(a[406] & b[78])^(a[405] & b[79])^(a[404] & b[80])^(a[403] & b[81])^(a[402] & b[82])^(a[401] & b[83])^(a[400] & b[84])^(a[399] & b[85])^(a[398] & b[86])^(a[397] & b[87])^(a[396] & b[88])^(a[395] & b[89])^(a[394] & b[90])^(a[393] & b[91])^(a[392] & b[92])^(a[391] & b[93])^(a[390] & b[94])^(a[389] & b[95])^(a[388] & b[96])^(a[387] & b[97])^(a[386] & b[98])^(a[385] & b[99])^(a[384] & b[100])^(a[383] & b[101])^(a[382] & b[102])^(a[381] & b[103])^(a[380] & b[104])^(a[379] & b[105])^(a[378] & b[106])^(a[377] & b[107])^(a[376] & b[108])^(a[375] & b[109])^(a[374] & b[110])^(a[373] & b[111])^(a[372] & b[112])^(a[371] & b[113])^(a[370] & b[114])^(a[369] & b[115])^(a[368] & b[116])^(a[367] & b[117])^(a[366] & b[118])^(a[365] & b[119])^(a[364] & b[120])^(a[363] & b[121])^(a[362] & b[122])^(a[361] & b[123])^(a[360] & b[124])^(a[359] & b[125])^(a[358] & b[126])^(a[357] & b[127])^(a[356] & b[128])^(a[355] & b[129])^(a[354] & b[130])^(a[353] & b[131])^(a[352] & b[132])^(a[351] & b[133])^(a[350] & b[134])^(a[349] & b[135])^(a[348] & b[136])^(a[347] & b[137])^(a[346] & b[138])^(a[345] & b[139])^(a[344] & b[140])^(a[343] & b[141])^(a[342] & b[142])^(a[341] & b[143])^(a[340] & b[144])^(a[339] & b[145])^(a[338] & b[146])^(a[337] & b[147])^(a[336] & b[148])^(a[335] & b[149])^(a[334] & b[150])^(a[333] & b[151])^(a[332] & b[152])^(a[331] & b[153])^(a[330] & b[154])^(a[329] & b[155])^(a[328] & b[156])^(a[327] & b[157])^(a[326] & b[158])^(a[325] & b[159])^(a[324] & b[160])^(a[323] & b[161])^(a[322] & b[162])^(a[321] & b[163])^(a[320] & b[164])^(a[319] & b[165])^(a[318] & b[166])^(a[317] & b[167])^(a[316] & b[168])^(a[315] & b[169])^(a[314] & b[170])^(a[313] & b[171])^(a[312] & b[172])^(a[311] & b[173])^(a[310] & b[174])^(a[309] & b[175])^(a[308] & b[176])^(a[307] & b[177])^(a[306] & b[178])^(a[305] & b[179])^(a[304] & b[180])^(a[303] & b[181])^(a[302] & b[182])^(a[301] & b[183])^(a[300] & b[184])^(a[299] & b[185])^(a[298] & b[186])^(a[297] & b[187])^(a[296] & b[188])^(a[295] & b[189])^(a[294] & b[190])^(a[293] & b[191])^(a[292] & b[192])^(a[291] & b[193])^(a[290] & b[194])^(a[289] & b[195])^(a[288] & b[196])^(a[287] & b[197])^(a[286] & b[198])^(a[285] & b[199])^(a[284] & b[200])^(a[283] & b[201])^(a[282] & b[202])^(a[281] & b[203])^(a[280] & b[204])^(a[279] & b[205])^(a[278] & b[206])^(a[277] & b[207])^(a[276] & b[208])^(a[275] & b[209])^(a[274] & b[210])^(a[273] & b[211])^(a[272] & b[212])^(a[271] & b[213])^(a[270] & b[214])^(a[269] & b[215])^(a[268] & b[216])^(a[267] & b[217])^(a[266] & b[218])^(a[265] & b[219])^(a[264] & b[220])^(a[263] & b[221])^(a[262] & b[222])^(a[261] & b[223])^(a[260] & b[224])^(a[259] & b[225])^(a[258] & b[226])^(a[257] & b[227])^(a[256] & b[228])^(a[255] & b[229])^(a[254] & b[230])^(a[253] & b[231])^(a[252] & b[232])^(a[251] & b[233])^(a[250] & b[234])^(a[249] & b[235])^(a[248] & b[236])^(a[247] & b[237])^(a[246] & b[238])^(a[245] & b[239])^(a[244] & b[240])^(a[243] & b[241])^(a[242] & b[242])^(a[241] & b[243])^(a[240] & b[244])^(a[239] & b[245])^(a[238] & b[246])^(a[237] & b[247])^(a[236] & b[248])^(a[235] & b[249])^(a[234] & b[250])^(a[233] & b[251])^(a[232] & b[252])^(a[231] & b[253])^(a[230] & b[254])^(a[229] & b[255])^(a[228] & b[256])^(a[227] & b[257])^(a[226] & b[258])^(a[225] & b[259])^(a[224] & b[260])^(a[223] & b[261])^(a[222] & b[262])^(a[221] & b[263])^(a[220] & b[264])^(a[219] & b[265])^(a[218] & b[266])^(a[217] & b[267])^(a[216] & b[268])^(a[215] & b[269])^(a[214] & b[270])^(a[213] & b[271])^(a[212] & b[272])^(a[211] & b[273])^(a[210] & b[274])^(a[209] & b[275])^(a[208] & b[276])^(a[207] & b[277])^(a[206] & b[278])^(a[205] & b[279])^(a[204] & b[280])^(a[203] & b[281])^(a[202] & b[282])^(a[201] & b[283])^(a[200] & b[284])^(a[199] & b[285])^(a[198] & b[286])^(a[197] & b[287])^(a[196] & b[288])^(a[195] & b[289])^(a[194] & b[290])^(a[193] & b[291])^(a[192] & b[292])^(a[191] & b[293])^(a[190] & b[294])^(a[189] & b[295])^(a[188] & b[296])^(a[187] & b[297])^(a[186] & b[298])^(a[185] & b[299])^(a[184] & b[300])^(a[183] & b[301])^(a[182] & b[302])^(a[181] & b[303])^(a[180] & b[304])^(a[179] & b[305])^(a[178] & b[306])^(a[177] & b[307])^(a[176] & b[308])^(a[175] & b[309])^(a[174] & b[310])^(a[173] & b[311])^(a[172] & b[312])^(a[171] & b[313])^(a[170] & b[314])^(a[169] & b[315])^(a[168] & b[316])^(a[167] & b[317])^(a[166] & b[318])^(a[165] & b[319])^(a[164] & b[320])^(a[163] & b[321])^(a[162] & b[322])^(a[161] & b[323])^(a[160] & b[324])^(a[159] & b[325])^(a[158] & b[326])^(a[157] & b[327])^(a[156] & b[328])^(a[155] & b[329])^(a[154] & b[330])^(a[153] & b[331])^(a[152] & b[332])^(a[151] & b[333])^(a[150] & b[334])^(a[149] & b[335])^(a[148] & b[336])^(a[147] & b[337])^(a[146] & b[338])^(a[145] & b[339])^(a[144] & b[340])^(a[143] & b[341])^(a[142] & b[342])^(a[141] & b[343])^(a[140] & b[344])^(a[139] & b[345])^(a[138] & b[346])^(a[137] & b[347])^(a[136] & b[348])^(a[135] & b[349])^(a[134] & b[350])^(a[133] & b[351])^(a[132] & b[352])^(a[131] & b[353])^(a[130] & b[354])^(a[129] & b[355])^(a[128] & b[356])^(a[127] & b[357])^(a[126] & b[358])^(a[125] & b[359])^(a[124] & b[360])^(a[123] & b[361])^(a[122] & b[362])^(a[121] & b[363])^(a[120] & b[364])^(a[119] & b[365])^(a[118] & b[366])^(a[117] & b[367])^(a[116] & b[368])^(a[115] & b[369])^(a[114] & b[370])^(a[113] & b[371])^(a[112] & b[372])^(a[111] & b[373])^(a[110] & b[374])^(a[109] & b[375])^(a[108] & b[376])^(a[107] & b[377])^(a[106] & b[378])^(a[105] & b[379])^(a[104] & b[380])^(a[103] & b[381])^(a[102] & b[382])^(a[101] & b[383])^(a[100] & b[384])^(a[99] & b[385])^(a[98] & b[386])^(a[97] & b[387])^(a[96] & b[388])^(a[95] & b[389])^(a[94] & b[390])^(a[93] & b[391])^(a[92] & b[392])^(a[91] & b[393])^(a[90] & b[394])^(a[89] & b[395])^(a[88] & b[396])^(a[87] & b[397])^(a[86] & b[398])^(a[85] & b[399])^(a[84] & b[400])^(a[83] & b[401])^(a[82] & b[402])^(a[81] & b[403])^(a[80] & b[404])^(a[79] & b[405])^(a[78] & b[406])^(a[77] & b[407])^(a[76] & b[408]);
assign y[485] = (a[408] & b[77])^(a[407] & b[78])^(a[406] & b[79])^(a[405] & b[80])^(a[404] & b[81])^(a[403] & b[82])^(a[402] & b[83])^(a[401] & b[84])^(a[400] & b[85])^(a[399] & b[86])^(a[398] & b[87])^(a[397] & b[88])^(a[396] & b[89])^(a[395] & b[90])^(a[394] & b[91])^(a[393] & b[92])^(a[392] & b[93])^(a[391] & b[94])^(a[390] & b[95])^(a[389] & b[96])^(a[388] & b[97])^(a[387] & b[98])^(a[386] & b[99])^(a[385] & b[100])^(a[384] & b[101])^(a[383] & b[102])^(a[382] & b[103])^(a[381] & b[104])^(a[380] & b[105])^(a[379] & b[106])^(a[378] & b[107])^(a[377] & b[108])^(a[376] & b[109])^(a[375] & b[110])^(a[374] & b[111])^(a[373] & b[112])^(a[372] & b[113])^(a[371] & b[114])^(a[370] & b[115])^(a[369] & b[116])^(a[368] & b[117])^(a[367] & b[118])^(a[366] & b[119])^(a[365] & b[120])^(a[364] & b[121])^(a[363] & b[122])^(a[362] & b[123])^(a[361] & b[124])^(a[360] & b[125])^(a[359] & b[126])^(a[358] & b[127])^(a[357] & b[128])^(a[356] & b[129])^(a[355] & b[130])^(a[354] & b[131])^(a[353] & b[132])^(a[352] & b[133])^(a[351] & b[134])^(a[350] & b[135])^(a[349] & b[136])^(a[348] & b[137])^(a[347] & b[138])^(a[346] & b[139])^(a[345] & b[140])^(a[344] & b[141])^(a[343] & b[142])^(a[342] & b[143])^(a[341] & b[144])^(a[340] & b[145])^(a[339] & b[146])^(a[338] & b[147])^(a[337] & b[148])^(a[336] & b[149])^(a[335] & b[150])^(a[334] & b[151])^(a[333] & b[152])^(a[332] & b[153])^(a[331] & b[154])^(a[330] & b[155])^(a[329] & b[156])^(a[328] & b[157])^(a[327] & b[158])^(a[326] & b[159])^(a[325] & b[160])^(a[324] & b[161])^(a[323] & b[162])^(a[322] & b[163])^(a[321] & b[164])^(a[320] & b[165])^(a[319] & b[166])^(a[318] & b[167])^(a[317] & b[168])^(a[316] & b[169])^(a[315] & b[170])^(a[314] & b[171])^(a[313] & b[172])^(a[312] & b[173])^(a[311] & b[174])^(a[310] & b[175])^(a[309] & b[176])^(a[308] & b[177])^(a[307] & b[178])^(a[306] & b[179])^(a[305] & b[180])^(a[304] & b[181])^(a[303] & b[182])^(a[302] & b[183])^(a[301] & b[184])^(a[300] & b[185])^(a[299] & b[186])^(a[298] & b[187])^(a[297] & b[188])^(a[296] & b[189])^(a[295] & b[190])^(a[294] & b[191])^(a[293] & b[192])^(a[292] & b[193])^(a[291] & b[194])^(a[290] & b[195])^(a[289] & b[196])^(a[288] & b[197])^(a[287] & b[198])^(a[286] & b[199])^(a[285] & b[200])^(a[284] & b[201])^(a[283] & b[202])^(a[282] & b[203])^(a[281] & b[204])^(a[280] & b[205])^(a[279] & b[206])^(a[278] & b[207])^(a[277] & b[208])^(a[276] & b[209])^(a[275] & b[210])^(a[274] & b[211])^(a[273] & b[212])^(a[272] & b[213])^(a[271] & b[214])^(a[270] & b[215])^(a[269] & b[216])^(a[268] & b[217])^(a[267] & b[218])^(a[266] & b[219])^(a[265] & b[220])^(a[264] & b[221])^(a[263] & b[222])^(a[262] & b[223])^(a[261] & b[224])^(a[260] & b[225])^(a[259] & b[226])^(a[258] & b[227])^(a[257] & b[228])^(a[256] & b[229])^(a[255] & b[230])^(a[254] & b[231])^(a[253] & b[232])^(a[252] & b[233])^(a[251] & b[234])^(a[250] & b[235])^(a[249] & b[236])^(a[248] & b[237])^(a[247] & b[238])^(a[246] & b[239])^(a[245] & b[240])^(a[244] & b[241])^(a[243] & b[242])^(a[242] & b[243])^(a[241] & b[244])^(a[240] & b[245])^(a[239] & b[246])^(a[238] & b[247])^(a[237] & b[248])^(a[236] & b[249])^(a[235] & b[250])^(a[234] & b[251])^(a[233] & b[252])^(a[232] & b[253])^(a[231] & b[254])^(a[230] & b[255])^(a[229] & b[256])^(a[228] & b[257])^(a[227] & b[258])^(a[226] & b[259])^(a[225] & b[260])^(a[224] & b[261])^(a[223] & b[262])^(a[222] & b[263])^(a[221] & b[264])^(a[220] & b[265])^(a[219] & b[266])^(a[218] & b[267])^(a[217] & b[268])^(a[216] & b[269])^(a[215] & b[270])^(a[214] & b[271])^(a[213] & b[272])^(a[212] & b[273])^(a[211] & b[274])^(a[210] & b[275])^(a[209] & b[276])^(a[208] & b[277])^(a[207] & b[278])^(a[206] & b[279])^(a[205] & b[280])^(a[204] & b[281])^(a[203] & b[282])^(a[202] & b[283])^(a[201] & b[284])^(a[200] & b[285])^(a[199] & b[286])^(a[198] & b[287])^(a[197] & b[288])^(a[196] & b[289])^(a[195] & b[290])^(a[194] & b[291])^(a[193] & b[292])^(a[192] & b[293])^(a[191] & b[294])^(a[190] & b[295])^(a[189] & b[296])^(a[188] & b[297])^(a[187] & b[298])^(a[186] & b[299])^(a[185] & b[300])^(a[184] & b[301])^(a[183] & b[302])^(a[182] & b[303])^(a[181] & b[304])^(a[180] & b[305])^(a[179] & b[306])^(a[178] & b[307])^(a[177] & b[308])^(a[176] & b[309])^(a[175] & b[310])^(a[174] & b[311])^(a[173] & b[312])^(a[172] & b[313])^(a[171] & b[314])^(a[170] & b[315])^(a[169] & b[316])^(a[168] & b[317])^(a[167] & b[318])^(a[166] & b[319])^(a[165] & b[320])^(a[164] & b[321])^(a[163] & b[322])^(a[162] & b[323])^(a[161] & b[324])^(a[160] & b[325])^(a[159] & b[326])^(a[158] & b[327])^(a[157] & b[328])^(a[156] & b[329])^(a[155] & b[330])^(a[154] & b[331])^(a[153] & b[332])^(a[152] & b[333])^(a[151] & b[334])^(a[150] & b[335])^(a[149] & b[336])^(a[148] & b[337])^(a[147] & b[338])^(a[146] & b[339])^(a[145] & b[340])^(a[144] & b[341])^(a[143] & b[342])^(a[142] & b[343])^(a[141] & b[344])^(a[140] & b[345])^(a[139] & b[346])^(a[138] & b[347])^(a[137] & b[348])^(a[136] & b[349])^(a[135] & b[350])^(a[134] & b[351])^(a[133] & b[352])^(a[132] & b[353])^(a[131] & b[354])^(a[130] & b[355])^(a[129] & b[356])^(a[128] & b[357])^(a[127] & b[358])^(a[126] & b[359])^(a[125] & b[360])^(a[124] & b[361])^(a[123] & b[362])^(a[122] & b[363])^(a[121] & b[364])^(a[120] & b[365])^(a[119] & b[366])^(a[118] & b[367])^(a[117] & b[368])^(a[116] & b[369])^(a[115] & b[370])^(a[114] & b[371])^(a[113] & b[372])^(a[112] & b[373])^(a[111] & b[374])^(a[110] & b[375])^(a[109] & b[376])^(a[108] & b[377])^(a[107] & b[378])^(a[106] & b[379])^(a[105] & b[380])^(a[104] & b[381])^(a[103] & b[382])^(a[102] & b[383])^(a[101] & b[384])^(a[100] & b[385])^(a[99] & b[386])^(a[98] & b[387])^(a[97] & b[388])^(a[96] & b[389])^(a[95] & b[390])^(a[94] & b[391])^(a[93] & b[392])^(a[92] & b[393])^(a[91] & b[394])^(a[90] & b[395])^(a[89] & b[396])^(a[88] & b[397])^(a[87] & b[398])^(a[86] & b[399])^(a[85] & b[400])^(a[84] & b[401])^(a[83] & b[402])^(a[82] & b[403])^(a[81] & b[404])^(a[80] & b[405])^(a[79] & b[406])^(a[78] & b[407])^(a[77] & b[408]);
assign y[486] = (a[408] & b[78])^(a[407] & b[79])^(a[406] & b[80])^(a[405] & b[81])^(a[404] & b[82])^(a[403] & b[83])^(a[402] & b[84])^(a[401] & b[85])^(a[400] & b[86])^(a[399] & b[87])^(a[398] & b[88])^(a[397] & b[89])^(a[396] & b[90])^(a[395] & b[91])^(a[394] & b[92])^(a[393] & b[93])^(a[392] & b[94])^(a[391] & b[95])^(a[390] & b[96])^(a[389] & b[97])^(a[388] & b[98])^(a[387] & b[99])^(a[386] & b[100])^(a[385] & b[101])^(a[384] & b[102])^(a[383] & b[103])^(a[382] & b[104])^(a[381] & b[105])^(a[380] & b[106])^(a[379] & b[107])^(a[378] & b[108])^(a[377] & b[109])^(a[376] & b[110])^(a[375] & b[111])^(a[374] & b[112])^(a[373] & b[113])^(a[372] & b[114])^(a[371] & b[115])^(a[370] & b[116])^(a[369] & b[117])^(a[368] & b[118])^(a[367] & b[119])^(a[366] & b[120])^(a[365] & b[121])^(a[364] & b[122])^(a[363] & b[123])^(a[362] & b[124])^(a[361] & b[125])^(a[360] & b[126])^(a[359] & b[127])^(a[358] & b[128])^(a[357] & b[129])^(a[356] & b[130])^(a[355] & b[131])^(a[354] & b[132])^(a[353] & b[133])^(a[352] & b[134])^(a[351] & b[135])^(a[350] & b[136])^(a[349] & b[137])^(a[348] & b[138])^(a[347] & b[139])^(a[346] & b[140])^(a[345] & b[141])^(a[344] & b[142])^(a[343] & b[143])^(a[342] & b[144])^(a[341] & b[145])^(a[340] & b[146])^(a[339] & b[147])^(a[338] & b[148])^(a[337] & b[149])^(a[336] & b[150])^(a[335] & b[151])^(a[334] & b[152])^(a[333] & b[153])^(a[332] & b[154])^(a[331] & b[155])^(a[330] & b[156])^(a[329] & b[157])^(a[328] & b[158])^(a[327] & b[159])^(a[326] & b[160])^(a[325] & b[161])^(a[324] & b[162])^(a[323] & b[163])^(a[322] & b[164])^(a[321] & b[165])^(a[320] & b[166])^(a[319] & b[167])^(a[318] & b[168])^(a[317] & b[169])^(a[316] & b[170])^(a[315] & b[171])^(a[314] & b[172])^(a[313] & b[173])^(a[312] & b[174])^(a[311] & b[175])^(a[310] & b[176])^(a[309] & b[177])^(a[308] & b[178])^(a[307] & b[179])^(a[306] & b[180])^(a[305] & b[181])^(a[304] & b[182])^(a[303] & b[183])^(a[302] & b[184])^(a[301] & b[185])^(a[300] & b[186])^(a[299] & b[187])^(a[298] & b[188])^(a[297] & b[189])^(a[296] & b[190])^(a[295] & b[191])^(a[294] & b[192])^(a[293] & b[193])^(a[292] & b[194])^(a[291] & b[195])^(a[290] & b[196])^(a[289] & b[197])^(a[288] & b[198])^(a[287] & b[199])^(a[286] & b[200])^(a[285] & b[201])^(a[284] & b[202])^(a[283] & b[203])^(a[282] & b[204])^(a[281] & b[205])^(a[280] & b[206])^(a[279] & b[207])^(a[278] & b[208])^(a[277] & b[209])^(a[276] & b[210])^(a[275] & b[211])^(a[274] & b[212])^(a[273] & b[213])^(a[272] & b[214])^(a[271] & b[215])^(a[270] & b[216])^(a[269] & b[217])^(a[268] & b[218])^(a[267] & b[219])^(a[266] & b[220])^(a[265] & b[221])^(a[264] & b[222])^(a[263] & b[223])^(a[262] & b[224])^(a[261] & b[225])^(a[260] & b[226])^(a[259] & b[227])^(a[258] & b[228])^(a[257] & b[229])^(a[256] & b[230])^(a[255] & b[231])^(a[254] & b[232])^(a[253] & b[233])^(a[252] & b[234])^(a[251] & b[235])^(a[250] & b[236])^(a[249] & b[237])^(a[248] & b[238])^(a[247] & b[239])^(a[246] & b[240])^(a[245] & b[241])^(a[244] & b[242])^(a[243] & b[243])^(a[242] & b[244])^(a[241] & b[245])^(a[240] & b[246])^(a[239] & b[247])^(a[238] & b[248])^(a[237] & b[249])^(a[236] & b[250])^(a[235] & b[251])^(a[234] & b[252])^(a[233] & b[253])^(a[232] & b[254])^(a[231] & b[255])^(a[230] & b[256])^(a[229] & b[257])^(a[228] & b[258])^(a[227] & b[259])^(a[226] & b[260])^(a[225] & b[261])^(a[224] & b[262])^(a[223] & b[263])^(a[222] & b[264])^(a[221] & b[265])^(a[220] & b[266])^(a[219] & b[267])^(a[218] & b[268])^(a[217] & b[269])^(a[216] & b[270])^(a[215] & b[271])^(a[214] & b[272])^(a[213] & b[273])^(a[212] & b[274])^(a[211] & b[275])^(a[210] & b[276])^(a[209] & b[277])^(a[208] & b[278])^(a[207] & b[279])^(a[206] & b[280])^(a[205] & b[281])^(a[204] & b[282])^(a[203] & b[283])^(a[202] & b[284])^(a[201] & b[285])^(a[200] & b[286])^(a[199] & b[287])^(a[198] & b[288])^(a[197] & b[289])^(a[196] & b[290])^(a[195] & b[291])^(a[194] & b[292])^(a[193] & b[293])^(a[192] & b[294])^(a[191] & b[295])^(a[190] & b[296])^(a[189] & b[297])^(a[188] & b[298])^(a[187] & b[299])^(a[186] & b[300])^(a[185] & b[301])^(a[184] & b[302])^(a[183] & b[303])^(a[182] & b[304])^(a[181] & b[305])^(a[180] & b[306])^(a[179] & b[307])^(a[178] & b[308])^(a[177] & b[309])^(a[176] & b[310])^(a[175] & b[311])^(a[174] & b[312])^(a[173] & b[313])^(a[172] & b[314])^(a[171] & b[315])^(a[170] & b[316])^(a[169] & b[317])^(a[168] & b[318])^(a[167] & b[319])^(a[166] & b[320])^(a[165] & b[321])^(a[164] & b[322])^(a[163] & b[323])^(a[162] & b[324])^(a[161] & b[325])^(a[160] & b[326])^(a[159] & b[327])^(a[158] & b[328])^(a[157] & b[329])^(a[156] & b[330])^(a[155] & b[331])^(a[154] & b[332])^(a[153] & b[333])^(a[152] & b[334])^(a[151] & b[335])^(a[150] & b[336])^(a[149] & b[337])^(a[148] & b[338])^(a[147] & b[339])^(a[146] & b[340])^(a[145] & b[341])^(a[144] & b[342])^(a[143] & b[343])^(a[142] & b[344])^(a[141] & b[345])^(a[140] & b[346])^(a[139] & b[347])^(a[138] & b[348])^(a[137] & b[349])^(a[136] & b[350])^(a[135] & b[351])^(a[134] & b[352])^(a[133] & b[353])^(a[132] & b[354])^(a[131] & b[355])^(a[130] & b[356])^(a[129] & b[357])^(a[128] & b[358])^(a[127] & b[359])^(a[126] & b[360])^(a[125] & b[361])^(a[124] & b[362])^(a[123] & b[363])^(a[122] & b[364])^(a[121] & b[365])^(a[120] & b[366])^(a[119] & b[367])^(a[118] & b[368])^(a[117] & b[369])^(a[116] & b[370])^(a[115] & b[371])^(a[114] & b[372])^(a[113] & b[373])^(a[112] & b[374])^(a[111] & b[375])^(a[110] & b[376])^(a[109] & b[377])^(a[108] & b[378])^(a[107] & b[379])^(a[106] & b[380])^(a[105] & b[381])^(a[104] & b[382])^(a[103] & b[383])^(a[102] & b[384])^(a[101] & b[385])^(a[100] & b[386])^(a[99] & b[387])^(a[98] & b[388])^(a[97] & b[389])^(a[96] & b[390])^(a[95] & b[391])^(a[94] & b[392])^(a[93] & b[393])^(a[92] & b[394])^(a[91] & b[395])^(a[90] & b[396])^(a[89] & b[397])^(a[88] & b[398])^(a[87] & b[399])^(a[86] & b[400])^(a[85] & b[401])^(a[84] & b[402])^(a[83] & b[403])^(a[82] & b[404])^(a[81] & b[405])^(a[80] & b[406])^(a[79] & b[407])^(a[78] & b[408]);
assign y[487] = (a[408] & b[79])^(a[407] & b[80])^(a[406] & b[81])^(a[405] & b[82])^(a[404] & b[83])^(a[403] & b[84])^(a[402] & b[85])^(a[401] & b[86])^(a[400] & b[87])^(a[399] & b[88])^(a[398] & b[89])^(a[397] & b[90])^(a[396] & b[91])^(a[395] & b[92])^(a[394] & b[93])^(a[393] & b[94])^(a[392] & b[95])^(a[391] & b[96])^(a[390] & b[97])^(a[389] & b[98])^(a[388] & b[99])^(a[387] & b[100])^(a[386] & b[101])^(a[385] & b[102])^(a[384] & b[103])^(a[383] & b[104])^(a[382] & b[105])^(a[381] & b[106])^(a[380] & b[107])^(a[379] & b[108])^(a[378] & b[109])^(a[377] & b[110])^(a[376] & b[111])^(a[375] & b[112])^(a[374] & b[113])^(a[373] & b[114])^(a[372] & b[115])^(a[371] & b[116])^(a[370] & b[117])^(a[369] & b[118])^(a[368] & b[119])^(a[367] & b[120])^(a[366] & b[121])^(a[365] & b[122])^(a[364] & b[123])^(a[363] & b[124])^(a[362] & b[125])^(a[361] & b[126])^(a[360] & b[127])^(a[359] & b[128])^(a[358] & b[129])^(a[357] & b[130])^(a[356] & b[131])^(a[355] & b[132])^(a[354] & b[133])^(a[353] & b[134])^(a[352] & b[135])^(a[351] & b[136])^(a[350] & b[137])^(a[349] & b[138])^(a[348] & b[139])^(a[347] & b[140])^(a[346] & b[141])^(a[345] & b[142])^(a[344] & b[143])^(a[343] & b[144])^(a[342] & b[145])^(a[341] & b[146])^(a[340] & b[147])^(a[339] & b[148])^(a[338] & b[149])^(a[337] & b[150])^(a[336] & b[151])^(a[335] & b[152])^(a[334] & b[153])^(a[333] & b[154])^(a[332] & b[155])^(a[331] & b[156])^(a[330] & b[157])^(a[329] & b[158])^(a[328] & b[159])^(a[327] & b[160])^(a[326] & b[161])^(a[325] & b[162])^(a[324] & b[163])^(a[323] & b[164])^(a[322] & b[165])^(a[321] & b[166])^(a[320] & b[167])^(a[319] & b[168])^(a[318] & b[169])^(a[317] & b[170])^(a[316] & b[171])^(a[315] & b[172])^(a[314] & b[173])^(a[313] & b[174])^(a[312] & b[175])^(a[311] & b[176])^(a[310] & b[177])^(a[309] & b[178])^(a[308] & b[179])^(a[307] & b[180])^(a[306] & b[181])^(a[305] & b[182])^(a[304] & b[183])^(a[303] & b[184])^(a[302] & b[185])^(a[301] & b[186])^(a[300] & b[187])^(a[299] & b[188])^(a[298] & b[189])^(a[297] & b[190])^(a[296] & b[191])^(a[295] & b[192])^(a[294] & b[193])^(a[293] & b[194])^(a[292] & b[195])^(a[291] & b[196])^(a[290] & b[197])^(a[289] & b[198])^(a[288] & b[199])^(a[287] & b[200])^(a[286] & b[201])^(a[285] & b[202])^(a[284] & b[203])^(a[283] & b[204])^(a[282] & b[205])^(a[281] & b[206])^(a[280] & b[207])^(a[279] & b[208])^(a[278] & b[209])^(a[277] & b[210])^(a[276] & b[211])^(a[275] & b[212])^(a[274] & b[213])^(a[273] & b[214])^(a[272] & b[215])^(a[271] & b[216])^(a[270] & b[217])^(a[269] & b[218])^(a[268] & b[219])^(a[267] & b[220])^(a[266] & b[221])^(a[265] & b[222])^(a[264] & b[223])^(a[263] & b[224])^(a[262] & b[225])^(a[261] & b[226])^(a[260] & b[227])^(a[259] & b[228])^(a[258] & b[229])^(a[257] & b[230])^(a[256] & b[231])^(a[255] & b[232])^(a[254] & b[233])^(a[253] & b[234])^(a[252] & b[235])^(a[251] & b[236])^(a[250] & b[237])^(a[249] & b[238])^(a[248] & b[239])^(a[247] & b[240])^(a[246] & b[241])^(a[245] & b[242])^(a[244] & b[243])^(a[243] & b[244])^(a[242] & b[245])^(a[241] & b[246])^(a[240] & b[247])^(a[239] & b[248])^(a[238] & b[249])^(a[237] & b[250])^(a[236] & b[251])^(a[235] & b[252])^(a[234] & b[253])^(a[233] & b[254])^(a[232] & b[255])^(a[231] & b[256])^(a[230] & b[257])^(a[229] & b[258])^(a[228] & b[259])^(a[227] & b[260])^(a[226] & b[261])^(a[225] & b[262])^(a[224] & b[263])^(a[223] & b[264])^(a[222] & b[265])^(a[221] & b[266])^(a[220] & b[267])^(a[219] & b[268])^(a[218] & b[269])^(a[217] & b[270])^(a[216] & b[271])^(a[215] & b[272])^(a[214] & b[273])^(a[213] & b[274])^(a[212] & b[275])^(a[211] & b[276])^(a[210] & b[277])^(a[209] & b[278])^(a[208] & b[279])^(a[207] & b[280])^(a[206] & b[281])^(a[205] & b[282])^(a[204] & b[283])^(a[203] & b[284])^(a[202] & b[285])^(a[201] & b[286])^(a[200] & b[287])^(a[199] & b[288])^(a[198] & b[289])^(a[197] & b[290])^(a[196] & b[291])^(a[195] & b[292])^(a[194] & b[293])^(a[193] & b[294])^(a[192] & b[295])^(a[191] & b[296])^(a[190] & b[297])^(a[189] & b[298])^(a[188] & b[299])^(a[187] & b[300])^(a[186] & b[301])^(a[185] & b[302])^(a[184] & b[303])^(a[183] & b[304])^(a[182] & b[305])^(a[181] & b[306])^(a[180] & b[307])^(a[179] & b[308])^(a[178] & b[309])^(a[177] & b[310])^(a[176] & b[311])^(a[175] & b[312])^(a[174] & b[313])^(a[173] & b[314])^(a[172] & b[315])^(a[171] & b[316])^(a[170] & b[317])^(a[169] & b[318])^(a[168] & b[319])^(a[167] & b[320])^(a[166] & b[321])^(a[165] & b[322])^(a[164] & b[323])^(a[163] & b[324])^(a[162] & b[325])^(a[161] & b[326])^(a[160] & b[327])^(a[159] & b[328])^(a[158] & b[329])^(a[157] & b[330])^(a[156] & b[331])^(a[155] & b[332])^(a[154] & b[333])^(a[153] & b[334])^(a[152] & b[335])^(a[151] & b[336])^(a[150] & b[337])^(a[149] & b[338])^(a[148] & b[339])^(a[147] & b[340])^(a[146] & b[341])^(a[145] & b[342])^(a[144] & b[343])^(a[143] & b[344])^(a[142] & b[345])^(a[141] & b[346])^(a[140] & b[347])^(a[139] & b[348])^(a[138] & b[349])^(a[137] & b[350])^(a[136] & b[351])^(a[135] & b[352])^(a[134] & b[353])^(a[133] & b[354])^(a[132] & b[355])^(a[131] & b[356])^(a[130] & b[357])^(a[129] & b[358])^(a[128] & b[359])^(a[127] & b[360])^(a[126] & b[361])^(a[125] & b[362])^(a[124] & b[363])^(a[123] & b[364])^(a[122] & b[365])^(a[121] & b[366])^(a[120] & b[367])^(a[119] & b[368])^(a[118] & b[369])^(a[117] & b[370])^(a[116] & b[371])^(a[115] & b[372])^(a[114] & b[373])^(a[113] & b[374])^(a[112] & b[375])^(a[111] & b[376])^(a[110] & b[377])^(a[109] & b[378])^(a[108] & b[379])^(a[107] & b[380])^(a[106] & b[381])^(a[105] & b[382])^(a[104] & b[383])^(a[103] & b[384])^(a[102] & b[385])^(a[101] & b[386])^(a[100] & b[387])^(a[99] & b[388])^(a[98] & b[389])^(a[97] & b[390])^(a[96] & b[391])^(a[95] & b[392])^(a[94] & b[393])^(a[93] & b[394])^(a[92] & b[395])^(a[91] & b[396])^(a[90] & b[397])^(a[89] & b[398])^(a[88] & b[399])^(a[87] & b[400])^(a[86] & b[401])^(a[85] & b[402])^(a[84] & b[403])^(a[83] & b[404])^(a[82] & b[405])^(a[81] & b[406])^(a[80] & b[407])^(a[79] & b[408]);
assign y[488] = (a[408] & b[80])^(a[407] & b[81])^(a[406] & b[82])^(a[405] & b[83])^(a[404] & b[84])^(a[403] & b[85])^(a[402] & b[86])^(a[401] & b[87])^(a[400] & b[88])^(a[399] & b[89])^(a[398] & b[90])^(a[397] & b[91])^(a[396] & b[92])^(a[395] & b[93])^(a[394] & b[94])^(a[393] & b[95])^(a[392] & b[96])^(a[391] & b[97])^(a[390] & b[98])^(a[389] & b[99])^(a[388] & b[100])^(a[387] & b[101])^(a[386] & b[102])^(a[385] & b[103])^(a[384] & b[104])^(a[383] & b[105])^(a[382] & b[106])^(a[381] & b[107])^(a[380] & b[108])^(a[379] & b[109])^(a[378] & b[110])^(a[377] & b[111])^(a[376] & b[112])^(a[375] & b[113])^(a[374] & b[114])^(a[373] & b[115])^(a[372] & b[116])^(a[371] & b[117])^(a[370] & b[118])^(a[369] & b[119])^(a[368] & b[120])^(a[367] & b[121])^(a[366] & b[122])^(a[365] & b[123])^(a[364] & b[124])^(a[363] & b[125])^(a[362] & b[126])^(a[361] & b[127])^(a[360] & b[128])^(a[359] & b[129])^(a[358] & b[130])^(a[357] & b[131])^(a[356] & b[132])^(a[355] & b[133])^(a[354] & b[134])^(a[353] & b[135])^(a[352] & b[136])^(a[351] & b[137])^(a[350] & b[138])^(a[349] & b[139])^(a[348] & b[140])^(a[347] & b[141])^(a[346] & b[142])^(a[345] & b[143])^(a[344] & b[144])^(a[343] & b[145])^(a[342] & b[146])^(a[341] & b[147])^(a[340] & b[148])^(a[339] & b[149])^(a[338] & b[150])^(a[337] & b[151])^(a[336] & b[152])^(a[335] & b[153])^(a[334] & b[154])^(a[333] & b[155])^(a[332] & b[156])^(a[331] & b[157])^(a[330] & b[158])^(a[329] & b[159])^(a[328] & b[160])^(a[327] & b[161])^(a[326] & b[162])^(a[325] & b[163])^(a[324] & b[164])^(a[323] & b[165])^(a[322] & b[166])^(a[321] & b[167])^(a[320] & b[168])^(a[319] & b[169])^(a[318] & b[170])^(a[317] & b[171])^(a[316] & b[172])^(a[315] & b[173])^(a[314] & b[174])^(a[313] & b[175])^(a[312] & b[176])^(a[311] & b[177])^(a[310] & b[178])^(a[309] & b[179])^(a[308] & b[180])^(a[307] & b[181])^(a[306] & b[182])^(a[305] & b[183])^(a[304] & b[184])^(a[303] & b[185])^(a[302] & b[186])^(a[301] & b[187])^(a[300] & b[188])^(a[299] & b[189])^(a[298] & b[190])^(a[297] & b[191])^(a[296] & b[192])^(a[295] & b[193])^(a[294] & b[194])^(a[293] & b[195])^(a[292] & b[196])^(a[291] & b[197])^(a[290] & b[198])^(a[289] & b[199])^(a[288] & b[200])^(a[287] & b[201])^(a[286] & b[202])^(a[285] & b[203])^(a[284] & b[204])^(a[283] & b[205])^(a[282] & b[206])^(a[281] & b[207])^(a[280] & b[208])^(a[279] & b[209])^(a[278] & b[210])^(a[277] & b[211])^(a[276] & b[212])^(a[275] & b[213])^(a[274] & b[214])^(a[273] & b[215])^(a[272] & b[216])^(a[271] & b[217])^(a[270] & b[218])^(a[269] & b[219])^(a[268] & b[220])^(a[267] & b[221])^(a[266] & b[222])^(a[265] & b[223])^(a[264] & b[224])^(a[263] & b[225])^(a[262] & b[226])^(a[261] & b[227])^(a[260] & b[228])^(a[259] & b[229])^(a[258] & b[230])^(a[257] & b[231])^(a[256] & b[232])^(a[255] & b[233])^(a[254] & b[234])^(a[253] & b[235])^(a[252] & b[236])^(a[251] & b[237])^(a[250] & b[238])^(a[249] & b[239])^(a[248] & b[240])^(a[247] & b[241])^(a[246] & b[242])^(a[245] & b[243])^(a[244] & b[244])^(a[243] & b[245])^(a[242] & b[246])^(a[241] & b[247])^(a[240] & b[248])^(a[239] & b[249])^(a[238] & b[250])^(a[237] & b[251])^(a[236] & b[252])^(a[235] & b[253])^(a[234] & b[254])^(a[233] & b[255])^(a[232] & b[256])^(a[231] & b[257])^(a[230] & b[258])^(a[229] & b[259])^(a[228] & b[260])^(a[227] & b[261])^(a[226] & b[262])^(a[225] & b[263])^(a[224] & b[264])^(a[223] & b[265])^(a[222] & b[266])^(a[221] & b[267])^(a[220] & b[268])^(a[219] & b[269])^(a[218] & b[270])^(a[217] & b[271])^(a[216] & b[272])^(a[215] & b[273])^(a[214] & b[274])^(a[213] & b[275])^(a[212] & b[276])^(a[211] & b[277])^(a[210] & b[278])^(a[209] & b[279])^(a[208] & b[280])^(a[207] & b[281])^(a[206] & b[282])^(a[205] & b[283])^(a[204] & b[284])^(a[203] & b[285])^(a[202] & b[286])^(a[201] & b[287])^(a[200] & b[288])^(a[199] & b[289])^(a[198] & b[290])^(a[197] & b[291])^(a[196] & b[292])^(a[195] & b[293])^(a[194] & b[294])^(a[193] & b[295])^(a[192] & b[296])^(a[191] & b[297])^(a[190] & b[298])^(a[189] & b[299])^(a[188] & b[300])^(a[187] & b[301])^(a[186] & b[302])^(a[185] & b[303])^(a[184] & b[304])^(a[183] & b[305])^(a[182] & b[306])^(a[181] & b[307])^(a[180] & b[308])^(a[179] & b[309])^(a[178] & b[310])^(a[177] & b[311])^(a[176] & b[312])^(a[175] & b[313])^(a[174] & b[314])^(a[173] & b[315])^(a[172] & b[316])^(a[171] & b[317])^(a[170] & b[318])^(a[169] & b[319])^(a[168] & b[320])^(a[167] & b[321])^(a[166] & b[322])^(a[165] & b[323])^(a[164] & b[324])^(a[163] & b[325])^(a[162] & b[326])^(a[161] & b[327])^(a[160] & b[328])^(a[159] & b[329])^(a[158] & b[330])^(a[157] & b[331])^(a[156] & b[332])^(a[155] & b[333])^(a[154] & b[334])^(a[153] & b[335])^(a[152] & b[336])^(a[151] & b[337])^(a[150] & b[338])^(a[149] & b[339])^(a[148] & b[340])^(a[147] & b[341])^(a[146] & b[342])^(a[145] & b[343])^(a[144] & b[344])^(a[143] & b[345])^(a[142] & b[346])^(a[141] & b[347])^(a[140] & b[348])^(a[139] & b[349])^(a[138] & b[350])^(a[137] & b[351])^(a[136] & b[352])^(a[135] & b[353])^(a[134] & b[354])^(a[133] & b[355])^(a[132] & b[356])^(a[131] & b[357])^(a[130] & b[358])^(a[129] & b[359])^(a[128] & b[360])^(a[127] & b[361])^(a[126] & b[362])^(a[125] & b[363])^(a[124] & b[364])^(a[123] & b[365])^(a[122] & b[366])^(a[121] & b[367])^(a[120] & b[368])^(a[119] & b[369])^(a[118] & b[370])^(a[117] & b[371])^(a[116] & b[372])^(a[115] & b[373])^(a[114] & b[374])^(a[113] & b[375])^(a[112] & b[376])^(a[111] & b[377])^(a[110] & b[378])^(a[109] & b[379])^(a[108] & b[380])^(a[107] & b[381])^(a[106] & b[382])^(a[105] & b[383])^(a[104] & b[384])^(a[103] & b[385])^(a[102] & b[386])^(a[101] & b[387])^(a[100] & b[388])^(a[99] & b[389])^(a[98] & b[390])^(a[97] & b[391])^(a[96] & b[392])^(a[95] & b[393])^(a[94] & b[394])^(a[93] & b[395])^(a[92] & b[396])^(a[91] & b[397])^(a[90] & b[398])^(a[89] & b[399])^(a[88] & b[400])^(a[87] & b[401])^(a[86] & b[402])^(a[85] & b[403])^(a[84] & b[404])^(a[83] & b[405])^(a[82] & b[406])^(a[81] & b[407])^(a[80] & b[408]);
assign y[489] = (a[408] & b[81])^(a[407] & b[82])^(a[406] & b[83])^(a[405] & b[84])^(a[404] & b[85])^(a[403] & b[86])^(a[402] & b[87])^(a[401] & b[88])^(a[400] & b[89])^(a[399] & b[90])^(a[398] & b[91])^(a[397] & b[92])^(a[396] & b[93])^(a[395] & b[94])^(a[394] & b[95])^(a[393] & b[96])^(a[392] & b[97])^(a[391] & b[98])^(a[390] & b[99])^(a[389] & b[100])^(a[388] & b[101])^(a[387] & b[102])^(a[386] & b[103])^(a[385] & b[104])^(a[384] & b[105])^(a[383] & b[106])^(a[382] & b[107])^(a[381] & b[108])^(a[380] & b[109])^(a[379] & b[110])^(a[378] & b[111])^(a[377] & b[112])^(a[376] & b[113])^(a[375] & b[114])^(a[374] & b[115])^(a[373] & b[116])^(a[372] & b[117])^(a[371] & b[118])^(a[370] & b[119])^(a[369] & b[120])^(a[368] & b[121])^(a[367] & b[122])^(a[366] & b[123])^(a[365] & b[124])^(a[364] & b[125])^(a[363] & b[126])^(a[362] & b[127])^(a[361] & b[128])^(a[360] & b[129])^(a[359] & b[130])^(a[358] & b[131])^(a[357] & b[132])^(a[356] & b[133])^(a[355] & b[134])^(a[354] & b[135])^(a[353] & b[136])^(a[352] & b[137])^(a[351] & b[138])^(a[350] & b[139])^(a[349] & b[140])^(a[348] & b[141])^(a[347] & b[142])^(a[346] & b[143])^(a[345] & b[144])^(a[344] & b[145])^(a[343] & b[146])^(a[342] & b[147])^(a[341] & b[148])^(a[340] & b[149])^(a[339] & b[150])^(a[338] & b[151])^(a[337] & b[152])^(a[336] & b[153])^(a[335] & b[154])^(a[334] & b[155])^(a[333] & b[156])^(a[332] & b[157])^(a[331] & b[158])^(a[330] & b[159])^(a[329] & b[160])^(a[328] & b[161])^(a[327] & b[162])^(a[326] & b[163])^(a[325] & b[164])^(a[324] & b[165])^(a[323] & b[166])^(a[322] & b[167])^(a[321] & b[168])^(a[320] & b[169])^(a[319] & b[170])^(a[318] & b[171])^(a[317] & b[172])^(a[316] & b[173])^(a[315] & b[174])^(a[314] & b[175])^(a[313] & b[176])^(a[312] & b[177])^(a[311] & b[178])^(a[310] & b[179])^(a[309] & b[180])^(a[308] & b[181])^(a[307] & b[182])^(a[306] & b[183])^(a[305] & b[184])^(a[304] & b[185])^(a[303] & b[186])^(a[302] & b[187])^(a[301] & b[188])^(a[300] & b[189])^(a[299] & b[190])^(a[298] & b[191])^(a[297] & b[192])^(a[296] & b[193])^(a[295] & b[194])^(a[294] & b[195])^(a[293] & b[196])^(a[292] & b[197])^(a[291] & b[198])^(a[290] & b[199])^(a[289] & b[200])^(a[288] & b[201])^(a[287] & b[202])^(a[286] & b[203])^(a[285] & b[204])^(a[284] & b[205])^(a[283] & b[206])^(a[282] & b[207])^(a[281] & b[208])^(a[280] & b[209])^(a[279] & b[210])^(a[278] & b[211])^(a[277] & b[212])^(a[276] & b[213])^(a[275] & b[214])^(a[274] & b[215])^(a[273] & b[216])^(a[272] & b[217])^(a[271] & b[218])^(a[270] & b[219])^(a[269] & b[220])^(a[268] & b[221])^(a[267] & b[222])^(a[266] & b[223])^(a[265] & b[224])^(a[264] & b[225])^(a[263] & b[226])^(a[262] & b[227])^(a[261] & b[228])^(a[260] & b[229])^(a[259] & b[230])^(a[258] & b[231])^(a[257] & b[232])^(a[256] & b[233])^(a[255] & b[234])^(a[254] & b[235])^(a[253] & b[236])^(a[252] & b[237])^(a[251] & b[238])^(a[250] & b[239])^(a[249] & b[240])^(a[248] & b[241])^(a[247] & b[242])^(a[246] & b[243])^(a[245] & b[244])^(a[244] & b[245])^(a[243] & b[246])^(a[242] & b[247])^(a[241] & b[248])^(a[240] & b[249])^(a[239] & b[250])^(a[238] & b[251])^(a[237] & b[252])^(a[236] & b[253])^(a[235] & b[254])^(a[234] & b[255])^(a[233] & b[256])^(a[232] & b[257])^(a[231] & b[258])^(a[230] & b[259])^(a[229] & b[260])^(a[228] & b[261])^(a[227] & b[262])^(a[226] & b[263])^(a[225] & b[264])^(a[224] & b[265])^(a[223] & b[266])^(a[222] & b[267])^(a[221] & b[268])^(a[220] & b[269])^(a[219] & b[270])^(a[218] & b[271])^(a[217] & b[272])^(a[216] & b[273])^(a[215] & b[274])^(a[214] & b[275])^(a[213] & b[276])^(a[212] & b[277])^(a[211] & b[278])^(a[210] & b[279])^(a[209] & b[280])^(a[208] & b[281])^(a[207] & b[282])^(a[206] & b[283])^(a[205] & b[284])^(a[204] & b[285])^(a[203] & b[286])^(a[202] & b[287])^(a[201] & b[288])^(a[200] & b[289])^(a[199] & b[290])^(a[198] & b[291])^(a[197] & b[292])^(a[196] & b[293])^(a[195] & b[294])^(a[194] & b[295])^(a[193] & b[296])^(a[192] & b[297])^(a[191] & b[298])^(a[190] & b[299])^(a[189] & b[300])^(a[188] & b[301])^(a[187] & b[302])^(a[186] & b[303])^(a[185] & b[304])^(a[184] & b[305])^(a[183] & b[306])^(a[182] & b[307])^(a[181] & b[308])^(a[180] & b[309])^(a[179] & b[310])^(a[178] & b[311])^(a[177] & b[312])^(a[176] & b[313])^(a[175] & b[314])^(a[174] & b[315])^(a[173] & b[316])^(a[172] & b[317])^(a[171] & b[318])^(a[170] & b[319])^(a[169] & b[320])^(a[168] & b[321])^(a[167] & b[322])^(a[166] & b[323])^(a[165] & b[324])^(a[164] & b[325])^(a[163] & b[326])^(a[162] & b[327])^(a[161] & b[328])^(a[160] & b[329])^(a[159] & b[330])^(a[158] & b[331])^(a[157] & b[332])^(a[156] & b[333])^(a[155] & b[334])^(a[154] & b[335])^(a[153] & b[336])^(a[152] & b[337])^(a[151] & b[338])^(a[150] & b[339])^(a[149] & b[340])^(a[148] & b[341])^(a[147] & b[342])^(a[146] & b[343])^(a[145] & b[344])^(a[144] & b[345])^(a[143] & b[346])^(a[142] & b[347])^(a[141] & b[348])^(a[140] & b[349])^(a[139] & b[350])^(a[138] & b[351])^(a[137] & b[352])^(a[136] & b[353])^(a[135] & b[354])^(a[134] & b[355])^(a[133] & b[356])^(a[132] & b[357])^(a[131] & b[358])^(a[130] & b[359])^(a[129] & b[360])^(a[128] & b[361])^(a[127] & b[362])^(a[126] & b[363])^(a[125] & b[364])^(a[124] & b[365])^(a[123] & b[366])^(a[122] & b[367])^(a[121] & b[368])^(a[120] & b[369])^(a[119] & b[370])^(a[118] & b[371])^(a[117] & b[372])^(a[116] & b[373])^(a[115] & b[374])^(a[114] & b[375])^(a[113] & b[376])^(a[112] & b[377])^(a[111] & b[378])^(a[110] & b[379])^(a[109] & b[380])^(a[108] & b[381])^(a[107] & b[382])^(a[106] & b[383])^(a[105] & b[384])^(a[104] & b[385])^(a[103] & b[386])^(a[102] & b[387])^(a[101] & b[388])^(a[100] & b[389])^(a[99] & b[390])^(a[98] & b[391])^(a[97] & b[392])^(a[96] & b[393])^(a[95] & b[394])^(a[94] & b[395])^(a[93] & b[396])^(a[92] & b[397])^(a[91] & b[398])^(a[90] & b[399])^(a[89] & b[400])^(a[88] & b[401])^(a[87] & b[402])^(a[86] & b[403])^(a[85] & b[404])^(a[84] & b[405])^(a[83] & b[406])^(a[82] & b[407])^(a[81] & b[408]);
assign y[490] = (a[408] & b[82])^(a[407] & b[83])^(a[406] & b[84])^(a[405] & b[85])^(a[404] & b[86])^(a[403] & b[87])^(a[402] & b[88])^(a[401] & b[89])^(a[400] & b[90])^(a[399] & b[91])^(a[398] & b[92])^(a[397] & b[93])^(a[396] & b[94])^(a[395] & b[95])^(a[394] & b[96])^(a[393] & b[97])^(a[392] & b[98])^(a[391] & b[99])^(a[390] & b[100])^(a[389] & b[101])^(a[388] & b[102])^(a[387] & b[103])^(a[386] & b[104])^(a[385] & b[105])^(a[384] & b[106])^(a[383] & b[107])^(a[382] & b[108])^(a[381] & b[109])^(a[380] & b[110])^(a[379] & b[111])^(a[378] & b[112])^(a[377] & b[113])^(a[376] & b[114])^(a[375] & b[115])^(a[374] & b[116])^(a[373] & b[117])^(a[372] & b[118])^(a[371] & b[119])^(a[370] & b[120])^(a[369] & b[121])^(a[368] & b[122])^(a[367] & b[123])^(a[366] & b[124])^(a[365] & b[125])^(a[364] & b[126])^(a[363] & b[127])^(a[362] & b[128])^(a[361] & b[129])^(a[360] & b[130])^(a[359] & b[131])^(a[358] & b[132])^(a[357] & b[133])^(a[356] & b[134])^(a[355] & b[135])^(a[354] & b[136])^(a[353] & b[137])^(a[352] & b[138])^(a[351] & b[139])^(a[350] & b[140])^(a[349] & b[141])^(a[348] & b[142])^(a[347] & b[143])^(a[346] & b[144])^(a[345] & b[145])^(a[344] & b[146])^(a[343] & b[147])^(a[342] & b[148])^(a[341] & b[149])^(a[340] & b[150])^(a[339] & b[151])^(a[338] & b[152])^(a[337] & b[153])^(a[336] & b[154])^(a[335] & b[155])^(a[334] & b[156])^(a[333] & b[157])^(a[332] & b[158])^(a[331] & b[159])^(a[330] & b[160])^(a[329] & b[161])^(a[328] & b[162])^(a[327] & b[163])^(a[326] & b[164])^(a[325] & b[165])^(a[324] & b[166])^(a[323] & b[167])^(a[322] & b[168])^(a[321] & b[169])^(a[320] & b[170])^(a[319] & b[171])^(a[318] & b[172])^(a[317] & b[173])^(a[316] & b[174])^(a[315] & b[175])^(a[314] & b[176])^(a[313] & b[177])^(a[312] & b[178])^(a[311] & b[179])^(a[310] & b[180])^(a[309] & b[181])^(a[308] & b[182])^(a[307] & b[183])^(a[306] & b[184])^(a[305] & b[185])^(a[304] & b[186])^(a[303] & b[187])^(a[302] & b[188])^(a[301] & b[189])^(a[300] & b[190])^(a[299] & b[191])^(a[298] & b[192])^(a[297] & b[193])^(a[296] & b[194])^(a[295] & b[195])^(a[294] & b[196])^(a[293] & b[197])^(a[292] & b[198])^(a[291] & b[199])^(a[290] & b[200])^(a[289] & b[201])^(a[288] & b[202])^(a[287] & b[203])^(a[286] & b[204])^(a[285] & b[205])^(a[284] & b[206])^(a[283] & b[207])^(a[282] & b[208])^(a[281] & b[209])^(a[280] & b[210])^(a[279] & b[211])^(a[278] & b[212])^(a[277] & b[213])^(a[276] & b[214])^(a[275] & b[215])^(a[274] & b[216])^(a[273] & b[217])^(a[272] & b[218])^(a[271] & b[219])^(a[270] & b[220])^(a[269] & b[221])^(a[268] & b[222])^(a[267] & b[223])^(a[266] & b[224])^(a[265] & b[225])^(a[264] & b[226])^(a[263] & b[227])^(a[262] & b[228])^(a[261] & b[229])^(a[260] & b[230])^(a[259] & b[231])^(a[258] & b[232])^(a[257] & b[233])^(a[256] & b[234])^(a[255] & b[235])^(a[254] & b[236])^(a[253] & b[237])^(a[252] & b[238])^(a[251] & b[239])^(a[250] & b[240])^(a[249] & b[241])^(a[248] & b[242])^(a[247] & b[243])^(a[246] & b[244])^(a[245] & b[245])^(a[244] & b[246])^(a[243] & b[247])^(a[242] & b[248])^(a[241] & b[249])^(a[240] & b[250])^(a[239] & b[251])^(a[238] & b[252])^(a[237] & b[253])^(a[236] & b[254])^(a[235] & b[255])^(a[234] & b[256])^(a[233] & b[257])^(a[232] & b[258])^(a[231] & b[259])^(a[230] & b[260])^(a[229] & b[261])^(a[228] & b[262])^(a[227] & b[263])^(a[226] & b[264])^(a[225] & b[265])^(a[224] & b[266])^(a[223] & b[267])^(a[222] & b[268])^(a[221] & b[269])^(a[220] & b[270])^(a[219] & b[271])^(a[218] & b[272])^(a[217] & b[273])^(a[216] & b[274])^(a[215] & b[275])^(a[214] & b[276])^(a[213] & b[277])^(a[212] & b[278])^(a[211] & b[279])^(a[210] & b[280])^(a[209] & b[281])^(a[208] & b[282])^(a[207] & b[283])^(a[206] & b[284])^(a[205] & b[285])^(a[204] & b[286])^(a[203] & b[287])^(a[202] & b[288])^(a[201] & b[289])^(a[200] & b[290])^(a[199] & b[291])^(a[198] & b[292])^(a[197] & b[293])^(a[196] & b[294])^(a[195] & b[295])^(a[194] & b[296])^(a[193] & b[297])^(a[192] & b[298])^(a[191] & b[299])^(a[190] & b[300])^(a[189] & b[301])^(a[188] & b[302])^(a[187] & b[303])^(a[186] & b[304])^(a[185] & b[305])^(a[184] & b[306])^(a[183] & b[307])^(a[182] & b[308])^(a[181] & b[309])^(a[180] & b[310])^(a[179] & b[311])^(a[178] & b[312])^(a[177] & b[313])^(a[176] & b[314])^(a[175] & b[315])^(a[174] & b[316])^(a[173] & b[317])^(a[172] & b[318])^(a[171] & b[319])^(a[170] & b[320])^(a[169] & b[321])^(a[168] & b[322])^(a[167] & b[323])^(a[166] & b[324])^(a[165] & b[325])^(a[164] & b[326])^(a[163] & b[327])^(a[162] & b[328])^(a[161] & b[329])^(a[160] & b[330])^(a[159] & b[331])^(a[158] & b[332])^(a[157] & b[333])^(a[156] & b[334])^(a[155] & b[335])^(a[154] & b[336])^(a[153] & b[337])^(a[152] & b[338])^(a[151] & b[339])^(a[150] & b[340])^(a[149] & b[341])^(a[148] & b[342])^(a[147] & b[343])^(a[146] & b[344])^(a[145] & b[345])^(a[144] & b[346])^(a[143] & b[347])^(a[142] & b[348])^(a[141] & b[349])^(a[140] & b[350])^(a[139] & b[351])^(a[138] & b[352])^(a[137] & b[353])^(a[136] & b[354])^(a[135] & b[355])^(a[134] & b[356])^(a[133] & b[357])^(a[132] & b[358])^(a[131] & b[359])^(a[130] & b[360])^(a[129] & b[361])^(a[128] & b[362])^(a[127] & b[363])^(a[126] & b[364])^(a[125] & b[365])^(a[124] & b[366])^(a[123] & b[367])^(a[122] & b[368])^(a[121] & b[369])^(a[120] & b[370])^(a[119] & b[371])^(a[118] & b[372])^(a[117] & b[373])^(a[116] & b[374])^(a[115] & b[375])^(a[114] & b[376])^(a[113] & b[377])^(a[112] & b[378])^(a[111] & b[379])^(a[110] & b[380])^(a[109] & b[381])^(a[108] & b[382])^(a[107] & b[383])^(a[106] & b[384])^(a[105] & b[385])^(a[104] & b[386])^(a[103] & b[387])^(a[102] & b[388])^(a[101] & b[389])^(a[100] & b[390])^(a[99] & b[391])^(a[98] & b[392])^(a[97] & b[393])^(a[96] & b[394])^(a[95] & b[395])^(a[94] & b[396])^(a[93] & b[397])^(a[92] & b[398])^(a[91] & b[399])^(a[90] & b[400])^(a[89] & b[401])^(a[88] & b[402])^(a[87] & b[403])^(a[86] & b[404])^(a[85] & b[405])^(a[84] & b[406])^(a[83] & b[407])^(a[82] & b[408]);
assign y[491] = (a[408] & b[83])^(a[407] & b[84])^(a[406] & b[85])^(a[405] & b[86])^(a[404] & b[87])^(a[403] & b[88])^(a[402] & b[89])^(a[401] & b[90])^(a[400] & b[91])^(a[399] & b[92])^(a[398] & b[93])^(a[397] & b[94])^(a[396] & b[95])^(a[395] & b[96])^(a[394] & b[97])^(a[393] & b[98])^(a[392] & b[99])^(a[391] & b[100])^(a[390] & b[101])^(a[389] & b[102])^(a[388] & b[103])^(a[387] & b[104])^(a[386] & b[105])^(a[385] & b[106])^(a[384] & b[107])^(a[383] & b[108])^(a[382] & b[109])^(a[381] & b[110])^(a[380] & b[111])^(a[379] & b[112])^(a[378] & b[113])^(a[377] & b[114])^(a[376] & b[115])^(a[375] & b[116])^(a[374] & b[117])^(a[373] & b[118])^(a[372] & b[119])^(a[371] & b[120])^(a[370] & b[121])^(a[369] & b[122])^(a[368] & b[123])^(a[367] & b[124])^(a[366] & b[125])^(a[365] & b[126])^(a[364] & b[127])^(a[363] & b[128])^(a[362] & b[129])^(a[361] & b[130])^(a[360] & b[131])^(a[359] & b[132])^(a[358] & b[133])^(a[357] & b[134])^(a[356] & b[135])^(a[355] & b[136])^(a[354] & b[137])^(a[353] & b[138])^(a[352] & b[139])^(a[351] & b[140])^(a[350] & b[141])^(a[349] & b[142])^(a[348] & b[143])^(a[347] & b[144])^(a[346] & b[145])^(a[345] & b[146])^(a[344] & b[147])^(a[343] & b[148])^(a[342] & b[149])^(a[341] & b[150])^(a[340] & b[151])^(a[339] & b[152])^(a[338] & b[153])^(a[337] & b[154])^(a[336] & b[155])^(a[335] & b[156])^(a[334] & b[157])^(a[333] & b[158])^(a[332] & b[159])^(a[331] & b[160])^(a[330] & b[161])^(a[329] & b[162])^(a[328] & b[163])^(a[327] & b[164])^(a[326] & b[165])^(a[325] & b[166])^(a[324] & b[167])^(a[323] & b[168])^(a[322] & b[169])^(a[321] & b[170])^(a[320] & b[171])^(a[319] & b[172])^(a[318] & b[173])^(a[317] & b[174])^(a[316] & b[175])^(a[315] & b[176])^(a[314] & b[177])^(a[313] & b[178])^(a[312] & b[179])^(a[311] & b[180])^(a[310] & b[181])^(a[309] & b[182])^(a[308] & b[183])^(a[307] & b[184])^(a[306] & b[185])^(a[305] & b[186])^(a[304] & b[187])^(a[303] & b[188])^(a[302] & b[189])^(a[301] & b[190])^(a[300] & b[191])^(a[299] & b[192])^(a[298] & b[193])^(a[297] & b[194])^(a[296] & b[195])^(a[295] & b[196])^(a[294] & b[197])^(a[293] & b[198])^(a[292] & b[199])^(a[291] & b[200])^(a[290] & b[201])^(a[289] & b[202])^(a[288] & b[203])^(a[287] & b[204])^(a[286] & b[205])^(a[285] & b[206])^(a[284] & b[207])^(a[283] & b[208])^(a[282] & b[209])^(a[281] & b[210])^(a[280] & b[211])^(a[279] & b[212])^(a[278] & b[213])^(a[277] & b[214])^(a[276] & b[215])^(a[275] & b[216])^(a[274] & b[217])^(a[273] & b[218])^(a[272] & b[219])^(a[271] & b[220])^(a[270] & b[221])^(a[269] & b[222])^(a[268] & b[223])^(a[267] & b[224])^(a[266] & b[225])^(a[265] & b[226])^(a[264] & b[227])^(a[263] & b[228])^(a[262] & b[229])^(a[261] & b[230])^(a[260] & b[231])^(a[259] & b[232])^(a[258] & b[233])^(a[257] & b[234])^(a[256] & b[235])^(a[255] & b[236])^(a[254] & b[237])^(a[253] & b[238])^(a[252] & b[239])^(a[251] & b[240])^(a[250] & b[241])^(a[249] & b[242])^(a[248] & b[243])^(a[247] & b[244])^(a[246] & b[245])^(a[245] & b[246])^(a[244] & b[247])^(a[243] & b[248])^(a[242] & b[249])^(a[241] & b[250])^(a[240] & b[251])^(a[239] & b[252])^(a[238] & b[253])^(a[237] & b[254])^(a[236] & b[255])^(a[235] & b[256])^(a[234] & b[257])^(a[233] & b[258])^(a[232] & b[259])^(a[231] & b[260])^(a[230] & b[261])^(a[229] & b[262])^(a[228] & b[263])^(a[227] & b[264])^(a[226] & b[265])^(a[225] & b[266])^(a[224] & b[267])^(a[223] & b[268])^(a[222] & b[269])^(a[221] & b[270])^(a[220] & b[271])^(a[219] & b[272])^(a[218] & b[273])^(a[217] & b[274])^(a[216] & b[275])^(a[215] & b[276])^(a[214] & b[277])^(a[213] & b[278])^(a[212] & b[279])^(a[211] & b[280])^(a[210] & b[281])^(a[209] & b[282])^(a[208] & b[283])^(a[207] & b[284])^(a[206] & b[285])^(a[205] & b[286])^(a[204] & b[287])^(a[203] & b[288])^(a[202] & b[289])^(a[201] & b[290])^(a[200] & b[291])^(a[199] & b[292])^(a[198] & b[293])^(a[197] & b[294])^(a[196] & b[295])^(a[195] & b[296])^(a[194] & b[297])^(a[193] & b[298])^(a[192] & b[299])^(a[191] & b[300])^(a[190] & b[301])^(a[189] & b[302])^(a[188] & b[303])^(a[187] & b[304])^(a[186] & b[305])^(a[185] & b[306])^(a[184] & b[307])^(a[183] & b[308])^(a[182] & b[309])^(a[181] & b[310])^(a[180] & b[311])^(a[179] & b[312])^(a[178] & b[313])^(a[177] & b[314])^(a[176] & b[315])^(a[175] & b[316])^(a[174] & b[317])^(a[173] & b[318])^(a[172] & b[319])^(a[171] & b[320])^(a[170] & b[321])^(a[169] & b[322])^(a[168] & b[323])^(a[167] & b[324])^(a[166] & b[325])^(a[165] & b[326])^(a[164] & b[327])^(a[163] & b[328])^(a[162] & b[329])^(a[161] & b[330])^(a[160] & b[331])^(a[159] & b[332])^(a[158] & b[333])^(a[157] & b[334])^(a[156] & b[335])^(a[155] & b[336])^(a[154] & b[337])^(a[153] & b[338])^(a[152] & b[339])^(a[151] & b[340])^(a[150] & b[341])^(a[149] & b[342])^(a[148] & b[343])^(a[147] & b[344])^(a[146] & b[345])^(a[145] & b[346])^(a[144] & b[347])^(a[143] & b[348])^(a[142] & b[349])^(a[141] & b[350])^(a[140] & b[351])^(a[139] & b[352])^(a[138] & b[353])^(a[137] & b[354])^(a[136] & b[355])^(a[135] & b[356])^(a[134] & b[357])^(a[133] & b[358])^(a[132] & b[359])^(a[131] & b[360])^(a[130] & b[361])^(a[129] & b[362])^(a[128] & b[363])^(a[127] & b[364])^(a[126] & b[365])^(a[125] & b[366])^(a[124] & b[367])^(a[123] & b[368])^(a[122] & b[369])^(a[121] & b[370])^(a[120] & b[371])^(a[119] & b[372])^(a[118] & b[373])^(a[117] & b[374])^(a[116] & b[375])^(a[115] & b[376])^(a[114] & b[377])^(a[113] & b[378])^(a[112] & b[379])^(a[111] & b[380])^(a[110] & b[381])^(a[109] & b[382])^(a[108] & b[383])^(a[107] & b[384])^(a[106] & b[385])^(a[105] & b[386])^(a[104] & b[387])^(a[103] & b[388])^(a[102] & b[389])^(a[101] & b[390])^(a[100] & b[391])^(a[99] & b[392])^(a[98] & b[393])^(a[97] & b[394])^(a[96] & b[395])^(a[95] & b[396])^(a[94] & b[397])^(a[93] & b[398])^(a[92] & b[399])^(a[91] & b[400])^(a[90] & b[401])^(a[89] & b[402])^(a[88] & b[403])^(a[87] & b[404])^(a[86] & b[405])^(a[85] & b[406])^(a[84] & b[407])^(a[83] & b[408]);
assign y[492] = (a[408] & b[84])^(a[407] & b[85])^(a[406] & b[86])^(a[405] & b[87])^(a[404] & b[88])^(a[403] & b[89])^(a[402] & b[90])^(a[401] & b[91])^(a[400] & b[92])^(a[399] & b[93])^(a[398] & b[94])^(a[397] & b[95])^(a[396] & b[96])^(a[395] & b[97])^(a[394] & b[98])^(a[393] & b[99])^(a[392] & b[100])^(a[391] & b[101])^(a[390] & b[102])^(a[389] & b[103])^(a[388] & b[104])^(a[387] & b[105])^(a[386] & b[106])^(a[385] & b[107])^(a[384] & b[108])^(a[383] & b[109])^(a[382] & b[110])^(a[381] & b[111])^(a[380] & b[112])^(a[379] & b[113])^(a[378] & b[114])^(a[377] & b[115])^(a[376] & b[116])^(a[375] & b[117])^(a[374] & b[118])^(a[373] & b[119])^(a[372] & b[120])^(a[371] & b[121])^(a[370] & b[122])^(a[369] & b[123])^(a[368] & b[124])^(a[367] & b[125])^(a[366] & b[126])^(a[365] & b[127])^(a[364] & b[128])^(a[363] & b[129])^(a[362] & b[130])^(a[361] & b[131])^(a[360] & b[132])^(a[359] & b[133])^(a[358] & b[134])^(a[357] & b[135])^(a[356] & b[136])^(a[355] & b[137])^(a[354] & b[138])^(a[353] & b[139])^(a[352] & b[140])^(a[351] & b[141])^(a[350] & b[142])^(a[349] & b[143])^(a[348] & b[144])^(a[347] & b[145])^(a[346] & b[146])^(a[345] & b[147])^(a[344] & b[148])^(a[343] & b[149])^(a[342] & b[150])^(a[341] & b[151])^(a[340] & b[152])^(a[339] & b[153])^(a[338] & b[154])^(a[337] & b[155])^(a[336] & b[156])^(a[335] & b[157])^(a[334] & b[158])^(a[333] & b[159])^(a[332] & b[160])^(a[331] & b[161])^(a[330] & b[162])^(a[329] & b[163])^(a[328] & b[164])^(a[327] & b[165])^(a[326] & b[166])^(a[325] & b[167])^(a[324] & b[168])^(a[323] & b[169])^(a[322] & b[170])^(a[321] & b[171])^(a[320] & b[172])^(a[319] & b[173])^(a[318] & b[174])^(a[317] & b[175])^(a[316] & b[176])^(a[315] & b[177])^(a[314] & b[178])^(a[313] & b[179])^(a[312] & b[180])^(a[311] & b[181])^(a[310] & b[182])^(a[309] & b[183])^(a[308] & b[184])^(a[307] & b[185])^(a[306] & b[186])^(a[305] & b[187])^(a[304] & b[188])^(a[303] & b[189])^(a[302] & b[190])^(a[301] & b[191])^(a[300] & b[192])^(a[299] & b[193])^(a[298] & b[194])^(a[297] & b[195])^(a[296] & b[196])^(a[295] & b[197])^(a[294] & b[198])^(a[293] & b[199])^(a[292] & b[200])^(a[291] & b[201])^(a[290] & b[202])^(a[289] & b[203])^(a[288] & b[204])^(a[287] & b[205])^(a[286] & b[206])^(a[285] & b[207])^(a[284] & b[208])^(a[283] & b[209])^(a[282] & b[210])^(a[281] & b[211])^(a[280] & b[212])^(a[279] & b[213])^(a[278] & b[214])^(a[277] & b[215])^(a[276] & b[216])^(a[275] & b[217])^(a[274] & b[218])^(a[273] & b[219])^(a[272] & b[220])^(a[271] & b[221])^(a[270] & b[222])^(a[269] & b[223])^(a[268] & b[224])^(a[267] & b[225])^(a[266] & b[226])^(a[265] & b[227])^(a[264] & b[228])^(a[263] & b[229])^(a[262] & b[230])^(a[261] & b[231])^(a[260] & b[232])^(a[259] & b[233])^(a[258] & b[234])^(a[257] & b[235])^(a[256] & b[236])^(a[255] & b[237])^(a[254] & b[238])^(a[253] & b[239])^(a[252] & b[240])^(a[251] & b[241])^(a[250] & b[242])^(a[249] & b[243])^(a[248] & b[244])^(a[247] & b[245])^(a[246] & b[246])^(a[245] & b[247])^(a[244] & b[248])^(a[243] & b[249])^(a[242] & b[250])^(a[241] & b[251])^(a[240] & b[252])^(a[239] & b[253])^(a[238] & b[254])^(a[237] & b[255])^(a[236] & b[256])^(a[235] & b[257])^(a[234] & b[258])^(a[233] & b[259])^(a[232] & b[260])^(a[231] & b[261])^(a[230] & b[262])^(a[229] & b[263])^(a[228] & b[264])^(a[227] & b[265])^(a[226] & b[266])^(a[225] & b[267])^(a[224] & b[268])^(a[223] & b[269])^(a[222] & b[270])^(a[221] & b[271])^(a[220] & b[272])^(a[219] & b[273])^(a[218] & b[274])^(a[217] & b[275])^(a[216] & b[276])^(a[215] & b[277])^(a[214] & b[278])^(a[213] & b[279])^(a[212] & b[280])^(a[211] & b[281])^(a[210] & b[282])^(a[209] & b[283])^(a[208] & b[284])^(a[207] & b[285])^(a[206] & b[286])^(a[205] & b[287])^(a[204] & b[288])^(a[203] & b[289])^(a[202] & b[290])^(a[201] & b[291])^(a[200] & b[292])^(a[199] & b[293])^(a[198] & b[294])^(a[197] & b[295])^(a[196] & b[296])^(a[195] & b[297])^(a[194] & b[298])^(a[193] & b[299])^(a[192] & b[300])^(a[191] & b[301])^(a[190] & b[302])^(a[189] & b[303])^(a[188] & b[304])^(a[187] & b[305])^(a[186] & b[306])^(a[185] & b[307])^(a[184] & b[308])^(a[183] & b[309])^(a[182] & b[310])^(a[181] & b[311])^(a[180] & b[312])^(a[179] & b[313])^(a[178] & b[314])^(a[177] & b[315])^(a[176] & b[316])^(a[175] & b[317])^(a[174] & b[318])^(a[173] & b[319])^(a[172] & b[320])^(a[171] & b[321])^(a[170] & b[322])^(a[169] & b[323])^(a[168] & b[324])^(a[167] & b[325])^(a[166] & b[326])^(a[165] & b[327])^(a[164] & b[328])^(a[163] & b[329])^(a[162] & b[330])^(a[161] & b[331])^(a[160] & b[332])^(a[159] & b[333])^(a[158] & b[334])^(a[157] & b[335])^(a[156] & b[336])^(a[155] & b[337])^(a[154] & b[338])^(a[153] & b[339])^(a[152] & b[340])^(a[151] & b[341])^(a[150] & b[342])^(a[149] & b[343])^(a[148] & b[344])^(a[147] & b[345])^(a[146] & b[346])^(a[145] & b[347])^(a[144] & b[348])^(a[143] & b[349])^(a[142] & b[350])^(a[141] & b[351])^(a[140] & b[352])^(a[139] & b[353])^(a[138] & b[354])^(a[137] & b[355])^(a[136] & b[356])^(a[135] & b[357])^(a[134] & b[358])^(a[133] & b[359])^(a[132] & b[360])^(a[131] & b[361])^(a[130] & b[362])^(a[129] & b[363])^(a[128] & b[364])^(a[127] & b[365])^(a[126] & b[366])^(a[125] & b[367])^(a[124] & b[368])^(a[123] & b[369])^(a[122] & b[370])^(a[121] & b[371])^(a[120] & b[372])^(a[119] & b[373])^(a[118] & b[374])^(a[117] & b[375])^(a[116] & b[376])^(a[115] & b[377])^(a[114] & b[378])^(a[113] & b[379])^(a[112] & b[380])^(a[111] & b[381])^(a[110] & b[382])^(a[109] & b[383])^(a[108] & b[384])^(a[107] & b[385])^(a[106] & b[386])^(a[105] & b[387])^(a[104] & b[388])^(a[103] & b[389])^(a[102] & b[390])^(a[101] & b[391])^(a[100] & b[392])^(a[99] & b[393])^(a[98] & b[394])^(a[97] & b[395])^(a[96] & b[396])^(a[95] & b[397])^(a[94] & b[398])^(a[93] & b[399])^(a[92] & b[400])^(a[91] & b[401])^(a[90] & b[402])^(a[89] & b[403])^(a[88] & b[404])^(a[87] & b[405])^(a[86] & b[406])^(a[85] & b[407])^(a[84] & b[408]);
assign y[493] = (a[408] & b[85])^(a[407] & b[86])^(a[406] & b[87])^(a[405] & b[88])^(a[404] & b[89])^(a[403] & b[90])^(a[402] & b[91])^(a[401] & b[92])^(a[400] & b[93])^(a[399] & b[94])^(a[398] & b[95])^(a[397] & b[96])^(a[396] & b[97])^(a[395] & b[98])^(a[394] & b[99])^(a[393] & b[100])^(a[392] & b[101])^(a[391] & b[102])^(a[390] & b[103])^(a[389] & b[104])^(a[388] & b[105])^(a[387] & b[106])^(a[386] & b[107])^(a[385] & b[108])^(a[384] & b[109])^(a[383] & b[110])^(a[382] & b[111])^(a[381] & b[112])^(a[380] & b[113])^(a[379] & b[114])^(a[378] & b[115])^(a[377] & b[116])^(a[376] & b[117])^(a[375] & b[118])^(a[374] & b[119])^(a[373] & b[120])^(a[372] & b[121])^(a[371] & b[122])^(a[370] & b[123])^(a[369] & b[124])^(a[368] & b[125])^(a[367] & b[126])^(a[366] & b[127])^(a[365] & b[128])^(a[364] & b[129])^(a[363] & b[130])^(a[362] & b[131])^(a[361] & b[132])^(a[360] & b[133])^(a[359] & b[134])^(a[358] & b[135])^(a[357] & b[136])^(a[356] & b[137])^(a[355] & b[138])^(a[354] & b[139])^(a[353] & b[140])^(a[352] & b[141])^(a[351] & b[142])^(a[350] & b[143])^(a[349] & b[144])^(a[348] & b[145])^(a[347] & b[146])^(a[346] & b[147])^(a[345] & b[148])^(a[344] & b[149])^(a[343] & b[150])^(a[342] & b[151])^(a[341] & b[152])^(a[340] & b[153])^(a[339] & b[154])^(a[338] & b[155])^(a[337] & b[156])^(a[336] & b[157])^(a[335] & b[158])^(a[334] & b[159])^(a[333] & b[160])^(a[332] & b[161])^(a[331] & b[162])^(a[330] & b[163])^(a[329] & b[164])^(a[328] & b[165])^(a[327] & b[166])^(a[326] & b[167])^(a[325] & b[168])^(a[324] & b[169])^(a[323] & b[170])^(a[322] & b[171])^(a[321] & b[172])^(a[320] & b[173])^(a[319] & b[174])^(a[318] & b[175])^(a[317] & b[176])^(a[316] & b[177])^(a[315] & b[178])^(a[314] & b[179])^(a[313] & b[180])^(a[312] & b[181])^(a[311] & b[182])^(a[310] & b[183])^(a[309] & b[184])^(a[308] & b[185])^(a[307] & b[186])^(a[306] & b[187])^(a[305] & b[188])^(a[304] & b[189])^(a[303] & b[190])^(a[302] & b[191])^(a[301] & b[192])^(a[300] & b[193])^(a[299] & b[194])^(a[298] & b[195])^(a[297] & b[196])^(a[296] & b[197])^(a[295] & b[198])^(a[294] & b[199])^(a[293] & b[200])^(a[292] & b[201])^(a[291] & b[202])^(a[290] & b[203])^(a[289] & b[204])^(a[288] & b[205])^(a[287] & b[206])^(a[286] & b[207])^(a[285] & b[208])^(a[284] & b[209])^(a[283] & b[210])^(a[282] & b[211])^(a[281] & b[212])^(a[280] & b[213])^(a[279] & b[214])^(a[278] & b[215])^(a[277] & b[216])^(a[276] & b[217])^(a[275] & b[218])^(a[274] & b[219])^(a[273] & b[220])^(a[272] & b[221])^(a[271] & b[222])^(a[270] & b[223])^(a[269] & b[224])^(a[268] & b[225])^(a[267] & b[226])^(a[266] & b[227])^(a[265] & b[228])^(a[264] & b[229])^(a[263] & b[230])^(a[262] & b[231])^(a[261] & b[232])^(a[260] & b[233])^(a[259] & b[234])^(a[258] & b[235])^(a[257] & b[236])^(a[256] & b[237])^(a[255] & b[238])^(a[254] & b[239])^(a[253] & b[240])^(a[252] & b[241])^(a[251] & b[242])^(a[250] & b[243])^(a[249] & b[244])^(a[248] & b[245])^(a[247] & b[246])^(a[246] & b[247])^(a[245] & b[248])^(a[244] & b[249])^(a[243] & b[250])^(a[242] & b[251])^(a[241] & b[252])^(a[240] & b[253])^(a[239] & b[254])^(a[238] & b[255])^(a[237] & b[256])^(a[236] & b[257])^(a[235] & b[258])^(a[234] & b[259])^(a[233] & b[260])^(a[232] & b[261])^(a[231] & b[262])^(a[230] & b[263])^(a[229] & b[264])^(a[228] & b[265])^(a[227] & b[266])^(a[226] & b[267])^(a[225] & b[268])^(a[224] & b[269])^(a[223] & b[270])^(a[222] & b[271])^(a[221] & b[272])^(a[220] & b[273])^(a[219] & b[274])^(a[218] & b[275])^(a[217] & b[276])^(a[216] & b[277])^(a[215] & b[278])^(a[214] & b[279])^(a[213] & b[280])^(a[212] & b[281])^(a[211] & b[282])^(a[210] & b[283])^(a[209] & b[284])^(a[208] & b[285])^(a[207] & b[286])^(a[206] & b[287])^(a[205] & b[288])^(a[204] & b[289])^(a[203] & b[290])^(a[202] & b[291])^(a[201] & b[292])^(a[200] & b[293])^(a[199] & b[294])^(a[198] & b[295])^(a[197] & b[296])^(a[196] & b[297])^(a[195] & b[298])^(a[194] & b[299])^(a[193] & b[300])^(a[192] & b[301])^(a[191] & b[302])^(a[190] & b[303])^(a[189] & b[304])^(a[188] & b[305])^(a[187] & b[306])^(a[186] & b[307])^(a[185] & b[308])^(a[184] & b[309])^(a[183] & b[310])^(a[182] & b[311])^(a[181] & b[312])^(a[180] & b[313])^(a[179] & b[314])^(a[178] & b[315])^(a[177] & b[316])^(a[176] & b[317])^(a[175] & b[318])^(a[174] & b[319])^(a[173] & b[320])^(a[172] & b[321])^(a[171] & b[322])^(a[170] & b[323])^(a[169] & b[324])^(a[168] & b[325])^(a[167] & b[326])^(a[166] & b[327])^(a[165] & b[328])^(a[164] & b[329])^(a[163] & b[330])^(a[162] & b[331])^(a[161] & b[332])^(a[160] & b[333])^(a[159] & b[334])^(a[158] & b[335])^(a[157] & b[336])^(a[156] & b[337])^(a[155] & b[338])^(a[154] & b[339])^(a[153] & b[340])^(a[152] & b[341])^(a[151] & b[342])^(a[150] & b[343])^(a[149] & b[344])^(a[148] & b[345])^(a[147] & b[346])^(a[146] & b[347])^(a[145] & b[348])^(a[144] & b[349])^(a[143] & b[350])^(a[142] & b[351])^(a[141] & b[352])^(a[140] & b[353])^(a[139] & b[354])^(a[138] & b[355])^(a[137] & b[356])^(a[136] & b[357])^(a[135] & b[358])^(a[134] & b[359])^(a[133] & b[360])^(a[132] & b[361])^(a[131] & b[362])^(a[130] & b[363])^(a[129] & b[364])^(a[128] & b[365])^(a[127] & b[366])^(a[126] & b[367])^(a[125] & b[368])^(a[124] & b[369])^(a[123] & b[370])^(a[122] & b[371])^(a[121] & b[372])^(a[120] & b[373])^(a[119] & b[374])^(a[118] & b[375])^(a[117] & b[376])^(a[116] & b[377])^(a[115] & b[378])^(a[114] & b[379])^(a[113] & b[380])^(a[112] & b[381])^(a[111] & b[382])^(a[110] & b[383])^(a[109] & b[384])^(a[108] & b[385])^(a[107] & b[386])^(a[106] & b[387])^(a[105] & b[388])^(a[104] & b[389])^(a[103] & b[390])^(a[102] & b[391])^(a[101] & b[392])^(a[100] & b[393])^(a[99] & b[394])^(a[98] & b[395])^(a[97] & b[396])^(a[96] & b[397])^(a[95] & b[398])^(a[94] & b[399])^(a[93] & b[400])^(a[92] & b[401])^(a[91] & b[402])^(a[90] & b[403])^(a[89] & b[404])^(a[88] & b[405])^(a[87] & b[406])^(a[86] & b[407])^(a[85] & b[408]);
assign y[494] = (a[408] & b[86])^(a[407] & b[87])^(a[406] & b[88])^(a[405] & b[89])^(a[404] & b[90])^(a[403] & b[91])^(a[402] & b[92])^(a[401] & b[93])^(a[400] & b[94])^(a[399] & b[95])^(a[398] & b[96])^(a[397] & b[97])^(a[396] & b[98])^(a[395] & b[99])^(a[394] & b[100])^(a[393] & b[101])^(a[392] & b[102])^(a[391] & b[103])^(a[390] & b[104])^(a[389] & b[105])^(a[388] & b[106])^(a[387] & b[107])^(a[386] & b[108])^(a[385] & b[109])^(a[384] & b[110])^(a[383] & b[111])^(a[382] & b[112])^(a[381] & b[113])^(a[380] & b[114])^(a[379] & b[115])^(a[378] & b[116])^(a[377] & b[117])^(a[376] & b[118])^(a[375] & b[119])^(a[374] & b[120])^(a[373] & b[121])^(a[372] & b[122])^(a[371] & b[123])^(a[370] & b[124])^(a[369] & b[125])^(a[368] & b[126])^(a[367] & b[127])^(a[366] & b[128])^(a[365] & b[129])^(a[364] & b[130])^(a[363] & b[131])^(a[362] & b[132])^(a[361] & b[133])^(a[360] & b[134])^(a[359] & b[135])^(a[358] & b[136])^(a[357] & b[137])^(a[356] & b[138])^(a[355] & b[139])^(a[354] & b[140])^(a[353] & b[141])^(a[352] & b[142])^(a[351] & b[143])^(a[350] & b[144])^(a[349] & b[145])^(a[348] & b[146])^(a[347] & b[147])^(a[346] & b[148])^(a[345] & b[149])^(a[344] & b[150])^(a[343] & b[151])^(a[342] & b[152])^(a[341] & b[153])^(a[340] & b[154])^(a[339] & b[155])^(a[338] & b[156])^(a[337] & b[157])^(a[336] & b[158])^(a[335] & b[159])^(a[334] & b[160])^(a[333] & b[161])^(a[332] & b[162])^(a[331] & b[163])^(a[330] & b[164])^(a[329] & b[165])^(a[328] & b[166])^(a[327] & b[167])^(a[326] & b[168])^(a[325] & b[169])^(a[324] & b[170])^(a[323] & b[171])^(a[322] & b[172])^(a[321] & b[173])^(a[320] & b[174])^(a[319] & b[175])^(a[318] & b[176])^(a[317] & b[177])^(a[316] & b[178])^(a[315] & b[179])^(a[314] & b[180])^(a[313] & b[181])^(a[312] & b[182])^(a[311] & b[183])^(a[310] & b[184])^(a[309] & b[185])^(a[308] & b[186])^(a[307] & b[187])^(a[306] & b[188])^(a[305] & b[189])^(a[304] & b[190])^(a[303] & b[191])^(a[302] & b[192])^(a[301] & b[193])^(a[300] & b[194])^(a[299] & b[195])^(a[298] & b[196])^(a[297] & b[197])^(a[296] & b[198])^(a[295] & b[199])^(a[294] & b[200])^(a[293] & b[201])^(a[292] & b[202])^(a[291] & b[203])^(a[290] & b[204])^(a[289] & b[205])^(a[288] & b[206])^(a[287] & b[207])^(a[286] & b[208])^(a[285] & b[209])^(a[284] & b[210])^(a[283] & b[211])^(a[282] & b[212])^(a[281] & b[213])^(a[280] & b[214])^(a[279] & b[215])^(a[278] & b[216])^(a[277] & b[217])^(a[276] & b[218])^(a[275] & b[219])^(a[274] & b[220])^(a[273] & b[221])^(a[272] & b[222])^(a[271] & b[223])^(a[270] & b[224])^(a[269] & b[225])^(a[268] & b[226])^(a[267] & b[227])^(a[266] & b[228])^(a[265] & b[229])^(a[264] & b[230])^(a[263] & b[231])^(a[262] & b[232])^(a[261] & b[233])^(a[260] & b[234])^(a[259] & b[235])^(a[258] & b[236])^(a[257] & b[237])^(a[256] & b[238])^(a[255] & b[239])^(a[254] & b[240])^(a[253] & b[241])^(a[252] & b[242])^(a[251] & b[243])^(a[250] & b[244])^(a[249] & b[245])^(a[248] & b[246])^(a[247] & b[247])^(a[246] & b[248])^(a[245] & b[249])^(a[244] & b[250])^(a[243] & b[251])^(a[242] & b[252])^(a[241] & b[253])^(a[240] & b[254])^(a[239] & b[255])^(a[238] & b[256])^(a[237] & b[257])^(a[236] & b[258])^(a[235] & b[259])^(a[234] & b[260])^(a[233] & b[261])^(a[232] & b[262])^(a[231] & b[263])^(a[230] & b[264])^(a[229] & b[265])^(a[228] & b[266])^(a[227] & b[267])^(a[226] & b[268])^(a[225] & b[269])^(a[224] & b[270])^(a[223] & b[271])^(a[222] & b[272])^(a[221] & b[273])^(a[220] & b[274])^(a[219] & b[275])^(a[218] & b[276])^(a[217] & b[277])^(a[216] & b[278])^(a[215] & b[279])^(a[214] & b[280])^(a[213] & b[281])^(a[212] & b[282])^(a[211] & b[283])^(a[210] & b[284])^(a[209] & b[285])^(a[208] & b[286])^(a[207] & b[287])^(a[206] & b[288])^(a[205] & b[289])^(a[204] & b[290])^(a[203] & b[291])^(a[202] & b[292])^(a[201] & b[293])^(a[200] & b[294])^(a[199] & b[295])^(a[198] & b[296])^(a[197] & b[297])^(a[196] & b[298])^(a[195] & b[299])^(a[194] & b[300])^(a[193] & b[301])^(a[192] & b[302])^(a[191] & b[303])^(a[190] & b[304])^(a[189] & b[305])^(a[188] & b[306])^(a[187] & b[307])^(a[186] & b[308])^(a[185] & b[309])^(a[184] & b[310])^(a[183] & b[311])^(a[182] & b[312])^(a[181] & b[313])^(a[180] & b[314])^(a[179] & b[315])^(a[178] & b[316])^(a[177] & b[317])^(a[176] & b[318])^(a[175] & b[319])^(a[174] & b[320])^(a[173] & b[321])^(a[172] & b[322])^(a[171] & b[323])^(a[170] & b[324])^(a[169] & b[325])^(a[168] & b[326])^(a[167] & b[327])^(a[166] & b[328])^(a[165] & b[329])^(a[164] & b[330])^(a[163] & b[331])^(a[162] & b[332])^(a[161] & b[333])^(a[160] & b[334])^(a[159] & b[335])^(a[158] & b[336])^(a[157] & b[337])^(a[156] & b[338])^(a[155] & b[339])^(a[154] & b[340])^(a[153] & b[341])^(a[152] & b[342])^(a[151] & b[343])^(a[150] & b[344])^(a[149] & b[345])^(a[148] & b[346])^(a[147] & b[347])^(a[146] & b[348])^(a[145] & b[349])^(a[144] & b[350])^(a[143] & b[351])^(a[142] & b[352])^(a[141] & b[353])^(a[140] & b[354])^(a[139] & b[355])^(a[138] & b[356])^(a[137] & b[357])^(a[136] & b[358])^(a[135] & b[359])^(a[134] & b[360])^(a[133] & b[361])^(a[132] & b[362])^(a[131] & b[363])^(a[130] & b[364])^(a[129] & b[365])^(a[128] & b[366])^(a[127] & b[367])^(a[126] & b[368])^(a[125] & b[369])^(a[124] & b[370])^(a[123] & b[371])^(a[122] & b[372])^(a[121] & b[373])^(a[120] & b[374])^(a[119] & b[375])^(a[118] & b[376])^(a[117] & b[377])^(a[116] & b[378])^(a[115] & b[379])^(a[114] & b[380])^(a[113] & b[381])^(a[112] & b[382])^(a[111] & b[383])^(a[110] & b[384])^(a[109] & b[385])^(a[108] & b[386])^(a[107] & b[387])^(a[106] & b[388])^(a[105] & b[389])^(a[104] & b[390])^(a[103] & b[391])^(a[102] & b[392])^(a[101] & b[393])^(a[100] & b[394])^(a[99] & b[395])^(a[98] & b[396])^(a[97] & b[397])^(a[96] & b[398])^(a[95] & b[399])^(a[94] & b[400])^(a[93] & b[401])^(a[92] & b[402])^(a[91] & b[403])^(a[90] & b[404])^(a[89] & b[405])^(a[88] & b[406])^(a[87] & b[407])^(a[86] & b[408]);
assign y[495] = (a[408] & b[87])^(a[407] & b[88])^(a[406] & b[89])^(a[405] & b[90])^(a[404] & b[91])^(a[403] & b[92])^(a[402] & b[93])^(a[401] & b[94])^(a[400] & b[95])^(a[399] & b[96])^(a[398] & b[97])^(a[397] & b[98])^(a[396] & b[99])^(a[395] & b[100])^(a[394] & b[101])^(a[393] & b[102])^(a[392] & b[103])^(a[391] & b[104])^(a[390] & b[105])^(a[389] & b[106])^(a[388] & b[107])^(a[387] & b[108])^(a[386] & b[109])^(a[385] & b[110])^(a[384] & b[111])^(a[383] & b[112])^(a[382] & b[113])^(a[381] & b[114])^(a[380] & b[115])^(a[379] & b[116])^(a[378] & b[117])^(a[377] & b[118])^(a[376] & b[119])^(a[375] & b[120])^(a[374] & b[121])^(a[373] & b[122])^(a[372] & b[123])^(a[371] & b[124])^(a[370] & b[125])^(a[369] & b[126])^(a[368] & b[127])^(a[367] & b[128])^(a[366] & b[129])^(a[365] & b[130])^(a[364] & b[131])^(a[363] & b[132])^(a[362] & b[133])^(a[361] & b[134])^(a[360] & b[135])^(a[359] & b[136])^(a[358] & b[137])^(a[357] & b[138])^(a[356] & b[139])^(a[355] & b[140])^(a[354] & b[141])^(a[353] & b[142])^(a[352] & b[143])^(a[351] & b[144])^(a[350] & b[145])^(a[349] & b[146])^(a[348] & b[147])^(a[347] & b[148])^(a[346] & b[149])^(a[345] & b[150])^(a[344] & b[151])^(a[343] & b[152])^(a[342] & b[153])^(a[341] & b[154])^(a[340] & b[155])^(a[339] & b[156])^(a[338] & b[157])^(a[337] & b[158])^(a[336] & b[159])^(a[335] & b[160])^(a[334] & b[161])^(a[333] & b[162])^(a[332] & b[163])^(a[331] & b[164])^(a[330] & b[165])^(a[329] & b[166])^(a[328] & b[167])^(a[327] & b[168])^(a[326] & b[169])^(a[325] & b[170])^(a[324] & b[171])^(a[323] & b[172])^(a[322] & b[173])^(a[321] & b[174])^(a[320] & b[175])^(a[319] & b[176])^(a[318] & b[177])^(a[317] & b[178])^(a[316] & b[179])^(a[315] & b[180])^(a[314] & b[181])^(a[313] & b[182])^(a[312] & b[183])^(a[311] & b[184])^(a[310] & b[185])^(a[309] & b[186])^(a[308] & b[187])^(a[307] & b[188])^(a[306] & b[189])^(a[305] & b[190])^(a[304] & b[191])^(a[303] & b[192])^(a[302] & b[193])^(a[301] & b[194])^(a[300] & b[195])^(a[299] & b[196])^(a[298] & b[197])^(a[297] & b[198])^(a[296] & b[199])^(a[295] & b[200])^(a[294] & b[201])^(a[293] & b[202])^(a[292] & b[203])^(a[291] & b[204])^(a[290] & b[205])^(a[289] & b[206])^(a[288] & b[207])^(a[287] & b[208])^(a[286] & b[209])^(a[285] & b[210])^(a[284] & b[211])^(a[283] & b[212])^(a[282] & b[213])^(a[281] & b[214])^(a[280] & b[215])^(a[279] & b[216])^(a[278] & b[217])^(a[277] & b[218])^(a[276] & b[219])^(a[275] & b[220])^(a[274] & b[221])^(a[273] & b[222])^(a[272] & b[223])^(a[271] & b[224])^(a[270] & b[225])^(a[269] & b[226])^(a[268] & b[227])^(a[267] & b[228])^(a[266] & b[229])^(a[265] & b[230])^(a[264] & b[231])^(a[263] & b[232])^(a[262] & b[233])^(a[261] & b[234])^(a[260] & b[235])^(a[259] & b[236])^(a[258] & b[237])^(a[257] & b[238])^(a[256] & b[239])^(a[255] & b[240])^(a[254] & b[241])^(a[253] & b[242])^(a[252] & b[243])^(a[251] & b[244])^(a[250] & b[245])^(a[249] & b[246])^(a[248] & b[247])^(a[247] & b[248])^(a[246] & b[249])^(a[245] & b[250])^(a[244] & b[251])^(a[243] & b[252])^(a[242] & b[253])^(a[241] & b[254])^(a[240] & b[255])^(a[239] & b[256])^(a[238] & b[257])^(a[237] & b[258])^(a[236] & b[259])^(a[235] & b[260])^(a[234] & b[261])^(a[233] & b[262])^(a[232] & b[263])^(a[231] & b[264])^(a[230] & b[265])^(a[229] & b[266])^(a[228] & b[267])^(a[227] & b[268])^(a[226] & b[269])^(a[225] & b[270])^(a[224] & b[271])^(a[223] & b[272])^(a[222] & b[273])^(a[221] & b[274])^(a[220] & b[275])^(a[219] & b[276])^(a[218] & b[277])^(a[217] & b[278])^(a[216] & b[279])^(a[215] & b[280])^(a[214] & b[281])^(a[213] & b[282])^(a[212] & b[283])^(a[211] & b[284])^(a[210] & b[285])^(a[209] & b[286])^(a[208] & b[287])^(a[207] & b[288])^(a[206] & b[289])^(a[205] & b[290])^(a[204] & b[291])^(a[203] & b[292])^(a[202] & b[293])^(a[201] & b[294])^(a[200] & b[295])^(a[199] & b[296])^(a[198] & b[297])^(a[197] & b[298])^(a[196] & b[299])^(a[195] & b[300])^(a[194] & b[301])^(a[193] & b[302])^(a[192] & b[303])^(a[191] & b[304])^(a[190] & b[305])^(a[189] & b[306])^(a[188] & b[307])^(a[187] & b[308])^(a[186] & b[309])^(a[185] & b[310])^(a[184] & b[311])^(a[183] & b[312])^(a[182] & b[313])^(a[181] & b[314])^(a[180] & b[315])^(a[179] & b[316])^(a[178] & b[317])^(a[177] & b[318])^(a[176] & b[319])^(a[175] & b[320])^(a[174] & b[321])^(a[173] & b[322])^(a[172] & b[323])^(a[171] & b[324])^(a[170] & b[325])^(a[169] & b[326])^(a[168] & b[327])^(a[167] & b[328])^(a[166] & b[329])^(a[165] & b[330])^(a[164] & b[331])^(a[163] & b[332])^(a[162] & b[333])^(a[161] & b[334])^(a[160] & b[335])^(a[159] & b[336])^(a[158] & b[337])^(a[157] & b[338])^(a[156] & b[339])^(a[155] & b[340])^(a[154] & b[341])^(a[153] & b[342])^(a[152] & b[343])^(a[151] & b[344])^(a[150] & b[345])^(a[149] & b[346])^(a[148] & b[347])^(a[147] & b[348])^(a[146] & b[349])^(a[145] & b[350])^(a[144] & b[351])^(a[143] & b[352])^(a[142] & b[353])^(a[141] & b[354])^(a[140] & b[355])^(a[139] & b[356])^(a[138] & b[357])^(a[137] & b[358])^(a[136] & b[359])^(a[135] & b[360])^(a[134] & b[361])^(a[133] & b[362])^(a[132] & b[363])^(a[131] & b[364])^(a[130] & b[365])^(a[129] & b[366])^(a[128] & b[367])^(a[127] & b[368])^(a[126] & b[369])^(a[125] & b[370])^(a[124] & b[371])^(a[123] & b[372])^(a[122] & b[373])^(a[121] & b[374])^(a[120] & b[375])^(a[119] & b[376])^(a[118] & b[377])^(a[117] & b[378])^(a[116] & b[379])^(a[115] & b[380])^(a[114] & b[381])^(a[113] & b[382])^(a[112] & b[383])^(a[111] & b[384])^(a[110] & b[385])^(a[109] & b[386])^(a[108] & b[387])^(a[107] & b[388])^(a[106] & b[389])^(a[105] & b[390])^(a[104] & b[391])^(a[103] & b[392])^(a[102] & b[393])^(a[101] & b[394])^(a[100] & b[395])^(a[99] & b[396])^(a[98] & b[397])^(a[97] & b[398])^(a[96] & b[399])^(a[95] & b[400])^(a[94] & b[401])^(a[93] & b[402])^(a[92] & b[403])^(a[91] & b[404])^(a[90] & b[405])^(a[89] & b[406])^(a[88] & b[407])^(a[87] & b[408]);
assign y[496] = (a[408] & b[88])^(a[407] & b[89])^(a[406] & b[90])^(a[405] & b[91])^(a[404] & b[92])^(a[403] & b[93])^(a[402] & b[94])^(a[401] & b[95])^(a[400] & b[96])^(a[399] & b[97])^(a[398] & b[98])^(a[397] & b[99])^(a[396] & b[100])^(a[395] & b[101])^(a[394] & b[102])^(a[393] & b[103])^(a[392] & b[104])^(a[391] & b[105])^(a[390] & b[106])^(a[389] & b[107])^(a[388] & b[108])^(a[387] & b[109])^(a[386] & b[110])^(a[385] & b[111])^(a[384] & b[112])^(a[383] & b[113])^(a[382] & b[114])^(a[381] & b[115])^(a[380] & b[116])^(a[379] & b[117])^(a[378] & b[118])^(a[377] & b[119])^(a[376] & b[120])^(a[375] & b[121])^(a[374] & b[122])^(a[373] & b[123])^(a[372] & b[124])^(a[371] & b[125])^(a[370] & b[126])^(a[369] & b[127])^(a[368] & b[128])^(a[367] & b[129])^(a[366] & b[130])^(a[365] & b[131])^(a[364] & b[132])^(a[363] & b[133])^(a[362] & b[134])^(a[361] & b[135])^(a[360] & b[136])^(a[359] & b[137])^(a[358] & b[138])^(a[357] & b[139])^(a[356] & b[140])^(a[355] & b[141])^(a[354] & b[142])^(a[353] & b[143])^(a[352] & b[144])^(a[351] & b[145])^(a[350] & b[146])^(a[349] & b[147])^(a[348] & b[148])^(a[347] & b[149])^(a[346] & b[150])^(a[345] & b[151])^(a[344] & b[152])^(a[343] & b[153])^(a[342] & b[154])^(a[341] & b[155])^(a[340] & b[156])^(a[339] & b[157])^(a[338] & b[158])^(a[337] & b[159])^(a[336] & b[160])^(a[335] & b[161])^(a[334] & b[162])^(a[333] & b[163])^(a[332] & b[164])^(a[331] & b[165])^(a[330] & b[166])^(a[329] & b[167])^(a[328] & b[168])^(a[327] & b[169])^(a[326] & b[170])^(a[325] & b[171])^(a[324] & b[172])^(a[323] & b[173])^(a[322] & b[174])^(a[321] & b[175])^(a[320] & b[176])^(a[319] & b[177])^(a[318] & b[178])^(a[317] & b[179])^(a[316] & b[180])^(a[315] & b[181])^(a[314] & b[182])^(a[313] & b[183])^(a[312] & b[184])^(a[311] & b[185])^(a[310] & b[186])^(a[309] & b[187])^(a[308] & b[188])^(a[307] & b[189])^(a[306] & b[190])^(a[305] & b[191])^(a[304] & b[192])^(a[303] & b[193])^(a[302] & b[194])^(a[301] & b[195])^(a[300] & b[196])^(a[299] & b[197])^(a[298] & b[198])^(a[297] & b[199])^(a[296] & b[200])^(a[295] & b[201])^(a[294] & b[202])^(a[293] & b[203])^(a[292] & b[204])^(a[291] & b[205])^(a[290] & b[206])^(a[289] & b[207])^(a[288] & b[208])^(a[287] & b[209])^(a[286] & b[210])^(a[285] & b[211])^(a[284] & b[212])^(a[283] & b[213])^(a[282] & b[214])^(a[281] & b[215])^(a[280] & b[216])^(a[279] & b[217])^(a[278] & b[218])^(a[277] & b[219])^(a[276] & b[220])^(a[275] & b[221])^(a[274] & b[222])^(a[273] & b[223])^(a[272] & b[224])^(a[271] & b[225])^(a[270] & b[226])^(a[269] & b[227])^(a[268] & b[228])^(a[267] & b[229])^(a[266] & b[230])^(a[265] & b[231])^(a[264] & b[232])^(a[263] & b[233])^(a[262] & b[234])^(a[261] & b[235])^(a[260] & b[236])^(a[259] & b[237])^(a[258] & b[238])^(a[257] & b[239])^(a[256] & b[240])^(a[255] & b[241])^(a[254] & b[242])^(a[253] & b[243])^(a[252] & b[244])^(a[251] & b[245])^(a[250] & b[246])^(a[249] & b[247])^(a[248] & b[248])^(a[247] & b[249])^(a[246] & b[250])^(a[245] & b[251])^(a[244] & b[252])^(a[243] & b[253])^(a[242] & b[254])^(a[241] & b[255])^(a[240] & b[256])^(a[239] & b[257])^(a[238] & b[258])^(a[237] & b[259])^(a[236] & b[260])^(a[235] & b[261])^(a[234] & b[262])^(a[233] & b[263])^(a[232] & b[264])^(a[231] & b[265])^(a[230] & b[266])^(a[229] & b[267])^(a[228] & b[268])^(a[227] & b[269])^(a[226] & b[270])^(a[225] & b[271])^(a[224] & b[272])^(a[223] & b[273])^(a[222] & b[274])^(a[221] & b[275])^(a[220] & b[276])^(a[219] & b[277])^(a[218] & b[278])^(a[217] & b[279])^(a[216] & b[280])^(a[215] & b[281])^(a[214] & b[282])^(a[213] & b[283])^(a[212] & b[284])^(a[211] & b[285])^(a[210] & b[286])^(a[209] & b[287])^(a[208] & b[288])^(a[207] & b[289])^(a[206] & b[290])^(a[205] & b[291])^(a[204] & b[292])^(a[203] & b[293])^(a[202] & b[294])^(a[201] & b[295])^(a[200] & b[296])^(a[199] & b[297])^(a[198] & b[298])^(a[197] & b[299])^(a[196] & b[300])^(a[195] & b[301])^(a[194] & b[302])^(a[193] & b[303])^(a[192] & b[304])^(a[191] & b[305])^(a[190] & b[306])^(a[189] & b[307])^(a[188] & b[308])^(a[187] & b[309])^(a[186] & b[310])^(a[185] & b[311])^(a[184] & b[312])^(a[183] & b[313])^(a[182] & b[314])^(a[181] & b[315])^(a[180] & b[316])^(a[179] & b[317])^(a[178] & b[318])^(a[177] & b[319])^(a[176] & b[320])^(a[175] & b[321])^(a[174] & b[322])^(a[173] & b[323])^(a[172] & b[324])^(a[171] & b[325])^(a[170] & b[326])^(a[169] & b[327])^(a[168] & b[328])^(a[167] & b[329])^(a[166] & b[330])^(a[165] & b[331])^(a[164] & b[332])^(a[163] & b[333])^(a[162] & b[334])^(a[161] & b[335])^(a[160] & b[336])^(a[159] & b[337])^(a[158] & b[338])^(a[157] & b[339])^(a[156] & b[340])^(a[155] & b[341])^(a[154] & b[342])^(a[153] & b[343])^(a[152] & b[344])^(a[151] & b[345])^(a[150] & b[346])^(a[149] & b[347])^(a[148] & b[348])^(a[147] & b[349])^(a[146] & b[350])^(a[145] & b[351])^(a[144] & b[352])^(a[143] & b[353])^(a[142] & b[354])^(a[141] & b[355])^(a[140] & b[356])^(a[139] & b[357])^(a[138] & b[358])^(a[137] & b[359])^(a[136] & b[360])^(a[135] & b[361])^(a[134] & b[362])^(a[133] & b[363])^(a[132] & b[364])^(a[131] & b[365])^(a[130] & b[366])^(a[129] & b[367])^(a[128] & b[368])^(a[127] & b[369])^(a[126] & b[370])^(a[125] & b[371])^(a[124] & b[372])^(a[123] & b[373])^(a[122] & b[374])^(a[121] & b[375])^(a[120] & b[376])^(a[119] & b[377])^(a[118] & b[378])^(a[117] & b[379])^(a[116] & b[380])^(a[115] & b[381])^(a[114] & b[382])^(a[113] & b[383])^(a[112] & b[384])^(a[111] & b[385])^(a[110] & b[386])^(a[109] & b[387])^(a[108] & b[388])^(a[107] & b[389])^(a[106] & b[390])^(a[105] & b[391])^(a[104] & b[392])^(a[103] & b[393])^(a[102] & b[394])^(a[101] & b[395])^(a[100] & b[396])^(a[99] & b[397])^(a[98] & b[398])^(a[97] & b[399])^(a[96] & b[400])^(a[95] & b[401])^(a[94] & b[402])^(a[93] & b[403])^(a[92] & b[404])^(a[91] & b[405])^(a[90] & b[406])^(a[89] & b[407])^(a[88] & b[408]);
assign y[497] = (a[408] & b[89])^(a[407] & b[90])^(a[406] & b[91])^(a[405] & b[92])^(a[404] & b[93])^(a[403] & b[94])^(a[402] & b[95])^(a[401] & b[96])^(a[400] & b[97])^(a[399] & b[98])^(a[398] & b[99])^(a[397] & b[100])^(a[396] & b[101])^(a[395] & b[102])^(a[394] & b[103])^(a[393] & b[104])^(a[392] & b[105])^(a[391] & b[106])^(a[390] & b[107])^(a[389] & b[108])^(a[388] & b[109])^(a[387] & b[110])^(a[386] & b[111])^(a[385] & b[112])^(a[384] & b[113])^(a[383] & b[114])^(a[382] & b[115])^(a[381] & b[116])^(a[380] & b[117])^(a[379] & b[118])^(a[378] & b[119])^(a[377] & b[120])^(a[376] & b[121])^(a[375] & b[122])^(a[374] & b[123])^(a[373] & b[124])^(a[372] & b[125])^(a[371] & b[126])^(a[370] & b[127])^(a[369] & b[128])^(a[368] & b[129])^(a[367] & b[130])^(a[366] & b[131])^(a[365] & b[132])^(a[364] & b[133])^(a[363] & b[134])^(a[362] & b[135])^(a[361] & b[136])^(a[360] & b[137])^(a[359] & b[138])^(a[358] & b[139])^(a[357] & b[140])^(a[356] & b[141])^(a[355] & b[142])^(a[354] & b[143])^(a[353] & b[144])^(a[352] & b[145])^(a[351] & b[146])^(a[350] & b[147])^(a[349] & b[148])^(a[348] & b[149])^(a[347] & b[150])^(a[346] & b[151])^(a[345] & b[152])^(a[344] & b[153])^(a[343] & b[154])^(a[342] & b[155])^(a[341] & b[156])^(a[340] & b[157])^(a[339] & b[158])^(a[338] & b[159])^(a[337] & b[160])^(a[336] & b[161])^(a[335] & b[162])^(a[334] & b[163])^(a[333] & b[164])^(a[332] & b[165])^(a[331] & b[166])^(a[330] & b[167])^(a[329] & b[168])^(a[328] & b[169])^(a[327] & b[170])^(a[326] & b[171])^(a[325] & b[172])^(a[324] & b[173])^(a[323] & b[174])^(a[322] & b[175])^(a[321] & b[176])^(a[320] & b[177])^(a[319] & b[178])^(a[318] & b[179])^(a[317] & b[180])^(a[316] & b[181])^(a[315] & b[182])^(a[314] & b[183])^(a[313] & b[184])^(a[312] & b[185])^(a[311] & b[186])^(a[310] & b[187])^(a[309] & b[188])^(a[308] & b[189])^(a[307] & b[190])^(a[306] & b[191])^(a[305] & b[192])^(a[304] & b[193])^(a[303] & b[194])^(a[302] & b[195])^(a[301] & b[196])^(a[300] & b[197])^(a[299] & b[198])^(a[298] & b[199])^(a[297] & b[200])^(a[296] & b[201])^(a[295] & b[202])^(a[294] & b[203])^(a[293] & b[204])^(a[292] & b[205])^(a[291] & b[206])^(a[290] & b[207])^(a[289] & b[208])^(a[288] & b[209])^(a[287] & b[210])^(a[286] & b[211])^(a[285] & b[212])^(a[284] & b[213])^(a[283] & b[214])^(a[282] & b[215])^(a[281] & b[216])^(a[280] & b[217])^(a[279] & b[218])^(a[278] & b[219])^(a[277] & b[220])^(a[276] & b[221])^(a[275] & b[222])^(a[274] & b[223])^(a[273] & b[224])^(a[272] & b[225])^(a[271] & b[226])^(a[270] & b[227])^(a[269] & b[228])^(a[268] & b[229])^(a[267] & b[230])^(a[266] & b[231])^(a[265] & b[232])^(a[264] & b[233])^(a[263] & b[234])^(a[262] & b[235])^(a[261] & b[236])^(a[260] & b[237])^(a[259] & b[238])^(a[258] & b[239])^(a[257] & b[240])^(a[256] & b[241])^(a[255] & b[242])^(a[254] & b[243])^(a[253] & b[244])^(a[252] & b[245])^(a[251] & b[246])^(a[250] & b[247])^(a[249] & b[248])^(a[248] & b[249])^(a[247] & b[250])^(a[246] & b[251])^(a[245] & b[252])^(a[244] & b[253])^(a[243] & b[254])^(a[242] & b[255])^(a[241] & b[256])^(a[240] & b[257])^(a[239] & b[258])^(a[238] & b[259])^(a[237] & b[260])^(a[236] & b[261])^(a[235] & b[262])^(a[234] & b[263])^(a[233] & b[264])^(a[232] & b[265])^(a[231] & b[266])^(a[230] & b[267])^(a[229] & b[268])^(a[228] & b[269])^(a[227] & b[270])^(a[226] & b[271])^(a[225] & b[272])^(a[224] & b[273])^(a[223] & b[274])^(a[222] & b[275])^(a[221] & b[276])^(a[220] & b[277])^(a[219] & b[278])^(a[218] & b[279])^(a[217] & b[280])^(a[216] & b[281])^(a[215] & b[282])^(a[214] & b[283])^(a[213] & b[284])^(a[212] & b[285])^(a[211] & b[286])^(a[210] & b[287])^(a[209] & b[288])^(a[208] & b[289])^(a[207] & b[290])^(a[206] & b[291])^(a[205] & b[292])^(a[204] & b[293])^(a[203] & b[294])^(a[202] & b[295])^(a[201] & b[296])^(a[200] & b[297])^(a[199] & b[298])^(a[198] & b[299])^(a[197] & b[300])^(a[196] & b[301])^(a[195] & b[302])^(a[194] & b[303])^(a[193] & b[304])^(a[192] & b[305])^(a[191] & b[306])^(a[190] & b[307])^(a[189] & b[308])^(a[188] & b[309])^(a[187] & b[310])^(a[186] & b[311])^(a[185] & b[312])^(a[184] & b[313])^(a[183] & b[314])^(a[182] & b[315])^(a[181] & b[316])^(a[180] & b[317])^(a[179] & b[318])^(a[178] & b[319])^(a[177] & b[320])^(a[176] & b[321])^(a[175] & b[322])^(a[174] & b[323])^(a[173] & b[324])^(a[172] & b[325])^(a[171] & b[326])^(a[170] & b[327])^(a[169] & b[328])^(a[168] & b[329])^(a[167] & b[330])^(a[166] & b[331])^(a[165] & b[332])^(a[164] & b[333])^(a[163] & b[334])^(a[162] & b[335])^(a[161] & b[336])^(a[160] & b[337])^(a[159] & b[338])^(a[158] & b[339])^(a[157] & b[340])^(a[156] & b[341])^(a[155] & b[342])^(a[154] & b[343])^(a[153] & b[344])^(a[152] & b[345])^(a[151] & b[346])^(a[150] & b[347])^(a[149] & b[348])^(a[148] & b[349])^(a[147] & b[350])^(a[146] & b[351])^(a[145] & b[352])^(a[144] & b[353])^(a[143] & b[354])^(a[142] & b[355])^(a[141] & b[356])^(a[140] & b[357])^(a[139] & b[358])^(a[138] & b[359])^(a[137] & b[360])^(a[136] & b[361])^(a[135] & b[362])^(a[134] & b[363])^(a[133] & b[364])^(a[132] & b[365])^(a[131] & b[366])^(a[130] & b[367])^(a[129] & b[368])^(a[128] & b[369])^(a[127] & b[370])^(a[126] & b[371])^(a[125] & b[372])^(a[124] & b[373])^(a[123] & b[374])^(a[122] & b[375])^(a[121] & b[376])^(a[120] & b[377])^(a[119] & b[378])^(a[118] & b[379])^(a[117] & b[380])^(a[116] & b[381])^(a[115] & b[382])^(a[114] & b[383])^(a[113] & b[384])^(a[112] & b[385])^(a[111] & b[386])^(a[110] & b[387])^(a[109] & b[388])^(a[108] & b[389])^(a[107] & b[390])^(a[106] & b[391])^(a[105] & b[392])^(a[104] & b[393])^(a[103] & b[394])^(a[102] & b[395])^(a[101] & b[396])^(a[100] & b[397])^(a[99] & b[398])^(a[98] & b[399])^(a[97] & b[400])^(a[96] & b[401])^(a[95] & b[402])^(a[94] & b[403])^(a[93] & b[404])^(a[92] & b[405])^(a[91] & b[406])^(a[90] & b[407])^(a[89] & b[408]);
assign y[498] = (a[408] & b[90])^(a[407] & b[91])^(a[406] & b[92])^(a[405] & b[93])^(a[404] & b[94])^(a[403] & b[95])^(a[402] & b[96])^(a[401] & b[97])^(a[400] & b[98])^(a[399] & b[99])^(a[398] & b[100])^(a[397] & b[101])^(a[396] & b[102])^(a[395] & b[103])^(a[394] & b[104])^(a[393] & b[105])^(a[392] & b[106])^(a[391] & b[107])^(a[390] & b[108])^(a[389] & b[109])^(a[388] & b[110])^(a[387] & b[111])^(a[386] & b[112])^(a[385] & b[113])^(a[384] & b[114])^(a[383] & b[115])^(a[382] & b[116])^(a[381] & b[117])^(a[380] & b[118])^(a[379] & b[119])^(a[378] & b[120])^(a[377] & b[121])^(a[376] & b[122])^(a[375] & b[123])^(a[374] & b[124])^(a[373] & b[125])^(a[372] & b[126])^(a[371] & b[127])^(a[370] & b[128])^(a[369] & b[129])^(a[368] & b[130])^(a[367] & b[131])^(a[366] & b[132])^(a[365] & b[133])^(a[364] & b[134])^(a[363] & b[135])^(a[362] & b[136])^(a[361] & b[137])^(a[360] & b[138])^(a[359] & b[139])^(a[358] & b[140])^(a[357] & b[141])^(a[356] & b[142])^(a[355] & b[143])^(a[354] & b[144])^(a[353] & b[145])^(a[352] & b[146])^(a[351] & b[147])^(a[350] & b[148])^(a[349] & b[149])^(a[348] & b[150])^(a[347] & b[151])^(a[346] & b[152])^(a[345] & b[153])^(a[344] & b[154])^(a[343] & b[155])^(a[342] & b[156])^(a[341] & b[157])^(a[340] & b[158])^(a[339] & b[159])^(a[338] & b[160])^(a[337] & b[161])^(a[336] & b[162])^(a[335] & b[163])^(a[334] & b[164])^(a[333] & b[165])^(a[332] & b[166])^(a[331] & b[167])^(a[330] & b[168])^(a[329] & b[169])^(a[328] & b[170])^(a[327] & b[171])^(a[326] & b[172])^(a[325] & b[173])^(a[324] & b[174])^(a[323] & b[175])^(a[322] & b[176])^(a[321] & b[177])^(a[320] & b[178])^(a[319] & b[179])^(a[318] & b[180])^(a[317] & b[181])^(a[316] & b[182])^(a[315] & b[183])^(a[314] & b[184])^(a[313] & b[185])^(a[312] & b[186])^(a[311] & b[187])^(a[310] & b[188])^(a[309] & b[189])^(a[308] & b[190])^(a[307] & b[191])^(a[306] & b[192])^(a[305] & b[193])^(a[304] & b[194])^(a[303] & b[195])^(a[302] & b[196])^(a[301] & b[197])^(a[300] & b[198])^(a[299] & b[199])^(a[298] & b[200])^(a[297] & b[201])^(a[296] & b[202])^(a[295] & b[203])^(a[294] & b[204])^(a[293] & b[205])^(a[292] & b[206])^(a[291] & b[207])^(a[290] & b[208])^(a[289] & b[209])^(a[288] & b[210])^(a[287] & b[211])^(a[286] & b[212])^(a[285] & b[213])^(a[284] & b[214])^(a[283] & b[215])^(a[282] & b[216])^(a[281] & b[217])^(a[280] & b[218])^(a[279] & b[219])^(a[278] & b[220])^(a[277] & b[221])^(a[276] & b[222])^(a[275] & b[223])^(a[274] & b[224])^(a[273] & b[225])^(a[272] & b[226])^(a[271] & b[227])^(a[270] & b[228])^(a[269] & b[229])^(a[268] & b[230])^(a[267] & b[231])^(a[266] & b[232])^(a[265] & b[233])^(a[264] & b[234])^(a[263] & b[235])^(a[262] & b[236])^(a[261] & b[237])^(a[260] & b[238])^(a[259] & b[239])^(a[258] & b[240])^(a[257] & b[241])^(a[256] & b[242])^(a[255] & b[243])^(a[254] & b[244])^(a[253] & b[245])^(a[252] & b[246])^(a[251] & b[247])^(a[250] & b[248])^(a[249] & b[249])^(a[248] & b[250])^(a[247] & b[251])^(a[246] & b[252])^(a[245] & b[253])^(a[244] & b[254])^(a[243] & b[255])^(a[242] & b[256])^(a[241] & b[257])^(a[240] & b[258])^(a[239] & b[259])^(a[238] & b[260])^(a[237] & b[261])^(a[236] & b[262])^(a[235] & b[263])^(a[234] & b[264])^(a[233] & b[265])^(a[232] & b[266])^(a[231] & b[267])^(a[230] & b[268])^(a[229] & b[269])^(a[228] & b[270])^(a[227] & b[271])^(a[226] & b[272])^(a[225] & b[273])^(a[224] & b[274])^(a[223] & b[275])^(a[222] & b[276])^(a[221] & b[277])^(a[220] & b[278])^(a[219] & b[279])^(a[218] & b[280])^(a[217] & b[281])^(a[216] & b[282])^(a[215] & b[283])^(a[214] & b[284])^(a[213] & b[285])^(a[212] & b[286])^(a[211] & b[287])^(a[210] & b[288])^(a[209] & b[289])^(a[208] & b[290])^(a[207] & b[291])^(a[206] & b[292])^(a[205] & b[293])^(a[204] & b[294])^(a[203] & b[295])^(a[202] & b[296])^(a[201] & b[297])^(a[200] & b[298])^(a[199] & b[299])^(a[198] & b[300])^(a[197] & b[301])^(a[196] & b[302])^(a[195] & b[303])^(a[194] & b[304])^(a[193] & b[305])^(a[192] & b[306])^(a[191] & b[307])^(a[190] & b[308])^(a[189] & b[309])^(a[188] & b[310])^(a[187] & b[311])^(a[186] & b[312])^(a[185] & b[313])^(a[184] & b[314])^(a[183] & b[315])^(a[182] & b[316])^(a[181] & b[317])^(a[180] & b[318])^(a[179] & b[319])^(a[178] & b[320])^(a[177] & b[321])^(a[176] & b[322])^(a[175] & b[323])^(a[174] & b[324])^(a[173] & b[325])^(a[172] & b[326])^(a[171] & b[327])^(a[170] & b[328])^(a[169] & b[329])^(a[168] & b[330])^(a[167] & b[331])^(a[166] & b[332])^(a[165] & b[333])^(a[164] & b[334])^(a[163] & b[335])^(a[162] & b[336])^(a[161] & b[337])^(a[160] & b[338])^(a[159] & b[339])^(a[158] & b[340])^(a[157] & b[341])^(a[156] & b[342])^(a[155] & b[343])^(a[154] & b[344])^(a[153] & b[345])^(a[152] & b[346])^(a[151] & b[347])^(a[150] & b[348])^(a[149] & b[349])^(a[148] & b[350])^(a[147] & b[351])^(a[146] & b[352])^(a[145] & b[353])^(a[144] & b[354])^(a[143] & b[355])^(a[142] & b[356])^(a[141] & b[357])^(a[140] & b[358])^(a[139] & b[359])^(a[138] & b[360])^(a[137] & b[361])^(a[136] & b[362])^(a[135] & b[363])^(a[134] & b[364])^(a[133] & b[365])^(a[132] & b[366])^(a[131] & b[367])^(a[130] & b[368])^(a[129] & b[369])^(a[128] & b[370])^(a[127] & b[371])^(a[126] & b[372])^(a[125] & b[373])^(a[124] & b[374])^(a[123] & b[375])^(a[122] & b[376])^(a[121] & b[377])^(a[120] & b[378])^(a[119] & b[379])^(a[118] & b[380])^(a[117] & b[381])^(a[116] & b[382])^(a[115] & b[383])^(a[114] & b[384])^(a[113] & b[385])^(a[112] & b[386])^(a[111] & b[387])^(a[110] & b[388])^(a[109] & b[389])^(a[108] & b[390])^(a[107] & b[391])^(a[106] & b[392])^(a[105] & b[393])^(a[104] & b[394])^(a[103] & b[395])^(a[102] & b[396])^(a[101] & b[397])^(a[100] & b[398])^(a[99] & b[399])^(a[98] & b[400])^(a[97] & b[401])^(a[96] & b[402])^(a[95] & b[403])^(a[94] & b[404])^(a[93] & b[405])^(a[92] & b[406])^(a[91] & b[407])^(a[90] & b[408]);
assign y[499] = (a[408] & b[91])^(a[407] & b[92])^(a[406] & b[93])^(a[405] & b[94])^(a[404] & b[95])^(a[403] & b[96])^(a[402] & b[97])^(a[401] & b[98])^(a[400] & b[99])^(a[399] & b[100])^(a[398] & b[101])^(a[397] & b[102])^(a[396] & b[103])^(a[395] & b[104])^(a[394] & b[105])^(a[393] & b[106])^(a[392] & b[107])^(a[391] & b[108])^(a[390] & b[109])^(a[389] & b[110])^(a[388] & b[111])^(a[387] & b[112])^(a[386] & b[113])^(a[385] & b[114])^(a[384] & b[115])^(a[383] & b[116])^(a[382] & b[117])^(a[381] & b[118])^(a[380] & b[119])^(a[379] & b[120])^(a[378] & b[121])^(a[377] & b[122])^(a[376] & b[123])^(a[375] & b[124])^(a[374] & b[125])^(a[373] & b[126])^(a[372] & b[127])^(a[371] & b[128])^(a[370] & b[129])^(a[369] & b[130])^(a[368] & b[131])^(a[367] & b[132])^(a[366] & b[133])^(a[365] & b[134])^(a[364] & b[135])^(a[363] & b[136])^(a[362] & b[137])^(a[361] & b[138])^(a[360] & b[139])^(a[359] & b[140])^(a[358] & b[141])^(a[357] & b[142])^(a[356] & b[143])^(a[355] & b[144])^(a[354] & b[145])^(a[353] & b[146])^(a[352] & b[147])^(a[351] & b[148])^(a[350] & b[149])^(a[349] & b[150])^(a[348] & b[151])^(a[347] & b[152])^(a[346] & b[153])^(a[345] & b[154])^(a[344] & b[155])^(a[343] & b[156])^(a[342] & b[157])^(a[341] & b[158])^(a[340] & b[159])^(a[339] & b[160])^(a[338] & b[161])^(a[337] & b[162])^(a[336] & b[163])^(a[335] & b[164])^(a[334] & b[165])^(a[333] & b[166])^(a[332] & b[167])^(a[331] & b[168])^(a[330] & b[169])^(a[329] & b[170])^(a[328] & b[171])^(a[327] & b[172])^(a[326] & b[173])^(a[325] & b[174])^(a[324] & b[175])^(a[323] & b[176])^(a[322] & b[177])^(a[321] & b[178])^(a[320] & b[179])^(a[319] & b[180])^(a[318] & b[181])^(a[317] & b[182])^(a[316] & b[183])^(a[315] & b[184])^(a[314] & b[185])^(a[313] & b[186])^(a[312] & b[187])^(a[311] & b[188])^(a[310] & b[189])^(a[309] & b[190])^(a[308] & b[191])^(a[307] & b[192])^(a[306] & b[193])^(a[305] & b[194])^(a[304] & b[195])^(a[303] & b[196])^(a[302] & b[197])^(a[301] & b[198])^(a[300] & b[199])^(a[299] & b[200])^(a[298] & b[201])^(a[297] & b[202])^(a[296] & b[203])^(a[295] & b[204])^(a[294] & b[205])^(a[293] & b[206])^(a[292] & b[207])^(a[291] & b[208])^(a[290] & b[209])^(a[289] & b[210])^(a[288] & b[211])^(a[287] & b[212])^(a[286] & b[213])^(a[285] & b[214])^(a[284] & b[215])^(a[283] & b[216])^(a[282] & b[217])^(a[281] & b[218])^(a[280] & b[219])^(a[279] & b[220])^(a[278] & b[221])^(a[277] & b[222])^(a[276] & b[223])^(a[275] & b[224])^(a[274] & b[225])^(a[273] & b[226])^(a[272] & b[227])^(a[271] & b[228])^(a[270] & b[229])^(a[269] & b[230])^(a[268] & b[231])^(a[267] & b[232])^(a[266] & b[233])^(a[265] & b[234])^(a[264] & b[235])^(a[263] & b[236])^(a[262] & b[237])^(a[261] & b[238])^(a[260] & b[239])^(a[259] & b[240])^(a[258] & b[241])^(a[257] & b[242])^(a[256] & b[243])^(a[255] & b[244])^(a[254] & b[245])^(a[253] & b[246])^(a[252] & b[247])^(a[251] & b[248])^(a[250] & b[249])^(a[249] & b[250])^(a[248] & b[251])^(a[247] & b[252])^(a[246] & b[253])^(a[245] & b[254])^(a[244] & b[255])^(a[243] & b[256])^(a[242] & b[257])^(a[241] & b[258])^(a[240] & b[259])^(a[239] & b[260])^(a[238] & b[261])^(a[237] & b[262])^(a[236] & b[263])^(a[235] & b[264])^(a[234] & b[265])^(a[233] & b[266])^(a[232] & b[267])^(a[231] & b[268])^(a[230] & b[269])^(a[229] & b[270])^(a[228] & b[271])^(a[227] & b[272])^(a[226] & b[273])^(a[225] & b[274])^(a[224] & b[275])^(a[223] & b[276])^(a[222] & b[277])^(a[221] & b[278])^(a[220] & b[279])^(a[219] & b[280])^(a[218] & b[281])^(a[217] & b[282])^(a[216] & b[283])^(a[215] & b[284])^(a[214] & b[285])^(a[213] & b[286])^(a[212] & b[287])^(a[211] & b[288])^(a[210] & b[289])^(a[209] & b[290])^(a[208] & b[291])^(a[207] & b[292])^(a[206] & b[293])^(a[205] & b[294])^(a[204] & b[295])^(a[203] & b[296])^(a[202] & b[297])^(a[201] & b[298])^(a[200] & b[299])^(a[199] & b[300])^(a[198] & b[301])^(a[197] & b[302])^(a[196] & b[303])^(a[195] & b[304])^(a[194] & b[305])^(a[193] & b[306])^(a[192] & b[307])^(a[191] & b[308])^(a[190] & b[309])^(a[189] & b[310])^(a[188] & b[311])^(a[187] & b[312])^(a[186] & b[313])^(a[185] & b[314])^(a[184] & b[315])^(a[183] & b[316])^(a[182] & b[317])^(a[181] & b[318])^(a[180] & b[319])^(a[179] & b[320])^(a[178] & b[321])^(a[177] & b[322])^(a[176] & b[323])^(a[175] & b[324])^(a[174] & b[325])^(a[173] & b[326])^(a[172] & b[327])^(a[171] & b[328])^(a[170] & b[329])^(a[169] & b[330])^(a[168] & b[331])^(a[167] & b[332])^(a[166] & b[333])^(a[165] & b[334])^(a[164] & b[335])^(a[163] & b[336])^(a[162] & b[337])^(a[161] & b[338])^(a[160] & b[339])^(a[159] & b[340])^(a[158] & b[341])^(a[157] & b[342])^(a[156] & b[343])^(a[155] & b[344])^(a[154] & b[345])^(a[153] & b[346])^(a[152] & b[347])^(a[151] & b[348])^(a[150] & b[349])^(a[149] & b[350])^(a[148] & b[351])^(a[147] & b[352])^(a[146] & b[353])^(a[145] & b[354])^(a[144] & b[355])^(a[143] & b[356])^(a[142] & b[357])^(a[141] & b[358])^(a[140] & b[359])^(a[139] & b[360])^(a[138] & b[361])^(a[137] & b[362])^(a[136] & b[363])^(a[135] & b[364])^(a[134] & b[365])^(a[133] & b[366])^(a[132] & b[367])^(a[131] & b[368])^(a[130] & b[369])^(a[129] & b[370])^(a[128] & b[371])^(a[127] & b[372])^(a[126] & b[373])^(a[125] & b[374])^(a[124] & b[375])^(a[123] & b[376])^(a[122] & b[377])^(a[121] & b[378])^(a[120] & b[379])^(a[119] & b[380])^(a[118] & b[381])^(a[117] & b[382])^(a[116] & b[383])^(a[115] & b[384])^(a[114] & b[385])^(a[113] & b[386])^(a[112] & b[387])^(a[111] & b[388])^(a[110] & b[389])^(a[109] & b[390])^(a[108] & b[391])^(a[107] & b[392])^(a[106] & b[393])^(a[105] & b[394])^(a[104] & b[395])^(a[103] & b[396])^(a[102] & b[397])^(a[101] & b[398])^(a[100] & b[399])^(a[99] & b[400])^(a[98] & b[401])^(a[97] & b[402])^(a[96] & b[403])^(a[95] & b[404])^(a[94] & b[405])^(a[93] & b[406])^(a[92] & b[407])^(a[91] & b[408]);
assign y[500] = (a[408] & b[92])^(a[407] & b[93])^(a[406] & b[94])^(a[405] & b[95])^(a[404] & b[96])^(a[403] & b[97])^(a[402] & b[98])^(a[401] & b[99])^(a[400] & b[100])^(a[399] & b[101])^(a[398] & b[102])^(a[397] & b[103])^(a[396] & b[104])^(a[395] & b[105])^(a[394] & b[106])^(a[393] & b[107])^(a[392] & b[108])^(a[391] & b[109])^(a[390] & b[110])^(a[389] & b[111])^(a[388] & b[112])^(a[387] & b[113])^(a[386] & b[114])^(a[385] & b[115])^(a[384] & b[116])^(a[383] & b[117])^(a[382] & b[118])^(a[381] & b[119])^(a[380] & b[120])^(a[379] & b[121])^(a[378] & b[122])^(a[377] & b[123])^(a[376] & b[124])^(a[375] & b[125])^(a[374] & b[126])^(a[373] & b[127])^(a[372] & b[128])^(a[371] & b[129])^(a[370] & b[130])^(a[369] & b[131])^(a[368] & b[132])^(a[367] & b[133])^(a[366] & b[134])^(a[365] & b[135])^(a[364] & b[136])^(a[363] & b[137])^(a[362] & b[138])^(a[361] & b[139])^(a[360] & b[140])^(a[359] & b[141])^(a[358] & b[142])^(a[357] & b[143])^(a[356] & b[144])^(a[355] & b[145])^(a[354] & b[146])^(a[353] & b[147])^(a[352] & b[148])^(a[351] & b[149])^(a[350] & b[150])^(a[349] & b[151])^(a[348] & b[152])^(a[347] & b[153])^(a[346] & b[154])^(a[345] & b[155])^(a[344] & b[156])^(a[343] & b[157])^(a[342] & b[158])^(a[341] & b[159])^(a[340] & b[160])^(a[339] & b[161])^(a[338] & b[162])^(a[337] & b[163])^(a[336] & b[164])^(a[335] & b[165])^(a[334] & b[166])^(a[333] & b[167])^(a[332] & b[168])^(a[331] & b[169])^(a[330] & b[170])^(a[329] & b[171])^(a[328] & b[172])^(a[327] & b[173])^(a[326] & b[174])^(a[325] & b[175])^(a[324] & b[176])^(a[323] & b[177])^(a[322] & b[178])^(a[321] & b[179])^(a[320] & b[180])^(a[319] & b[181])^(a[318] & b[182])^(a[317] & b[183])^(a[316] & b[184])^(a[315] & b[185])^(a[314] & b[186])^(a[313] & b[187])^(a[312] & b[188])^(a[311] & b[189])^(a[310] & b[190])^(a[309] & b[191])^(a[308] & b[192])^(a[307] & b[193])^(a[306] & b[194])^(a[305] & b[195])^(a[304] & b[196])^(a[303] & b[197])^(a[302] & b[198])^(a[301] & b[199])^(a[300] & b[200])^(a[299] & b[201])^(a[298] & b[202])^(a[297] & b[203])^(a[296] & b[204])^(a[295] & b[205])^(a[294] & b[206])^(a[293] & b[207])^(a[292] & b[208])^(a[291] & b[209])^(a[290] & b[210])^(a[289] & b[211])^(a[288] & b[212])^(a[287] & b[213])^(a[286] & b[214])^(a[285] & b[215])^(a[284] & b[216])^(a[283] & b[217])^(a[282] & b[218])^(a[281] & b[219])^(a[280] & b[220])^(a[279] & b[221])^(a[278] & b[222])^(a[277] & b[223])^(a[276] & b[224])^(a[275] & b[225])^(a[274] & b[226])^(a[273] & b[227])^(a[272] & b[228])^(a[271] & b[229])^(a[270] & b[230])^(a[269] & b[231])^(a[268] & b[232])^(a[267] & b[233])^(a[266] & b[234])^(a[265] & b[235])^(a[264] & b[236])^(a[263] & b[237])^(a[262] & b[238])^(a[261] & b[239])^(a[260] & b[240])^(a[259] & b[241])^(a[258] & b[242])^(a[257] & b[243])^(a[256] & b[244])^(a[255] & b[245])^(a[254] & b[246])^(a[253] & b[247])^(a[252] & b[248])^(a[251] & b[249])^(a[250] & b[250])^(a[249] & b[251])^(a[248] & b[252])^(a[247] & b[253])^(a[246] & b[254])^(a[245] & b[255])^(a[244] & b[256])^(a[243] & b[257])^(a[242] & b[258])^(a[241] & b[259])^(a[240] & b[260])^(a[239] & b[261])^(a[238] & b[262])^(a[237] & b[263])^(a[236] & b[264])^(a[235] & b[265])^(a[234] & b[266])^(a[233] & b[267])^(a[232] & b[268])^(a[231] & b[269])^(a[230] & b[270])^(a[229] & b[271])^(a[228] & b[272])^(a[227] & b[273])^(a[226] & b[274])^(a[225] & b[275])^(a[224] & b[276])^(a[223] & b[277])^(a[222] & b[278])^(a[221] & b[279])^(a[220] & b[280])^(a[219] & b[281])^(a[218] & b[282])^(a[217] & b[283])^(a[216] & b[284])^(a[215] & b[285])^(a[214] & b[286])^(a[213] & b[287])^(a[212] & b[288])^(a[211] & b[289])^(a[210] & b[290])^(a[209] & b[291])^(a[208] & b[292])^(a[207] & b[293])^(a[206] & b[294])^(a[205] & b[295])^(a[204] & b[296])^(a[203] & b[297])^(a[202] & b[298])^(a[201] & b[299])^(a[200] & b[300])^(a[199] & b[301])^(a[198] & b[302])^(a[197] & b[303])^(a[196] & b[304])^(a[195] & b[305])^(a[194] & b[306])^(a[193] & b[307])^(a[192] & b[308])^(a[191] & b[309])^(a[190] & b[310])^(a[189] & b[311])^(a[188] & b[312])^(a[187] & b[313])^(a[186] & b[314])^(a[185] & b[315])^(a[184] & b[316])^(a[183] & b[317])^(a[182] & b[318])^(a[181] & b[319])^(a[180] & b[320])^(a[179] & b[321])^(a[178] & b[322])^(a[177] & b[323])^(a[176] & b[324])^(a[175] & b[325])^(a[174] & b[326])^(a[173] & b[327])^(a[172] & b[328])^(a[171] & b[329])^(a[170] & b[330])^(a[169] & b[331])^(a[168] & b[332])^(a[167] & b[333])^(a[166] & b[334])^(a[165] & b[335])^(a[164] & b[336])^(a[163] & b[337])^(a[162] & b[338])^(a[161] & b[339])^(a[160] & b[340])^(a[159] & b[341])^(a[158] & b[342])^(a[157] & b[343])^(a[156] & b[344])^(a[155] & b[345])^(a[154] & b[346])^(a[153] & b[347])^(a[152] & b[348])^(a[151] & b[349])^(a[150] & b[350])^(a[149] & b[351])^(a[148] & b[352])^(a[147] & b[353])^(a[146] & b[354])^(a[145] & b[355])^(a[144] & b[356])^(a[143] & b[357])^(a[142] & b[358])^(a[141] & b[359])^(a[140] & b[360])^(a[139] & b[361])^(a[138] & b[362])^(a[137] & b[363])^(a[136] & b[364])^(a[135] & b[365])^(a[134] & b[366])^(a[133] & b[367])^(a[132] & b[368])^(a[131] & b[369])^(a[130] & b[370])^(a[129] & b[371])^(a[128] & b[372])^(a[127] & b[373])^(a[126] & b[374])^(a[125] & b[375])^(a[124] & b[376])^(a[123] & b[377])^(a[122] & b[378])^(a[121] & b[379])^(a[120] & b[380])^(a[119] & b[381])^(a[118] & b[382])^(a[117] & b[383])^(a[116] & b[384])^(a[115] & b[385])^(a[114] & b[386])^(a[113] & b[387])^(a[112] & b[388])^(a[111] & b[389])^(a[110] & b[390])^(a[109] & b[391])^(a[108] & b[392])^(a[107] & b[393])^(a[106] & b[394])^(a[105] & b[395])^(a[104] & b[396])^(a[103] & b[397])^(a[102] & b[398])^(a[101] & b[399])^(a[100] & b[400])^(a[99] & b[401])^(a[98] & b[402])^(a[97] & b[403])^(a[96] & b[404])^(a[95] & b[405])^(a[94] & b[406])^(a[93] & b[407])^(a[92] & b[408]);
assign y[501] = (a[408] & b[93])^(a[407] & b[94])^(a[406] & b[95])^(a[405] & b[96])^(a[404] & b[97])^(a[403] & b[98])^(a[402] & b[99])^(a[401] & b[100])^(a[400] & b[101])^(a[399] & b[102])^(a[398] & b[103])^(a[397] & b[104])^(a[396] & b[105])^(a[395] & b[106])^(a[394] & b[107])^(a[393] & b[108])^(a[392] & b[109])^(a[391] & b[110])^(a[390] & b[111])^(a[389] & b[112])^(a[388] & b[113])^(a[387] & b[114])^(a[386] & b[115])^(a[385] & b[116])^(a[384] & b[117])^(a[383] & b[118])^(a[382] & b[119])^(a[381] & b[120])^(a[380] & b[121])^(a[379] & b[122])^(a[378] & b[123])^(a[377] & b[124])^(a[376] & b[125])^(a[375] & b[126])^(a[374] & b[127])^(a[373] & b[128])^(a[372] & b[129])^(a[371] & b[130])^(a[370] & b[131])^(a[369] & b[132])^(a[368] & b[133])^(a[367] & b[134])^(a[366] & b[135])^(a[365] & b[136])^(a[364] & b[137])^(a[363] & b[138])^(a[362] & b[139])^(a[361] & b[140])^(a[360] & b[141])^(a[359] & b[142])^(a[358] & b[143])^(a[357] & b[144])^(a[356] & b[145])^(a[355] & b[146])^(a[354] & b[147])^(a[353] & b[148])^(a[352] & b[149])^(a[351] & b[150])^(a[350] & b[151])^(a[349] & b[152])^(a[348] & b[153])^(a[347] & b[154])^(a[346] & b[155])^(a[345] & b[156])^(a[344] & b[157])^(a[343] & b[158])^(a[342] & b[159])^(a[341] & b[160])^(a[340] & b[161])^(a[339] & b[162])^(a[338] & b[163])^(a[337] & b[164])^(a[336] & b[165])^(a[335] & b[166])^(a[334] & b[167])^(a[333] & b[168])^(a[332] & b[169])^(a[331] & b[170])^(a[330] & b[171])^(a[329] & b[172])^(a[328] & b[173])^(a[327] & b[174])^(a[326] & b[175])^(a[325] & b[176])^(a[324] & b[177])^(a[323] & b[178])^(a[322] & b[179])^(a[321] & b[180])^(a[320] & b[181])^(a[319] & b[182])^(a[318] & b[183])^(a[317] & b[184])^(a[316] & b[185])^(a[315] & b[186])^(a[314] & b[187])^(a[313] & b[188])^(a[312] & b[189])^(a[311] & b[190])^(a[310] & b[191])^(a[309] & b[192])^(a[308] & b[193])^(a[307] & b[194])^(a[306] & b[195])^(a[305] & b[196])^(a[304] & b[197])^(a[303] & b[198])^(a[302] & b[199])^(a[301] & b[200])^(a[300] & b[201])^(a[299] & b[202])^(a[298] & b[203])^(a[297] & b[204])^(a[296] & b[205])^(a[295] & b[206])^(a[294] & b[207])^(a[293] & b[208])^(a[292] & b[209])^(a[291] & b[210])^(a[290] & b[211])^(a[289] & b[212])^(a[288] & b[213])^(a[287] & b[214])^(a[286] & b[215])^(a[285] & b[216])^(a[284] & b[217])^(a[283] & b[218])^(a[282] & b[219])^(a[281] & b[220])^(a[280] & b[221])^(a[279] & b[222])^(a[278] & b[223])^(a[277] & b[224])^(a[276] & b[225])^(a[275] & b[226])^(a[274] & b[227])^(a[273] & b[228])^(a[272] & b[229])^(a[271] & b[230])^(a[270] & b[231])^(a[269] & b[232])^(a[268] & b[233])^(a[267] & b[234])^(a[266] & b[235])^(a[265] & b[236])^(a[264] & b[237])^(a[263] & b[238])^(a[262] & b[239])^(a[261] & b[240])^(a[260] & b[241])^(a[259] & b[242])^(a[258] & b[243])^(a[257] & b[244])^(a[256] & b[245])^(a[255] & b[246])^(a[254] & b[247])^(a[253] & b[248])^(a[252] & b[249])^(a[251] & b[250])^(a[250] & b[251])^(a[249] & b[252])^(a[248] & b[253])^(a[247] & b[254])^(a[246] & b[255])^(a[245] & b[256])^(a[244] & b[257])^(a[243] & b[258])^(a[242] & b[259])^(a[241] & b[260])^(a[240] & b[261])^(a[239] & b[262])^(a[238] & b[263])^(a[237] & b[264])^(a[236] & b[265])^(a[235] & b[266])^(a[234] & b[267])^(a[233] & b[268])^(a[232] & b[269])^(a[231] & b[270])^(a[230] & b[271])^(a[229] & b[272])^(a[228] & b[273])^(a[227] & b[274])^(a[226] & b[275])^(a[225] & b[276])^(a[224] & b[277])^(a[223] & b[278])^(a[222] & b[279])^(a[221] & b[280])^(a[220] & b[281])^(a[219] & b[282])^(a[218] & b[283])^(a[217] & b[284])^(a[216] & b[285])^(a[215] & b[286])^(a[214] & b[287])^(a[213] & b[288])^(a[212] & b[289])^(a[211] & b[290])^(a[210] & b[291])^(a[209] & b[292])^(a[208] & b[293])^(a[207] & b[294])^(a[206] & b[295])^(a[205] & b[296])^(a[204] & b[297])^(a[203] & b[298])^(a[202] & b[299])^(a[201] & b[300])^(a[200] & b[301])^(a[199] & b[302])^(a[198] & b[303])^(a[197] & b[304])^(a[196] & b[305])^(a[195] & b[306])^(a[194] & b[307])^(a[193] & b[308])^(a[192] & b[309])^(a[191] & b[310])^(a[190] & b[311])^(a[189] & b[312])^(a[188] & b[313])^(a[187] & b[314])^(a[186] & b[315])^(a[185] & b[316])^(a[184] & b[317])^(a[183] & b[318])^(a[182] & b[319])^(a[181] & b[320])^(a[180] & b[321])^(a[179] & b[322])^(a[178] & b[323])^(a[177] & b[324])^(a[176] & b[325])^(a[175] & b[326])^(a[174] & b[327])^(a[173] & b[328])^(a[172] & b[329])^(a[171] & b[330])^(a[170] & b[331])^(a[169] & b[332])^(a[168] & b[333])^(a[167] & b[334])^(a[166] & b[335])^(a[165] & b[336])^(a[164] & b[337])^(a[163] & b[338])^(a[162] & b[339])^(a[161] & b[340])^(a[160] & b[341])^(a[159] & b[342])^(a[158] & b[343])^(a[157] & b[344])^(a[156] & b[345])^(a[155] & b[346])^(a[154] & b[347])^(a[153] & b[348])^(a[152] & b[349])^(a[151] & b[350])^(a[150] & b[351])^(a[149] & b[352])^(a[148] & b[353])^(a[147] & b[354])^(a[146] & b[355])^(a[145] & b[356])^(a[144] & b[357])^(a[143] & b[358])^(a[142] & b[359])^(a[141] & b[360])^(a[140] & b[361])^(a[139] & b[362])^(a[138] & b[363])^(a[137] & b[364])^(a[136] & b[365])^(a[135] & b[366])^(a[134] & b[367])^(a[133] & b[368])^(a[132] & b[369])^(a[131] & b[370])^(a[130] & b[371])^(a[129] & b[372])^(a[128] & b[373])^(a[127] & b[374])^(a[126] & b[375])^(a[125] & b[376])^(a[124] & b[377])^(a[123] & b[378])^(a[122] & b[379])^(a[121] & b[380])^(a[120] & b[381])^(a[119] & b[382])^(a[118] & b[383])^(a[117] & b[384])^(a[116] & b[385])^(a[115] & b[386])^(a[114] & b[387])^(a[113] & b[388])^(a[112] & b[389])^(a[111] & b[390])^(a[110] & b[391])^(a[109] & b[392])^(a[108] & b[393])^(a[107] & b[394])^(a[106] & b[395])^(a[105] & b[396])^(a[104] & b[397])^(a[103] & b[398])^(a[102] & b[399])^(a[101] & b[400])^(a[100] & b[401])^(a[99] & b[402])^(a[98] & b[403])^(a[97] & b[404])^(a[96] & b[405])^(a[95] & b[406])^(a[94] & b[407])^(a[93] & b[408]);
assign y[502] = (a[408] & b[94])^(a[407] & b[95])^(a[406] & b[96])^(a[405] & b[97])^(a[404] & b[98])^(a[403] & b[99])^(a[402] & b[100])^(a[401] & b[101])^(a[400] & b[102])^(a[399] & b[103])^(a[398] & b[104])^(a[397] & b[105])^(a[396] & b[106])^(a[395] & b[107])^(a[394] & b[108])^(a[393] & b[109])^(a[392] & b[110])^(a[391] & b[111])^(a[390] & b[112])^(a[389] & b[113])^(a[388] & b[114])^(a[387] & b[115])^(a[386] & b[116])^(a[385] & b[117])^(a[384] & b[118])^(a[383] & b[119])^(a[382] & b[120])^(a[381] & b[121])^(a[380] & b[122])^(a[379] & b[123])^(a[378] & b[124])^(a[377] & b[125])^(a[376] & b[126])^(a[375] & b[127])^(a[374] & b[128])^(a[373] & b[129])^(a[372] & b[130])^(a[371] & b[131])^(a[370] & b[132])^(a[369] & b[133])^(a[368] & b[134])^(a[367] & b[135])^(a[366] & b[136])^(a[365] & b[137])^(a[364] & b[138])^(a[363] & b[139])^(a[362] & b[140])^(a[361] & b[141])^(a[360] & b[142])^(a[359] & b[143])^(a[358] & b[144])^(a[357] & b[145])^(a[356] & b[146])^(a[355] & b[147])^(a[354] & b[148])^(a[353] & b[149])^(a[352] & b[150])^(a[351] & b[151])^(a[350] & b[152])^(a[349] & b[153])^(a[348] & b[154])^(a[347] & b[155])^(a[346] & b[156])^(a[345] & b[157])^(a[344] & b[158])^(a[343] & b[159])^(a[342] & b[160])^(a[341] & b[161])^(a[340] & b[162])^(a[339] & b[163])^(a[338] & b[164])^(a[337] & b[165])^(a[336] & b[166])^(a[335] & b[167])^(a[334] & b[168])^(a[333] & b[169])^(a[332] & b[170])^(a[331] & b[171])^(a[330] & b[172])^(a[329] & b[173])^(a[328] & b[174])^(a[327] & b[175])^(a[326] & b[176])^(a[325] & b[177])^(a[324] & b[178])^(a[323] & b[179])^(a[322] & b[180])^(a[321] & b[181])^(a[320] & b[182])^(a[319] & b[183])^(a[318] & b[184])^(a[317] & b[185])^(a[316] & b[186])^(a[315] & b[187])^(a[314] & b[188])^(a[313] & b[189])^(a[312] & b[190])^(a[311] & b[191])^(a[310] & b[192])^(a[309] & b[193])^(a[308] & b[194])^(a[307] & b[195])^(a[306] & b[196])^(a[305] & b[197])^(a[304] & b[198])^(a[303] & b[199])^(a[302] & b[200])^(a[301] & b[201])^(a[300] & b[202])^(a[299] & b[203])^(a[298] & b[204])^(a[297] & b[205])^(a[296] & b[206])^(a[295] & b[207])^(a[294] & b[208])^(a[293] & b[209])^(a[292] & b[210])^(a[291] & b[211])^(a[290] & b[212])^(a[289] & b[213])^(a[288] & b[214])^(a[287] & b[215])^(a[286] & b[216])^(a[285] & b[217])^(a[284] & b[218])^(a[283] & b[219])^(a[282] & b[220])^(a[281] & b[221])^(a[280] & b[222])^(a[279] & b[223])^(a[278] & b[224])^(a[277] & b[225])^(a[276] & b[226])^(a[275] & b[227])^(a[274] & b[228])^(a[273] & b[229])^(a[272] & b[230])^(a[271] & b[231])^(a[270] & b[232])^(a[269] & b[233])^(a[268] & b[234])^(a[267] & b[235])^(a[266] & b[236])^(a[265] & b[237])^(a[264] & b[238])^(a[263] & b[239])^(a[262] & b[240])^(a[261] & b[241])^(a[260] & b[242])^(a[259] & b[243])^(a[258] & b[244])^(a[257] & b[245])^(a[256] & b[246])^(a[255] & b[247])^(a[254] & b[248])^(a[253] & b[249])^(a[252] & b[250])^(a[251] & b[251])^(a[250] & b[252])^(a[249] & b[253])^(a[248] & b[254])^(a[247] & b[255])^(a[246] & b[256])^(a[245] & b[257])^(a[244] & b[258])^(a[243] & b[259])^(a[242] & b[260])^(a[241] & b[261])^(a[240] & b[262])^(a[239] & b[263])^(a[238] & b[264])^(a[237] & b[265])^(a[236] & b[266])^(a[235] & b[267])^(a[234] & b[268])^(a[233] & b[269])^(a[232] & b[270])^(a[231] & b[271])^(a[230] & b[272])^(a[229] & b[273])^(a[228] & b[274])^(a[227] & b[275])^(a[226] & b[276])^(a[225] & b[277])^(a[224] & b[278])^(a[223] & b[279])^(a[222] & b[280])^(a[221] & b[281])^(a[220] & b[282])^(a[219] & b[283])^(a[218] & b[284])^(a[217] & b[285])^(a[216] & b[286])^(a[215] & b[287])^(a[214] & b[288])^(a[213] & b[289])^(a[212] & b[290])^(a[211] & b[291])^(a[210] & b[292])^(a[209] & b[293])^(a[208] & b[294])^(a[207] & b[295])^(a[206] & b[296])^(a[205] & b[297])^(a[204] & b[298])^(a[203] & b[299])^(a[202] & b[300])^(a[201] & b[301])^(a[200] & b[302])^(a[199] & b[303])^(a[198] & b[304])^(a[197] & b[305])^(a[196] & b[306])^(a[195] & b[307])^(a[194] & b[308])^(a[193] & b[309])^(a[192] & b[310])^(a[191] & b[311])^(a[190] & b[312])^(a[189] & b[313])^(a[188] & b[314])^(a[187] & b[315])^(a[186] & b[316])^(a[185] & b[317])^(a[184] & b[318])^(a[183] & b[319])^(a[182] & b[320])^(a[181] & b[321])^(a[180] & b[322])^(a[179] & b[323])^(a[178] & b[324])^(a[177] & b[325])^(a[176] & b[326])^(a[175] & b[327])^(a[174] & b[328])^(a[173] & b[329])^(a[172] & b[330])^(a[171] & b[331])^(a[170] & b[332])^(a[169] & b[333])^(a[168] & b[334])^(a[167] & b[335])^(a[166] & b[336])^(a[165] & b[337])^(a[164] & b[338])^(a[163] & b[339])^(a[162] & b[340])^(a[161] & b[341])^(a[160] & b[342])^(a[159] & b[343])^(a[158] & b[344])^(a[157] & b[345])^(a[156] & b[346])^(a[155] & b[347])^(a[154] & b[348])^(a[153] & b[349])^(a[152] & b[350])^(a[151] & b[351])^(a[150] & b[352])^(a[149] & b[353])^(a[148] & b[354])^(a[147] & b[355])^(a[146] & b[356])^(a[145] & b[357])^(a[144] & b[358])^(a[143] & b[359])^(a[142] & b[360])^(a[141] & b[361])^(a[140] & b[362])^(a[139] & b[363])^(a[138] & b[364])^(a[137] & b[365])^(a[136] & b[366])^(a[135] & b[367])^(a[134] & b[368])^(a[133] & b[369])^(a[132] & b[370])^(a[131] & b[371])^(a[130] & b[372])^(a[129] & b[373])^(a[128] & b[374])^(a[127] & b[375])^(a[126] & b[376])^(a[125] & b[377])^(a[124] & b[378])^(a[123] & b[379])^(a[122] & b[380])^(a[121] & b[381])^(a[120] & b[382])^(a[119] & b[383])^(a[118] & b[384])^(a[117] & b[385])^(a[116] & b[386])^(a[115] & b[387])^(a[114] & b[388])^(a[113] & b[389])^(a[112] & b[390])^(a[111] & b[391])^(a[110] & b[392])^(a[109] & b[393])^(a[108] & b[394])^(a[107] & b[395])^(a[106] & b[396])^(a[105] & b[397])^(a[104] & b[398])^(a[103] & b[399])^(a[102] & b[400])^(a[101] & b[401])^(a[100] & b[402])^(a[99] & b[403])^(a[98] & b[404])^(a[97] & b[405])^(a[96] & b[406])^(a[95] & b[407])^(a[94] & b[408]);
assign y[503] = (a[408] & b[95])^(a[407] & b[96])^(a[406] & b[97])^(a[405] & b[98])^(a[404] & b[99])^(a[403] & b[100])^(a[402] & b[101])^(a[401] & b[102])^(a[400] & b[103])^(a[399] & b[104])^(a[398] & b[105])^(a[397] & b[106])^(a[396] & b[107])^(a[395] & b[108])^(a[394] & b[109])^(a[393] & b[110])^(a[392] & b[111])^(a[391] & b[112])^(a[390] & b[113])^(a[389] & b[114])^(a[388] & b[115])^(a[387] & b[116])^(a[386] & b[117])^(a[385] & b[118])^(a[384] & b[119])^(a[383] & b[120])^(a[382] & b[121])^(a[381] & b[122])^(a[380] & b[123])^(a[379] & b[124])^(a[378] & b[125])^(a[377] & b[126])^(a[376] & b[127])^(a[375] & b[128])^(a[374] & b[129])^(a[373] & b[130])^(a[372] & b[131])^(a[371] & b[132])^(a[370] & b[133])^(a[369] & b[134])^(a[368] & b[135])^(a[367] & b[136])^(a[366] & b[137])^(a[365] & b[138])^(a[364] & b[139])^(a[363] & b[140])^(a[362] & b[141])^(a[361] & b[142])^(a[360] & b[143])^(a[359] & b[144])^(a[358] & b[145])^(a[357] & b[146])^(a[356] & b[147])^(a[355] & b[148])^(a[354] & b[149])^(a[353] & b[150])^(a[352] & b[151])^(a[351] & b[152])^(a[350] & b[153])^(a[349] & b[154])^(a[348] & b[155])^(a[347] & b[156])^(a[346] & b[157])^(a[345] & b[158])^(a[344] & b[159])^(a[343] & b[160])^(a[342] & b[161])^(a[341] & b[162])^(a[340] & b[163])^(a[339] & b[164])^(a[338] & b[165])^(a[337] & b[166])^(a[336] & b[167])^(a[335] & b[168])^(a[334] & b[169])^(a[333] & b[170])^(a[332] & b[171])^(a[331] & b[172])^(a[330] & b[173])^(a[329] & b[174])^(a[328] & b[175])^(a[327] & b[176])^(a[326] & b[177])^(a[325] & b[178])^(a[324] & b[179])^(a[323] & b[180])^(a[322] & b[181])^(a[321] & b[182])^(a[320] & b[183])^(a[319] & b[184])^(a[318] & b[185])^(a[317] & b[186])^(a[316] & b[187])^(a[315] & b[188])^(a[314] & b[189])^(a[313] & b[190])^(a[312] & b[191])^(a[311] & b[192])^(a[310] & b[193])^(a[309] & b[194])^(a[308] & b[195])^(a[307] & b[196])^(a[306] & b[197])^(a[305] & b[198])^(a[304] & b[199])^(a[303] & b[200])^(a[302] & b[201])^(a[301] & b[202])^(a[300] & b[203])^(a[299] & b[204])^(a[298] & b[205])^(a[297] & b[206])^(a[296] & b[207])^(a[295] & b[208])^(a[294] & b[209])^(a[293] & b[210])^(a[292] & b[211])^(a[291] & b[212])^(a[290] & b[213])^(a[289] & b[214])^(a[288] & b[215])^(a[287] & b[216])^(a[286] & b[217])^(a[285] & b[218])^(a[284] & b[219])^(a[283] & b[220])^(a[282] & b[221])^(a[281] & b[222])^(a[280] & b[223])^(a[279] & b[224])^(a[278] & b[225])^(a[277] & b[226])^(a[276] & b[227])^(a[275] & b[228])^(a[274] & b[229])^(a[273] & b[230])^(a[272] & b[231])^(a[271] & b[232])^(a[270] & b[233])^(a[269] & b[234])^(a[268] & b[235])^(a[267] & b[236])^(a[266] & b[237])^(a[265] & b[238])^(a[264] & b[239])^(a[263] & b[240])^(a[262] & b[241])^(a[261] & b[242])^(a[260] & b[243])^(a[259] & b[244])^(a[258] & b[245])^(a[257] & b[246])^(a[256] & b[247])^(a[255] & b[248])^(a[254] & b[249])^(a[253] & b[250])^(a[252] & b[251])^(a[251] & b[252])^(a[250] & b[253])^(a[249] & b[254])^(a[248] & b[255])^(a[247] & b[256])^(a[246] & b[257])^(a[245] & b[258])^(a[244] & b[259])^(a[243] & b[260])^(a[242] & b[261])^(a[241] & b[262])^(a[240] & b[263])^(a[239] & b[264])^(a[238] & b[265])^(a[237] & b[266])^(a[236] & b[267])^(a[235] & b[268])^(a[234] & b[269])^(a[233] & b[270])^(a[232] & b[271])^(a[231] & b[272])^(a[230] & b[273])^(a[229] & b[274])^(a[228] & b[275])^(a[227] & b[276])^(a[226] & b[277])^(a[225] & b[278])^(a[224] & b[279])^(a[223] & b[280])^(a[222] & b[281])^(a[221] & b[282])^(a[220] & b[283])^(a[219] & b[284])^(a[218] & b[285])^(a[217] & b[286])^(a[216] & b[287])^(a[215] & b[288])^(a[214] & b[289])^(a[213] & b[290])^(a[212] & b[291])^(a[211] & b[292])^(a[210] & b[293])^(a[209] & b[294])^(a[208] & b[295])^(a[207] & b[296])^(a[206] & b[297])^(a[205] & b[298])^(a[204] & b[299])^(a[203] & b[300])^(a[202] & b[301])^(a[201] & b[302])^(a[200] & b[303])^(a[199] & b[304])^(a[198] & b[305])^(a[197] & b[306])^(a[196] & b[307])^(a[195] & b[308])^(a[194] & b[309])^(a[193] & b[310])^(a[192] & b[311])^(a[191] & b[312])^(a[190] & b[313])^(a[189] & b[314])^(a[188] & b[315])^(a[187] & b[316])^(a[186] & b[317])^(a[185] & b[318])^(a[184] & b[319])^(a[183] & b[320])^(a[182] & b[321])^(a[181] & b[322])^(a[180] & b[323])^(a[179] & b[324])^(a[178] & b[325])^(a[177] & b[326])^(a[176] & b[327])^(a[175] & b[328])^(a[174] & b[329])^(a[173] & b[330])^(a[172] & b[331])^(a[171] & b[332])^(a[170] & b[333])^(a[169] & b[334])^(a[168] & b[335])^(a[167] & b[336])^(a[166] & b[337])^(a[165] & b[338])^(a[164] & b[339])^(a[163] & b[340])^(a[162] & b[341])^(a[161] & b[342])^(a[160] & b[343])^(a[159] & b[344])^(a[158] & b[345])^(a[157] & b[346])^(a[156] & b[347])^(a[155] & b[348])^(a[154] & b[349])^(a[153] & b[350])^(a[152] & b[351])^(a[151] & b[352])^(a[150] & b[353])^(a[149] & b[354])^(a[148] & b[355])^(a[147] & b[356])^(a[146] & b[357])^(a[145] & b[358])^(a[144] & b[359])^(a[143] & b[360])^(a[142] & b[361])^(a[141] & b[362])^(a[140] & b[363])^(a[139] & b[364])^(a[138] & b[365])^(a[137] & b[366])^(a[136] & b[367])^(a[135] & b[368])^(a[134] & b[369])^(a[133] & b[370])^(a[132] & b[371])^(a[131] & b[372])^(a[130] & b[373])^(a[129] & b[374])^(a[128] & b[375])^(a[127] & b[376])^(a[126] & b[377])^(a[125] & b[378])^(a[124] & b[379])^(a[123] & b[380])^(a[122] & b[381])^(a[121] & b[382])^(a[120] & b[383])^(a[119] & b[384])^(a[118] & b[385])^(a[117] & b[386])^(a[116] & b[387])^(a[115] & b[388])^(a[114] & b[389])^(a[113] & b[390])^(a[112] & b[391])^(a[111] & b[392])^(a[110] & b[393])^(a[109] & b[394])^(a[108] & b[395])^(a[107] & b[396])^(a[106] & b[397])^(a[105] & b[398])^(a[104] & b[399])^(a[103] & b[400])^(a[102] & b[401])^(a[101] & b[402])^(a[100] & b[403])^(a[99] & b[404])^(a[98] & b[405])^(a[97] & b[406])^(a[96] & b[407])^(a[95] & b[408]);
assign y[504] = (a[408] & b[96])^(a[407] & b[97])^(a[406] & b[98])^(a[405] & b[99])^(a[404] & b[100])^(a[403] & b[101])^(a[402] & b[102])^(a[401] & b[103])^(a[400] & b[104])^(a[399] & b[105])^(a[398] & b[106])^(a[397] & b[107])^(a[396] & b[108])^(a[395] & b[109])^(a[394] & b[110])^(a[393] & b[111])^(a[392] & b[112])^(a[391] & b[113])^(a[390] & b[114])^(a[389] & b[115])^(a[388] & b[116])^(a[387] & b[117])^(a[386] & b[118])^(a[385] & b[119])^(a[384] & b[120])^(a[383] & b[121])^(a[382] & b[122])^(a[381] & b[123])^(a[380] & b[124])^(a[379] & b[125])^(a[378] & b[126])^(a[377] & b[127])^(a[376] & b[128])^(a[375] & b[129])^(a[374] & b[130])^(a[373] & b[131])^(a[372] & b[132])^(a[371] & b[133])^(a[370] & b[134])^(a[369] & b[135])^(a[368] & b[136])^(a[367] & b[137])^(a[366] & b[138])^(a[365] & b[139])^(a[364] & b[140])^(a[363] & b[141])^(a[362] & b[142])^(a[361] & b[143])^(a[360] & b[144])^(a[359] & b[145])^(a[358] & b[146])^(a[357] & b[147])^(a[356] & b[148])^(a[355] & b[149])^(a[354] & b[150])^(a[353] & b[151])^(a[352] & b[152])^(a[351] & b[153])^(a[350] & b[154])^(a[349] & b[155])^(a[348] & b[156])^(a[347] & b[157])^(a[346] & b[158])^(a[345] & b[159])^(a[344] & b[160])^(a[343] & b[161])^(a[342] & b[162])^(a[341] & b[163])^(a[340] & b[164])^(a[339] & b[165])^(a[338] & b[166])^(a[337] & b[167])^(a[336] & b[168])^(a[335] & b[169])^(a[334] & b[170])^(a[333] & b[171])^(a[332] & b[172])^(a[331] & b[173])^(a[330] & b[174])^(a[329] & b[175])^(a[328] & b[176])^(a[327] & b[177])^(a[326] & b[178])^(a[325] & b[179])^(a[324] & b[180])^(a[323] & b[181])^(a[322] & b[182])^(a[321] & b[183])^(a[320] & b[184])^(a[319] & b[185])^(a[318] & b[186])^(a[317] & b[187])^(a[316] & b[188])^(a[315] & b[189])^(a[314] & b[190])^(a[313] & b[191])^(a[312] & b[192])^(a[311] & b[193])^(a[310] & b[194])^(a[309] & b[195])^(a[308] & b[196])^(a[307] & b[197])^(a[306] & b[198])^(a[305] & b[199])^(a[304] & b[200])^(a[303] & b[201])^(a[302] & b[202])^(a[301] & b[203])^(a[300] & b[204])^(a[299] & b[205])^(a[298] & b[206])^(a[297] & b[207])^(a[296] & b[208])^(a[295] & b[209])^(a[294] & b[210])^(a[293] & b[211])^(a[292] & b[212])^(a[291] & b[213])^(a[290] & b[214])^(a[289] & b[215])^(a[288] & b[216])^(a[287] & b[217])^(a[286] & b[218])^(a[285] & b[219])^(a[284] & b[220])^(a[283] & b[221])^(a[282] & b[222])^(a[281] & b[223])^(a[280] & b[224])^(a[279] & b[225])^(a[278] & b[226])^(a[277] & b[227])^(a[276] & b[228])^(a[275] & b[229])^(a[274] & b[230])^(a[273] & b[231])^(a[272] & b[232])^(a[271] & b[233])^(a[270] & b[234])^(a[269] & b[235])^(a[268] & b[236])^(a[267] & b[237])^(a[266] & b[238])^(a[265] & b[239])^(a[264] & b[240])^(a[263] & b[241])^(a[262] & b[242])^(a[261] & b[243])^(a[260] & b[244])^(a[259] & b[245])^(a[258] & b[246])^(a[257] & b[247])^(a[256] & b[248])^(a[255] & b[249])^(a[254] & b[250])^(a[253] & b[251])^(a[252] & b[252])^(a[251] & b[253])^(a[250] & b[254])^(a[249] & b[255])^(a[248] & b[256])^(a[247] & b[257])^(a[246] & b[258])^(a[245] & b[259])^(a[244] & b[260])^(a[243] & b[261])^(a[242] & b[262])^(a[241] & b[263])^(a[240] & b[264])^(a[239] & b[265])^(a[238] & b[266])^(a[237] & b[267])^(a[236] & b[268])^(a[235] & b[269])^(a[234] & b[270])^(a[233] & b[271])^(a[232] & b[272])^(a[231] & b[273])^(a[230] & b[274])^(a[229] & b[275])^(a[228] & b[276])^(a[227] & b[277])^(a[226] & b[278])^(a[225] & b[279])^(a[224] & b[280])^(a[223] & b[281])^(a[222] & b[282])^(a[221] & b[283])^(a[220] & b[284])^(a[219] & b[285])^(a[218] & b[286])^(a[217] & b[287])^(a[216] & b[288])^(a[215] & b[289])^(a[214] & b[290])^(a[213] & b[291])^(a[212] & b[292])^(a[211] & b[293])^(a[210] & b[294])^(a[209] & b[295])^(a[208] & b[296])^(a[207] & b[297])^(a[206] & b[298])^(a[205] & b[299])^(a[204] & b[300])^(a[203] & b[301])^(a[202] & b[302])^(a[201] & b[303])^(a[200] & b[304])^(a[199] & b[305])^(a[198] & b[306])^(a[197] & b[307])^(a[196] & b[308])^(a[195] & b[309])^(a[194] & b[310])^(a[193] & b[311])^(a[192] & b[312])^(a[191] & b[313])^(a[190] & b[314])^(a[189] & b[315])^(a[188] & b[316])^(a[187] & b[317])^(a[186] & b[318])^(a[185] & b[319])^(a[184] & b[320])^(a[183] & b[321])^(a[182] & b[322])^(a[181] & b[323])^(a[180] & b[324])^(a[179] & b[325])^(a[178] & b[326])^(a[177] & b[327])^(a[176] & b[328])^(a[175] & b[329])^(a[174] & b[330])^(a[173] & b[331])^(a[172] & b[332])^(a[171] & b[333])^(a[170] & b[334])^(a[169] & b[335])^(a[168] & b[336])^(a[167] & b[337])^(a[166] & b[338])^(a[165] & b[339])^(a[164] & b[340])^(a[163] & b[341])^(a[162] & b[342])^(a[161] & b[343])^(a[160] & b[344])^(a[159] & b[345])^(a[158] & b[346])^(a[157] & b[347])^(a[156] & b[348])^(a[155] & b[349])^(a[154] & b[350])^(a[153] & b[351])^(a[152] & b[352])^(a[151] & b[353])^(a[150] & b[354])^(a[149] & b[355])^(a[148] & b[356])^(a[147] & b[357])^(a[146] & b[358])^(a[145] & b[359])^(a[144] & b[360])^(a[143] & b[361])^(a[142] & b[362])^(a[141] & b[363])^(a[140] & b[364])^(a[139] & b[365])^(a[138] & b[366])^(a[137] & b[367])^(a[136] & b[368])^(a[135] & b[369])^(a[134] & b[370])^(a[133] & b[371])^(a[132] & b[372])^(a[131] & b[373])^(a[130] & b[374])^(a[129] & b[375])^(a[128] & b[376])^(a[127] & b[377])^(a[126] & b[378])^(a[125] & b[379])^(a[124] & b[380])^(a[123] & b[381])^(a[122] & b[382])^(a[121] & b[383])^(a[120] & b[384])^(a[119] & b[385])^(a[118] & b[386])^(a[117] & b[387])^(a[116] & b[388])^(a[115] & b[389])^(a[114] & b[390])^(a[113] & b[391])^(a[112] & b[392])^(a[111] & b[393])^(a[110] & b[394])^(a[109] & b[395])^(a[108] & b[396])^(a[107] & b[397])^(a[106] & b[398])^(a[105] & b[399])^(a[104] & b[400])^(a[103] & b[401])^(a[102] & b[402])^(a[101] & b[403])^(a[100] & b[404])^(a[99] & b[405])^(a[98] & b[406])^(a[97] & b[407])^(a[96] & b[408]);
assign y[505] = (a[408] & b[97])^(a[407] & b[98])^(a[406] & b[99])^(a[405] & b[100])^(a[404] & b[101])^(a[403] & b[102])^(a[402] & b[103])^(a[401] & b[104])^(a[400] & b[105])^(a[399] & b[106])^(a[398] & b[107])^(a[397] & b[108])^(a[396] & b[109])^(a[395] & b[110])^(a[394] & b[111])^(a[393] & b[112])^(a[392] & b[113])^(a[391] & b[114])^(a[390] & b[115])^(a[389] & b[116])^(a[388] & b[117])^(a[387] & b[118])^(a[386] & b[119])^(a[385] & b[120])^(a[384] & b[121])^(a[383] & b[122])^(a[382] & b[123])^(a[381] & b[124])^(a[380] & b[125])^(a[379] & b[126])^(a[378] & b[127])^(a[377] & b[128])^(a[376] & b[129])^(a[375] & b[130])^(a[374] & b[131])^(a[373] & b[132])^(a[372] & b[133])^(a[371] & b[134])^(a[370] & b[135])^(a[369] & b[136])^(a[368] & b[137])^(a[367] & b[138])^(a[366] & b[139])^(a[365] & b[140])^(a[364] & b[141])^(a[363] & b[142])^(a[362] & b[143])^(a[361] & b[144])^(a[360] & b[145])^(a[359] & b[146])^(a[358] & b[147])^(a[357] & b[148])^(a[356] & b[149])^(a[355] & b[150])^(a[354] & b[151])^(a[353] & b[152])^(a[352] & b[153])^(a[351] & b[154])^(a[350] & b[155])^(a[349] & b[156])^(a[348] & b[157])^(a[347] & b[158])^(a[346] & b[159])^(a[345] & b[160])^(a[344] & b[161])^(a[343] & b[162])^(a[342] & b[163])^(a[341] & b[164])^(a[340] & b[165])^(a[339] & b[166])^(a[338] & b[167])^(a[337] & b[168])^(a[336] & b[169])^(a[335] & b[170])^(a[334] & b[171])^(a[333] & b[172])^(a[332] & b[173])^(a[331] & b[174])^(a[330] & b[175])^(a[329] & b[176])^(a[328] & b[177])^(a[327] & b[178])^(a[326] & b[179])^(a[325] & b[180])^(a[324] & b[181])^(a[323] & b[182])^(a[322] & b[183])^(a[321] & b[184])^(a[320] & b[185])^(a[319] & b[186])^(a[318] & b[187])^(a[317] & b[188])^(a[316] & b[189])^(a[315] & b[190])^(a[314] & b[191])^(a[313] & b[192])^(a[312] & b[193])^(a[311] & b[194])^(a[310] & b[195])^(a[309] & b[196])^(a[308] & b[197])^(a[307] & b[198])^(a[306] & b[199])^(a[305] & b[200])^(a[304] & b[201])^(a[303] & b[202])^(a[302] & b[203])^(a[301] & b[204])^(a[300] & b[205])^(a[299] & b[206])^(a[298] & b[207])^(a[297] & b[208])^(a[296] & b[209])^(a[295] & b[210])^(a[294] & b[211])^(a[293] & b[212])^(a[292] & b[213])^(a[291] & b[214])^(a[290] & b[215])^(a[289] & b[216])^(a[288] & b[217])^(a[287] & b[218])^(a[286] & b[219])^(a[285] & b[220])^(a[284] & b[221])^(a[283] & b[222])^(a[282] & b[223])^(a[281] & b[224])^(a[280] & b[225])^(a[279] & b[226])^(a[278] & b[227])^(a[277] & b[228])^(a[276] & b[229])^(a[275] & b[230])^(a[274] & b[231])^(a[273] & b[232])^(a[272] & b[233])^(a[271] & b[234])^(a[270] & b[235])^(a[269] & b[236])^(a[268] & b[237])^(a[267] & b[238])^(a[266] & b[239])^(a[265] & b[240])^(a[264] & b[241])^(a[263] & b[242])^(a[262] & b[243])^(a[261] & b[244])^(a[260] & b[245])^(a[259] & b[246])^(a[258] & b[247])^(a[257] & b[248])^(a[256] & b[249])^(a[255] & b[250])^(a[254] & b[251])^(a[253] & b[252])^(a[252] & b[253])^(a[251] & b[254])^(a[250] & b[255])^(a[249] & b[256])^(a[248] & b[257])^(a[247] & b[258])^(a[246] & b[259])^(a[245] & b[260])^(a[244] & b[261])^(a[243] & b[262])^(a[242] & b[263])^(a[241] & b[264])^(a[240] & b[265])^(a[239] & b[266])^(a[238] & b[267])^(a[237] & b[268])^(a[236] & b[269])^(a[235] & b[270])^(a[234] & b[271])^(a[233] & b[272])^(a[232] & b[273])^(a[231] & b[274])^(a[230] & b[275])^(a[229] & b[276])^(a[228] & b[277])^(a[227] & b[278])^(a[226] & b[279])^(a[225] & b[280])^(a[224] & b[281])^(a[223] & b[282])^(a[222] & b[283])^(a[221] & b[284])^(a[220] & b[285])^(a[219] & b[286])^(a[218] & b[287])^(a[217] & b[288])^(a[216] & b[289])^(a[215] & b[290])^(a[214] & b[291])^(a[213] & b[292])^(a[212] & b[293])^(a[211] & b[294])^(a[210] & b[295])^(a[209] & b[296])^(a[208] & b[297])^(a[207] & b[298])^(a[206] & b[299])^(a[205] & b[300])^(a[204] & b[301])^(a[203] & b[302])^(a[202] & b[303])^(a[201] & b[304])^(a[200] & b[305])^(a[199] & b[306])^(a[198] & b[307])^(a[197] & b[308])^(a[196] & b[309])^(a[195] & b[310])^(a[194] & b[311])^(a[193] & b[312])^(a[192] & b[313])^(a[191] & b[314])^(a[190] & b[315])^(a[189] & b[316])^(a[188] & b[317])^(a[187] & b[318])^(a[186] & b[319])^(a[185] & b[320])^(a[184] & b[321])^(a[183] & b[322])^(a[182] & b[323])^(a[181] & b[324])^(a[180] & b[325])^(a[179] & b[326])^(a[178] & b[327])^(a[177] & b[328])^(a[176] & b[329])^(a[175] & b[330])^(a[174] & b[331])^(a[173] & b[332])^(a[172] & b[333])^(a[171] & b[334])^(a[170] & b[335])^(a[169] & b[336])^(a[168] & b[337])^(a[167] & b[338])^(a[166] & b[339])^(a[165] & b[340])^(a[164] & b[341])^(a[163] & b[342])^(a[162] & b[343])^(a[161] & b[344])^(a[160] & b[345])^(a[159] & b[346])^(a[158] & b[347])^(a[157] & b[348])^(a[156] & b[349])^(a[155] & b[350])^(a[154] & b[351])^(a[153] & b[352])^(a[152] & b[353])^(a[151] & b[354])^(a[150] & b[355])^(a[149] & b[356])^(a[148] & b[357])^(a[147] & b[358])^(a[146] & b[359])^(a[145] & b[360])^(a[144] & b[361])^(a[143] & b[362])^(a[142] & b[363])^(a[141] & b[364])^(a[140] & b[365])^(a[139] & b[366])^(a[138] & b[367])^(a[137] & b[368])^(a[136] & b[369])^(a[135] & b[370])^(a[134] & b[371])^(a[133] & b[372])^(a[132] & b[373])^(a[131] & b[374])^(a[130] & b[375])^(a[129] & b[376])^(a[128] & b[377])^(a[127] & b[378])^(a[126] & b[379])^(a[125] & b[380])^(a[124] & b[381])^(a[123] & b[382])^(a[122] & b[383])^(a[121] & b[384])^(a[120] & b[385])^(a[119] & b[386])^(a[118] & b[387])^(a[117] & b[388])^(a[116] & b[389])^(a[115] & b[390])^(a[114] & b[391])^(a[113] & b[392])^(a[112] & b[393])^(a[111] & b[394])^(a[110] & b[395])^(a[109] & b[396])^(a[108] & b[397])^(a[107] & b[398])^(a[106] & b[399])^(a[105] & b[400])^(a[104] & b[401])^(a[103] & b[402])^(a[102] & b[403])^(a[101] & b[404])^(a[100] & b[405])^(a[99] & b[406])^(a[98] & b[407])^(a[97] & b[408]);
assign y[506] = (a[408] & b[98])^(a[407] & b[99])^(a[406] & b[100])^(a[405] & b[101])^(a[404] & b[102])^(a[403] & b[103])^(a[402] & b[104])^(a[401] & b[105])^(a[400] & b[106])^(a[399] & b[107])^(a[398] & b[108])^(a[397] & b[109])^(a[396] & b[110])^(a[395] & b[111])^(a[394] & b[112])^(a[393] & b[113])^(a[392] & b[114])^(a[391] & b[115])^(a[390] & b[116])^(a[389] & b[117])^(a[388] & b[118])^(a[387] & b[119])^(a[386] & b[120])^(a[385] & b[121])^(a[384] & b[122])^(a[383] & b[123])^(a[382] & b[124])^(a[381] & b[125])^(a[380] & b[126])^(a[379] & b[127])^(a[378] & b[128])^(a[377] & b[129])^(a[376] & b[130])^(a[375] & b[131])^(a[374] & b[132])^(a[373] & b[133])^(a[372] & b[134])^(a[371] & b[135])^(a[370] & b[136])^(a[369] & b[137])^(a[368] & b[138])^(a[367] & b[139])^(a[366] & b[140])^(a[365] & b[141])^(a[364] & b[142])^(a[363] & b[143])^(a[362] & b[144])^(a[361] & b[145])^(a[360] & b[146])^(a[359] & b[147])^(a[358] & b[148])^(a[357] & b[149])^(a[356] & b[150])^(a[355] & b[151])^(a[354] & b[152])^(a[353] & b[153])^(a[352] & b[154])^(a[351] & b[155])^(a[350] & b[156])^(a[349] & b[157])^(a[348] & b[158])^(a[347] & b[159])^(a[346] & b[160])^(a[345] & b[161])^(a[344] & b[162])^(a[343] & b[163])^(a[342] & b[164])^(a[341] & b[165])^(a[340] & b[166])^(a[339] & b[167])^(a[338] & b[168])^(a[337] & b[169])^(a[336] & b[170])^(a[335] & b[171])^(a[334] & b[172])^(a[333] & b[173])^(a[332] & b[174])^(a[331] & b[175])^(a[330] & b[176])^(a[329] & b[177])^(a[328] & b[178])^(a[327] & b[179])^(a[326] & b[180])^(a[325] & b[181])^(a[324] & b[182])^(a[323] & b[183])^(a[322] & b[184])^(a[321] & b[185])^(a[320] & b[186])^(a[319] & b[187])^(a[318] & b[188])^(a[317] & b[189])^(a[316] & b[190])^(a[315] & b[191])^(a[314] & b[192])^(a[313] & b[193])^(a[312] & b[194])^(a[311] & b[195])^(a[310] & b[196])^(a[309] & b[197])^(a[308] & b[198])^(a[307] & b[199])^(a[306] & b[200])^(a[305] & b[201])^(a[304] & b[202])^(a[303] & b[203])^(a[302] & b[204])^(a[301] & b[205])^(a[300] & b[206])^(a[299] & b[207])^(a[298] & b[208])^(a[297] & b[209])^(a[296] & b[210])^(a[295] & b[211])^(a[294] & b[212])^(a[293] & b[213])^(a[292] & b[214])^(a[291] & b[215])^(a[290] & b[216])^(a[289] & b[217])^(a[288] & b[218])^(a[287] & b[219])^(a[286] & b[220])^(a[285] & b[221])^(a[284] & b[222])^(a[283] & b[223])^(a[282] & b[224])^(a[281] & b[225])^(a[280] & b[226])^(a[279] & b[227])^(a[278] & b[228])^(a[277] & b[229])^(a[276] & b[230])^(a[275] & b[231])^(a[274] & b[232])^(a[273] & b[233])^(a[272] & b[234])^(a[271] & b[235])^(a[270] & b[236])^(a[269] & b[237])^(a[268] & b[238])^(a[267] & b[239])^(a[266] & b[240])^(a[265] & b[241])^(a[264] & b[242])^(a[263] & b[243])^(a[262] & b[244])^(a[261] & b[245])^(a[260] & b[246])^(a[259] & b[247])^(a[258] & b[248])^(a[257] & b[249])^(a[256] & b[250])^(a[255] & b[251])^(a[254] & b[252])^(a[253] & b[253])^(a[252] & b[254])^(a[251] & b[255])^(a[250] & b[256])^(a[249] & b[257])^(a[248] & b[258])^(a[247] & b[259])^(a[246] & b[260])^(a[245] & b[261])^(a[244] & b[262])^(a[243] & b[263])^(a[242] & b[264])^(a[241] & b[265])^(a[240] & b[266])^(a[239] & b[267])^(a[238] & b[268])^(a[237] & b[269])^(a[236] & b[270])^(a[235] & b[271])^(a[234] & b[272])^(a[233] & b[273])^(a[232] & b[274])^(a[231] & b[275])^(a[230] & b[276])^(a[229] & b[277])^(a[228] & b[278])^(a[227] & b[279])^(a[226] & b[280])^(a[225] & b[281])^(a[224] & b[282])^(a[223] & b[283])^(a[222] & b[284])^(a[221] & b[285])^(a[220] & b[286])^(a[219] & b[287])^(a[218] & b[288])^(a[217] & b[289])^(a[216] & b[290])^(a[215] & b[291])^(a[214] & b[292])^(a[213] & b[293])^(a[212] & b[294])^(a[211] & b[295])^(a[210] & b[296])^(a[209] & b[297])^(a[208] & b[298])^(a[207] & b[299])^(a[206] & b[300])^(a[205] & b[301])^(a[204] & b[302])^(a[203] & b[303])^(a[202] & b[304])^(a[201] & b[305])^(a[200] & b[306])^(a[199] & b[307])^(a[198] & b[308])^(a[197] & b[309])^(a[196] & b[310])^(a[195] & b[311])^(a[194] & b[312])^(a[193] & b[313])^(a[192] & b[314])^(a[191] & b[315])^(a[190] & b[316])^(a[189] & b[317])^(a[188] & b[318])^(a[187] & b[319])^(a[186] & b[320])^(a[185] & b[321])^(a[184] & b[322])^(a[183] & b[323])^(a[182] & b[324])^(a[181] & b[325])^(a[180] & b[326])^(a[179] & b[327])^(a[178] & b[328])^(a[177] & b[329])^(a[176] & b[330])^(a[175] & b[331])^(a[174] & b[332])^(a[173] & b[333])^(a[172] & b[334])^(a[171] & b[335])^(a[170] & b[336])^(a[169] & b[337])^(a[168] & b[338])^(a[167] & b[339])^(a[166] & b[340])^(a[165] & b[341])^(a[164] & b[342])^(a[163] & b[343])^(a[162] & b[344])^(a[161] & b[345])^(a[160] & b[346])^(a[159] & b[347])^(a[158] & b[348])^(a[157] & b[349])^(a[156] & b[350])^(a[155] & b[351])^(a[154] & b[352])^(a[153] & b[353])^(a[152] & b[354])^(a[151] & b[355])^(a[150] & b[356])^(a[149] & b[357])^(a[148] & b[358])^(a[147] & b[359])^(a[146] & b[360])^(a[145] & b[361])^(a[144] & b[362])^(a[143] & b[363])^(a[142] & b[364])^(a[141] & b[365])^(a[140] & b[366])^(a[139] & b[367])^(a[138] & b[368])^(a[137] & b[369])^(a[136] & b[370])^(a[135] & b[371])^(a[134] & b[372])^(a[133] & b[373])^(a[132] & b[374])^(a[131] & b[375])^(a[130] & b[376])^(a[129] & b[377])^(a[128] & b[378])^(a[127] & b[379])^(a[126] & b[380])^(a[125] & b[381])^(a[124] & b[382])^(a[123] & b[383])^(a[122] & b[384])^(a[121] & b[385])^(a[120] & b[386])^(a[119] & b[387])^(a[118] & b[388])^(a[117] & b[389])^(a[116] & b[390])^(a[115] & b[391])^(a[114] & b[392])^(a[113] & b[393])^(a[112] & b[394])^(a[111] & b[395])^(a[110] & b[396])^(a[109] & b[397])^(a[108] & b[398])^(a[107] & b[399])^(a[106] & b[400])^(a[105] & b[401])^(a[104] & b[402])^(a[103] & b[403])^(a[102] & b[404])^(a[101] & b[405])^(a[100] & b[406])^(a[99] & b[407])^(a[98] & b[408]);
assign y[507] = (a[408] & b[99])^(a[407] & b[100])^(a[406] & b[101])^(a[405] & b[102])^(a[404] & b[103])^(a[403] & b[104])^(a[402] & b[105])^(a[401] & b[106])^(a[400] & b[107])^(a[399] & b[108])^(a[398] & b[109])^(a[397] & b[110])^(a[396] & b[111])^(a[395] & b[112])^(a[394] & b[113])^(a[393] & b[114])^(a[392] & b[115])^(a[391] & b[116])^(a[390] & b[117])^(a[389] & b[118])^(a[388] & b[119])^(a[387] & b[120])^(a[386] & b[121])^(a[385] & b[122])^(a[384] & b[123])^(a[383] & b[124])^(a[382] & b[125])^(a[381] & b[126])^(a[380] & b[127])^(a[379] & b[128])^(a[378] & b[129])^(a[377] & b[130])^(a[376] & b[131])^(a[375] & b[132])^(a[374] & b[133])^(a[373] & b[134])^(a[372] & b[135])^(a[371] & b[136])^(a[370] & b[137])^(a[369] & b[138])^(a[368] & b[139])^(a[367] & b[140])^(a[366] & b[141])^(a[365] & b[142])^(a[364] & b[143])^(a[363] & b[144])^(a[362] & b[145])^(a[361] & b[146])^(a[360] & b[147])^(a[359] & b[148])^(a[358] & b[149])^(a[357] & b[150])^(a[356] & b[151])^(a[355] & b[152])^(a[354] & b[153])^(a[353] & b[154])^(a[352] & b[155])^(a[351] & b[156])^(a[350] & b[157])^(a[349] & b[158])^(a[348] & b[159])^(a[347] & b[160])^(a[346] & b[161])^(a[345] & b[162])^(a[344] & b[163])^(a[343] & b[164])^(a[342] & b[165])^(a[341] & b[166])^(a[340] & b[167])^(a[339] & b[168])^(a[338] & b[169])^(a[337] & b[170])^(a[336] & b[171])^(a[335] & b[172])^(a[334] & b[173])^(a[333] & b[174])^(a[332] & b[175])^(a[331] & b[176])^(a[330] & b[177])^(a[329] & b[178])^(a[328] & b[179])^(a[327] & b[180])^(a[326] & b[181])^(a[325] & b[182])^(a[324] & b[183])^(a[323] & b[184])^(a[322] & b[185])^(a[321] & b[186])^(a[320] & b[187])^(a[319] & b[188])^(a[318] & b[189])^(a[317] & b[190])^(a[316] & b[191])^(a[315] & b[192])^(a[314] & b[193])^(a[313] & b[194])^(a[312] & b[195])^(a[311] & b[196])^(a[310] & b[197])^(a[309] & b[198])^(a[308] & b[199])^(a[307] & b[200])^(a[306] & b[201])^(a[305] & b[202])^(a[304] & b[203])^(a[303] & b[204])^(a[302] & b[205])^(a[301] & b[206])^(a[300] & b[207])^(a[299] & b[208])^(a[298] & b[209])^(a[297] & b[210])^(a[296] & b[211])^(a[295] & b[212])^(a[294] & b[213])^(a[293] & b[214])^(a[292] & b[215])^(a[291] & b[216])^(a[290] & b[217])^(a[289] & b[218])^(a[288] & b[219])^(a[287] & b[220])^(a[286] & b[221])^(a[285] & b[222])^(a[284] & b[223])^(a[283] & b[224])^(a[282] & b[225])^(a[281] & b[226])^(a[280] & b[227])^(a[279] & b[228])^(a[278] & b[229])^(a[277] & b[230])^(a[276] & b[231])^(a[275] & b[232])^(a[274] & b[233])^(a[273] & b[234])^(a[272] & b[235])^(a[271] & b[236])^(a[270] & b[237])^(a[269] & b[238])^(a[268] & b[239])^(a[267] & b[240])^(a[266] & b[241])^(a[265] & b[242])^(a[264] & b[243])^(a[263] & b[244])^(a[262] & b[245])^(a[261] & b[246])^(a[260] & b[247])^(a[259] & b[248])^(a[258] & b[249])^(a[257] & b[250])^(a[256] & b[251])^(a[255] & b[252])^(a[254] & b[253])^(a[253] & b[254])^(a[252] & b[255])^(a[251] & b[256])^(a[250] & b[257])^(a[249] & b[258])^(a[248] & b[259])^(a[247] & b[260])^(a[246] & b[261])^(a[245] & b[262])^(a[244] & b[263])^(a[243] & b[264])^(a[242] & b[265])^(a[241] & b[266])^(a[240] & b[267])^(a[239] & b[268])^(a[238] & b[269])^(a[237] & b[270])^(a[236] & b[271])^(a[235] & b[272])^(a[234] & b[273])^(a[233] & b[274])^(a[232] & b[275])^(a[231] & b[276])^(a[230] & b[277])^(a[229] & b[278])^(a[228] & b[279])^(a[227] & b[280])^(a[226] & b[281])^(a[225] & b[282])^(a[224] & b[283])^(a[223] & b[284])^(a[222] & b[285])^(a[221] & b[286])^(a[220] & b[287])^(a[219] & b[288])^(a[218] & b[289])^(a[217] & b[290])^(a[216] & b[291])^(a[215] & b[292])^(a[214] & b[293])^(a[213] & b[294])^(a[212] & b[295])^(a[211] & b[296])^(a[210] & b[297])^(a[209] & b[298])^(a[208] & b[299])^(a[207] & b[300])^(a[206] & b[301])^(a[205] & b[302])^(a[204] & b[303])^(a[203] & b[304])^(a[202] & b[305])^(a[201] & b[306])^(a[200] & b[307])^(a[199] & b[308])^(a[198] & b[309])^(a[197] & b[310])^(a[196] & b[311])^(a[195] & b[312])^(a[194] & b[313])^(a[193] & b[314])^(a[192] & b[315])^(a[191] & b[316])^(a[190] & b[317])^(a[189] & b[318])^(a[188] & b[319])^(a[187] & b[320])^(a[186] & b[321])^(a[185] & b[322])^(a[184] & b[323])^(a[183] & b[324])^(a[182] & b[325])^(a[181] & b[326])^(a[180] & b[327])^(a[179] & b[328])^(a[178] & b[329])^(a[177] & b[330])^(a[176] & b[331])^(a[175] & b[332])^(a[174] & b[333])^(a[173] & b[334])^(a[172] & b[335])^(a[171] & b[336])^(a[170] & b[337])^(a[169] & b[338])^(a[168] & b[339])^(a[167] & b[340])^(a[166] & b[341])^(a[165] & b[342])^(a[164] & b[343])^(a[163] & b[344])^(a[162] & b[345])^(a[161] & b[346])^(a[160] & b[347])^(a[159] & b[348])^(a[158] & b[349])^(a[157] & b[350])^(a[156] & b[351])^(a[155] & b[352])^(a[154] & b[353])^(a[153] & b[354])^(a[152] & b[355])^(a[151] & b[356])^(a[150] & b[357])^(a[149] & b[358])^(a[148] & b[359])^(a[147] & b[360])^(a[146] & b[361])^(a[145] & b[362])^(a[144] & b[363])^(a[143] & b[364])^(a[142] & b[365])^(a[141] & b[366])^(a[140] & b[367])^(a[139] & b[368])^(a[138] & b[369])^(a[137] & b[370])^(a[136] & b[371])^(a[135] & b[372])^(a[134] & b[373])^(a[133] & b[374])^(a[132] & b[375])^(a[131] & b[376])^(a[130] & b[377])^(a[129] & b[378])^(a[128] & b[379])^(a[127] & b[380])^(a[126] & b[381])^(a[125] & b[382])^(a[124] & b[383])^(a[123] & b[384])^(a[122] & b[385])^(a[121] & b[386])^(a[120] & b[387])^(a[119] & b[388])^(a[118] & b[389])^(a[117] & b[390])^(a[116] & b[391])^(a[115] & b[392])^(a[114] & b[393])^(a[113] & b[394])^(a[112] & b[395])^(a[111] & b[396])^(a[110] & b[397])^(a[109] & b[398])^(a[108] & b[399])^(a[107] & b[400])^(a[106] & b[401])^(a[105] & b[402])^(a[104] & b[403])^(a[103] & b[404])^(a[102] & b[405])^(a[101] & b[406])^(a[100] & b[407])^(a[99] & b[408]);
assign y[508] = (a[408] & b[100])^(a[407] & b[101])^(a[406] & b[102])^(a[405] & b[103])^(a[404] & b[104])^(a[403] & b[105])^(a[402] & b[106])^(a[401] & b[107])^(a[400] & b[108])^(a[399] & b[109])^(a[398] & b[110])^(a[397] & b[111])^(a[396] & b[112])^(a[395] & b[113])^(a[394] & b[114])^(a[393] & b[115])^(a[392] & b[116])^(a[391] & b[117])^(a[390] & b[118])^(a[389] & b[119])^(a[388] & b[120])^(a[387] & b[121])^(a[386] & b[122])^(a[385] & b[123])^(a[384] & b[124])^(a[383] & b[125])^(a[382] & b[126])^(a[381] & b[127])^(a[380] & b[128])^(a[379] & b[129])^(a[378] & b[130])^(a[377] & b[131])^(a[376] & b[132])^(a[375] & b[133])^(a[374] & b[134])^(a[373] & b[135])^(a[372] & b[136])^(a[371] & b[137])^(a[370] & b[138])^(a[369] & b[139])^(a[368] & b[140])^(a[367] & b[141])^(a[366] & b[142])^(a[365] & b[143])^(a[364] & b[144])^(a[363] & b[145])^(a[362] & b[146])^(a[361] & b[147])^(a[360] & b[148])^(a[359] & b[149])^(a[358] & b[150])^(a[357] & b[151])^(a[356] & b[152])^(a[355] & b[153])^(a[354] & b[154])^(a[353] & b[155])^(a[352] & b[156])^(a[351] & b[157])^(a[350] & b[158])^(a[349] & b[159])^(a[348] & b[160])^(a[347] & b[161])^(a[346] & b[162])^(a[345] & b[163])^(a[344] & b[164])^(a[343] & b[165])^(a[342] & b[166])^(a[341] & b[167])^(a[340] & b[168])^(a[339] & b[169])^(a[338] & b[170])^(a[337] & b[171])^(a[336] & b[172])^(a[335] & b[173])^(a[334] & b[174])^(a[333] & b[175])^(a[332] & b[176])^(a[331] & b[177])^(a[330] & b[178])^(a[329] & b[179])^(a[328] & b[180])^(a[327] & b[181])^(a[326] & b[182])^(a[325] & b[183])^(a[324] & b[184])^(a[323] & b[185])^(a[322] & b[186])^(a[321] & b[187])^(a[320] & b[188])^(a[319] & b[189])^(a[318] & b[190])^(a[317] & b[191])^(a[316] & b[192])^(a[315] & b[193])^(a[314] & b[194])^(a[313] & b[195])^(a[312] & b[196])^(a[311] & b[197])^(a[310] & b[198])^(a[309] & b[199])^(a[308] & b[200])^(a[307] & b[201])^(a[306] & b[202])^(a[305] & b[203])^(a[304] & b[204])^(a[303] & b[205])^(a[302] & b[206])^(a[301] & b[207])^(a[300] & b[208])^(a[299] & b[209])^(a[298] & b[210])^(a[297] & b[211])^(a[296] & b[212])^(a[295] & b[213])^(a[294] & b[214])^(a[293] & b[215])^(a[292] & b[216])^(a[291] & b[217])^(a[290] & b[218])^(a[289] & b[219])^(a[288] & b[220])^(a[287] & b[221])^(a[286] & b[222])^(a[285] & b[223])^(a[284] & b[224])^(a[283] & b[225])^(a[282] & b[226])^(a[281] & b[227])^(a[280] & b[228])^(a[279] & b[229])^(a[278] & b[230])^(a[277] & b[231])^(a[276] & b[232])^(a[275] & b[233])^(a[274] & b[234])^(a[273] & b[235])^(a[272] & b[236])^(a[271] & b[237])^(a[270] & b[238])^(a[269] & b[239])^(a[268] & b[240])^(a[267] & b[241])^(a[266] & b[242])^(a[265] & b[243])^(a[264] & b[244])^(a[263] & b[245])^(a[262] & b[246])^(a[261] & b[247])^(a[260] & b[248])^(a[259] & b[249])^(a[258] & b[250])^(a[257] & b[251])^(a[256] & b[252])^(a[255] & b[253])^(a[254] & b[254])^(a[253] & b[255])^(a[252] & b[256])^(a[251] & b[257])^(a[250] & b[258])^(a[249] & b[259])^(a[248] & b[260])^(a[247] & b[261])^(a[246] & b[262])^(a[245] & b[263])^(a[244] & b[264])^(a[243] & b[265])^(a[242] & b[266])^(a[241] & b[267])^(a[240] & b[268])^(a[239] & b[269])^(a[238] & b[270])^(a[237] & b[271])^(a[236] & b[272])^(a[235] & b[273])^(a[234] & b[274])^(a[233] & b[275])^(a[232] & b[276])^(a[231] & b[277])^(a[230] & b[278])^(a[229] & b[279])^(a[228] & b[280])^(a[227] & b[281])^(a[226] & b[282])^(a[225] & b[283])^(a[224] & b[284])^(a[223] & b[285])^(a[222] & b[286])^(a[221] & b[287])^(a[220] & b[288])^(a[219] & b[289])^(a[218] & b[290])^(a[217] & b[291])^(a[216] & b[292])^(a[215] & b[293])^(a[214] & b[294])^(a[213] & b[295])^(a[212] & b[296])^(a[211] & b[297])^(a[210] & b[298])^(a[209] & b[299])^(a[208] & b[300])^(a[207] & b[301])^(a[206] & b[302])^(a[205] & b[303])^(a[204] & b[304])^(a[203] & b[305])^(a[202] & b[306])^(a[201] & b[307])^(a[200] & b[308])^(a[199] & b[309])^(a[198] & b[310])^(a[197] & b[311])^(a[196] & b[312])^(a[195] & b[313])^(a[194] & b[314])^(a[193] & b[315])^(a[192] & b[316])^(a[191] & b[317])^(a[190] & b[318])^(a[189] & b[319])^(a[188] & b[320])^(a[187] & b[321])^(a[186] & b[322])^(a[185] & b[323])^(a[184] & b[324])^(a[183] & b[325])^(a[182] & b[326])^(a[181] & b[327])^(a[180] & b[328])^(a[179] & b[329])^(a[178] & b[330])^(a[177] & b[331])^(a[176] & b[332])^(a[175] & b[333])^(a[174] & b[334])^(a[173] & b[335])^(a[172] & b[336])^(a[171] & b[337])^(a[170] & b[338])^(a[169] & b[339])^(a[168] & b[340])^(a[167] & b[341])^(a[166] & b[342])^(a[165] & b[343])^(a[164] & b[344])^(a[163] & b[345])^(a[162] & b[346])^(a[161] & b[347])^(a[160] & b[348])^(a[159] & b[349])^(a[158] & b[350])^(a[157] & b[351])^(a[156] & b[352])^(a[155] & b[353])^(a[154] & b[354])^(a[153] & b[355])^(a[152] & b[356])^(a[151] & b[357])^(a[150] & b[358])^(a[149] & b[359])^(a[148] & b[360])^(a[147] & b[361])^(a[146] & b[362])^(a[145] & b[363])^(a[144] & b[364])^(a[143] & b[365])^(a[142] & b[366])^(a[141] & b[367])^(a[140] & b[368])^(a[139] & b[369])^(a[138] & b[370])^(a[137] & b[371])^(a[136] & b[372])^(a[135] & b[373])^(a[134] & b[374])^(a[133] & b[375])^(a[132] & b[376])^(a[131] & b[377])^(a[130] & b[378])^(a[129] & b[379])^(a[128] & b[380])^(a[127] & b[381])^(a[126] & b[382])^(a[125] & b[383])^(a[124] & b[384])^(a[123] & b[385])^(a[122] & b[386])^(a[121] & b[387])^(a[120] & b[388])^(a[119] & b[389])^(a[118] & b[390])^(a[117] & b[391])^(a[116] & b[392])^(a[115] & b[393])^(a[114] & b[394])^(a[113] & b[395])^(a[112] & b[396])^(a[111] & b[397])^(a[110] & b[398])^(a[109] & b[399])^(a[108] & b[400])^(a[107] & b[401])^(a[106] & b[402])^(a[105] & b[403])^(a[104] & b[404])^(a[103] & b[405])^(a[102] & b[406])^(a[101] & b[407])^(a[100] & b[408]);
assign y[509] = (a[408] & b[101])^(a[407] & b[102])^(a[406] & b[103])^(a[405] & b[104])^(a[404] & b[105])^(a[403] & b[106])^(a[402] & b[107])^(a[401] & b[108])^(a[400] & b[109])^(a[399] & b[110])^(a[398] & b[111])^(a[397] & b[112])^(a[396] & b[113])^(a[395] & b[114])^(a[394] & b[115])^(a[393] & b[116])^(a[392] & b[117])^(a[391] & b[118])^(a[390] & b[119])^(a[389] & b[120])^(a[388] & b[121])^(a[387] & b[122])^(a[386] & b[123])^(a[385] & b[124])^(a[384] & b[125])^(a[383] & b[126])^(a[382] & b[127])^(a[381] & b[128])^(a[380] & b[129])^(a[379] & b[130])^(a[378] & b[131])^(a[377] & b[132])^(a[376] & b[133])^(a[375] & b[134])^(a[374] & b[135])^(a[373] & b[136])^(a[372] & b[137])^(a[371] & b[138])^(a[370] & b[139])^(a[369] & b[140])^(a[368] & b[141])^(a[367] & b[142])^(a[366] & b[143])^(a[365] & b[144])^(a[364] & b[145])^(a[363] & b[146])^(a[362] & b[147])^(a[361] & b[148])^(a[360] & b[149])^(a[359] & b[150])^(a[358] & b[151])^(a[357] & b[152])^(a[356] & b[153])^(a[355] & b[154])^(a[354] & b[155])^(a[353] & b[156])^(a[352] & b[157])^(a[351] & b[158])^(a[350] & b[159])^(a[349] & b[160])^(a[348] & b[161])^(a[347] & b[162])^(a[346] & b[163])^(a[345] & b[164])^(a[344] & b[165])^(a[343] & b[166])^(a[342] & b[167])^(a[341] & b[168])^(a[340] & b[169])^(a[339] & b[170])^(a[338] & b[171])^(a[337] & b[172])^(a[336] & b[173])^(a[335] & b[174])^(a[334] & b[175])^(a[333] & b[176])^(a[332] & b[177])^(a[331] & b[178])^(a[330] & b[179])^(a[329] & b[180])^(a[328] & b[181])^(a[327] & b[182])^(a[326] & b[183])^(a[325] & b[184])^(a[324] & b[185])^(a[323] & b[186])^(a[322] & b[187])^(a[321] & b[188])^(a[320] & b[189])^(a[319] & b[190])^(a[318] & b[191])^(a[317] & b[192])^(a[316] & b[193])^(a[315] & b[194])^(a[314] & b[195])^(a[313] & b[196])^(a[312] & b[197])^(a[311] & b[198])^(a[310] & b[199])^(a[309] & b[200])^(a[308] & b[201])^(a[307] & b[202])^(a[306] & b[203])^(a[305] & b[204])^(a[304] & b[205])^(a[303] & b[206])^(a[302] & b[207])^(a[301] & b[208])^(a[300] & b[209])^(a[299] & b[210])^(a[298] & b[211])^(a[297] & b[212])^(a[296] & b[213])^(a[295] & b[214])^(a[294] & b[215])^(a[293] & b[216])^(a[292] & b[217])^(a[291] & b[218])^(a[290] & b[219])^(a[289] & b[220])^(a[288] & b[221])^(a[287] & b[222])^(a[286] & b[223])^(a[285] & b[224])^(a[284] & b[225])^(a[283] & b[226])^(a[282] & b[227])^(a[281] & b[228])^(a[280] & b[229])^(a[279] & b[230])^(a[278] & b[231])^(a[277] & b[232])^(a[276] & b[233])^(a[275] & b[234])^(a[274] & b[235])^(a[273] & b[236])^(a[272] & b[237])^(a[271] & b[238])^(a[270] & b[239])^(a[269] & b[240])^(a[268] & b[241])^(a[267] & b[242])^(a[266] & b[243])^(a[265] & b[244])^(a[264] & b[245])^(a[263] & b[246])^(a[262] & b[247])^(a[261] & b[248])^(a[260] & b[249])^(a[259] & b[250])^(a[258] & b[251])^(a[257] & b[252])^(a[256] & b[253])^(a[255] & b[254])^(a[254] & b[255])^(a[253] & b[256])^(a[252] & b[257])^(a[251] & b[258])^(a[250] & b[259])^(a[249] & b[260])^(a[248] & b[261])^(a[247] & b[262])^(a[246] & b[263])^(a[245] & b[264])^(a[244] & b[265])^(a[243] & b[266])^(a[242] & b[267])^(a[241] & b[268])^(a[240] & b[269])^(a[239] & b[270])^(a[238] & b[271])^(a[237] & b[272])^(a[236] & b[273])^(a[235] & b[274])^(a[234] & b[275])^(a[233] & b[276])^(a[232] & b[277])^(a[231] & b[278])^(a[230] & b[279])^(a[229] & b[280])^(a[228] & b[281])^(a[227] & b[282])^(a[226] & b[283])^(a[225] & b[284])^(a[224] & b[285])^(a[223] & b[286])^(a[222] & b[287])^(a[221] & b[288])^(a[220] & b[289])^(a[219] & b[290])^(a[218] & b[291])^(a[217] & b[292])^(a[216] & b[293])^(a[215] & b[294])^(a[214] & b[295])^(a[213] & b[296])^(a[212] & b[297])^(a[211] & b[298])^(a[210] & b[299])^(a[209] & b[300])^(a[208] & b[301])^(a[207] & b[302])^(a[206] & b[303])^(a[205] & b[304])^(a[204] & b[305])^(a[203] & b[306])^(a[202] & b[307])^(a[201] & b[308])^(a[200] & b[309])^(a[199] & b[310])^(a[198] & b[311])^(a[197] & b[312])^(a[196] & b[313])^(a[195] & b[314])^(a[194] & b[315])^(a[193] & b[316])^(a[192] & b[317])^(a[191] & b[318])^(a[190] & b[319])^(a[189] & b[320])^(a[188] & b[321])^(a[187] & b[322])^(a[186] & b[323])^(a[185] & b[324])^(a[184] & b[325])^(a[183] & b[326])^(a[182] & b[327])^(a[181] & b[328])^(a[180] & b[329])^(a[179] & b[330])^(a[178] & b[331])^(a[177] & b[332])^(a[176] & b[333])^(a[175] & b[334])^(a[174] & b[335])^(a[173] & b[336])^(a[172] & b[337])^(a[171] & b[338])^(a[170] & b[339])^(a[169] & b[340])^(a[168] & b[341])^(a[167] & b[342])^(a[166] & b[343])^(a[165] & b[344])^(a[164] & b[345])^(a[163] & b[346])^(a[162] & b[347])^(a[161] & b[348])^(a[160] & b[349])^(a[159] & b[350])^(a[158] & b[351])^(a[157] & b[352])^(a[156] & b[353])^(a[155] & b[354])^(a[154] & b[355])^(a[153] & b[356])^(a[152] & b[357])^(a[151] & b[358])^(a[150] & b[359])^(a[149] & b[360])^(a[148] & b[361])^(a[147] & b[362])^(a[146] & b[363])^(a[145] & b[364])^(a[144] & b[365])^(a[143] & b[366])^(a[142] & b[367])^(a[141] & b[368])^(a[140] & b[369])^(a[139] & b[370])^(a[138] & b[371])^(a[137] & b[372])^(a[136] & b[373])^(a[135] & b[374])^(a[134] & b[375])^(a[133] & b[376])^(a[132] & b[377])^(a[131] & b[378])^(a[130] & b[379])^(a[129] & b[380])^(a[128] & b[381])^(a[127] & b[382])^(a[126] & b[383])^(a[125] & b[384])^(a[124] & b[385])^(a[123] & b[386])^(a[122] & b[387])^(a[121] & b[388])^(a[120] & b[389])^(a[119] & b[390])^(a[118] & b[391])^(a[117] & b[392])^(a[116] & b[393])^(a[115] & b[394])^(a[114] & b[395])^(a[113] & b[396])^(a[112] & b[397])^(a[111] & b[398])^(a[110] & b[399])^(a[109] & b[400])^(a[108] & b[401])^(a[107] & b[402])^(a[106] & b[403])^(a[105] & b[404])^(a[104] & b[405])^(a[103] & b[406])^(a[102] & b[407])^(a[101] & b[408]);
assign y[510] = (a[408] & b[102])^(a[407] & b[103])^(a[406] & b[104])^(a[405] & b[105])^(a[404] & b[106])^(a[403] & b[107])^(a[402] & b[108])^(a[401] & b[109])^(a[400] & b[110])^(a[399] & b[111])^(a[398] & b[112])^(a[397] & b[113])^(a[396] & b[114])^(a[395] & b[115])^(a[394] & b[116])^(a[393] & b[117])^(a[392] & b[118])^(a[391] & b[119])^(a[390] & b[120])^(a[389] & b[121])^(a[388] & b[122])^(a[387] & b[123])^(a[386] & b[124])^(a[385] & b[125])^(a[384] & b[126])^(a[383] & b[127])^(a[382] & b[128])^(a[381] & b[129])^(a[380] & b[130])^(a[379] & b[131])^(a[378] & b[132])^(a[377] & b[133])^(a[376] & b[134])^(a[375] & b[135])^(a[374] & b[136])^(a[373] & b[137])^(a[372] & b[138])^(a[371] & b[139])^(a[370] & b[140])^(a[369] & b[141])^(a[368] & b[142])^(a[367] & b[143])^(a[366] & b[144])^(a[365] & b[145])^(a[364] & b[146])^(a[363] & b[147])^(a[362] & b[148])^(a[361] & b[149])^(a[360] & b[150])^(a[359] & b[151])^(a[358] & b[152])^(a[357] & b[153])^(a[356] & b[154])^(a[355] & b[155])^(a[354] & b[156])^(a[353] & b[157])^(a[352] & b[158])^(a[351] & b[159])^(a[350] & b[160])^(a[349] & b[161])^(a[348] & b[162])^(a[347] & b[163])^(a[346] & b[164])^(a[345] & b[165])^(a[344] & b[166])^(a[343] & b[167])^(a[342] & b[168])^(a[341] & b[169])^(a[340] & b[170])^(a[339] & b[171])^(a[338] & b[172])^(a[337] & b[173])^(a[336] & b[174])^(a[335] & b[175])^(a[334] & b[176])^(a[333] & b[177])^(a[332] & b[178])^(a[331] & b[179])^(a[330] & b[180])^(a[329] & b[181])^(a[328] & b[182])^(a[327] & b[183])^(a[326] & b[184])^(a[325] & b[185])^(a[324] & b[186])^(a[323] & b[187])^(a[322] & b[188])^(a[321] & b[189])^(a[320] & b[190])^(a[319] & b[191])^(a[318] & b[192])^(a[317] & b[193])^(a[316] & b[194])^(a[315] & b[195])^(a[314] & b[196])^(a[313] & b[197])^(a[312] & b[198])^(a[311] & b[199])^(a[310] & b[200])^(a[309] & b[201])^(a[308] & b[202])^(a[307] & b[203])^(a[306] & b[204])^(a[305] & b[205])^(a[304] & b[206])^(a[303] & b[207])^(a[302] & b[208])^(a[301] & b[209])^(a[300] & b[210])^(a[299] & b[211])^(a[298] & b[212])^(a[297] & b[213])^(a[296] & b[214])^(a[295] & b[215])^(a[294] & b[216])^(a[293] & b[217])^(a[292] & b[218])^(a[291] & b[219])^(a[290] & b[220])^(a[289] & b[221])^(a[288] & b[222])^(a[287] & b[223])^(a[286] & b[224])^(a[285] & b[225])^(a[284] & b[226])^(a[283] & b[227])^(a[282] & b[228])^(a[281] & b[229])^(a[280] & b[230])^(a[279] & b[231])^(a[278] & b[232])^(a[277] & b[233])^(a[276] & b[234])^(a[275] & b[235])^(a[274] & b[236])^(a[273] & b[237])^(a[272] & b[238])^(a[271] & b[239])^(a[270] & b[240])^(a[269] & b[241])^(a[268] & b[242])^(a[267] & b[243])^(a[266] & b[244])^(a[265] & b[245])^(a[264] & b[246])^(a[263] & b[247])^(a[262] & b[248])^(a[261] & b[249])^(a[260] & b[250])^(a[259] & b[251])^(a[258] & b[252])^(a[257] & b[253])^(a[256] & b[254])^(a[255] & b[255])^(a[254] & b[256])^(a[253] & b[257])^(a[252] & b[258])^(a[251] & b[259])^(a[250] & b[260])^(a[249] & b[261])^(a[248] & b[262])^(a[247] & b[263])^(a[246] & b[264])^(a[245] & b[265])^(a[244] & b[266])^(a[243] & b[267])^(a[242] & b[268])^(a[241] & b[269])^(a[240] & b[270])^(a[239] & b[271])^(a[238] & b[272])^(a[237] & b[273])^(a[236] & b[274])^(a[235] & b[275])^(a[234] & b[276])^(a[233] & b[277])^(a[232] & b[278])^(a[231] & b[279])^(a[230] & b[280])^(a[229] & b[281])^(a[228] & b[282])^(a[227] & b[283])^(a[226] & b[284])^(a[225] & b[285])^(a[224] & b[286])^(a[223] & b[287])^(a[222] & b[288])^(a[221] & b[289])^(a[220] & b[290])^(a[219] & b[291])^(a[218] & b[292])^(a[217] & b[293])^(a[216] & b[294])^(a[215] & b[295])^(a[214] & b[296])^(a[213] & b[297])^(a[212] & b[298])^(a[211] & b[299])^(a[210] & b[300])^(a[209] & b[301])^(a[208] & b[302])^(a[207] & b[303])^(a[206] & b[304])^(a[205] & b[305])^(a[204] & b[306])^(a[203] & b[307])^(a[202] & b[308])^(a[201] & b[309])^(a[200] & b[310])^(a[199] & b[311])^(a[198] & b[312])^(a[197] & b[313])^(a[196] & b[314])^(a[195] & b[315])^(a[194] & b[316])^(a[193] & b[317])^(a[192] & b[318])^(a[191] & b[319])^(a[190] & b[320])^(a[189] & b[321])^(a[188] & b[322])^(a[187] & b[323])^(a[186] & b[324])^(a[185] & b[325])^(a[184] & b[326])^(a[183] & b[327])^(a[182] & b[328])^(a[181] & b[329])^(a[180] & b[330])^(a[179] & b[331])^(a[178] & b[332])^(a[177] & b[333])^(a[176] & b[334])^(a[175] & b[335])^(a[174] & b[336])^(a[173] & b[337])^(a[172] & b[338])^(a[171] & b[339])^(a[170] & b[340])^(a[169] & b[341])^(a[168] & b[342])^(a[167] & b[343])^(a[166] & b[344])^(a[165] & b[345])^(a[164] & b[346])^(a[163] & b[347])^(a[162] & b[348])^(a[161] & b[349])^(a[160] & b[350])^(a[159] & b[351])^(a[158] & b[352])^(a[157] & b[353])^(a[156] & b[354])^(a[155] & b[355])^(a[154] & b[356])^(a[153] & b[357])^(a[152] & b[358])^(a[151] & b[359])^(a[150] & b[360])^(a[149] & b[361])^(a[148] & b[362])^(a[147] & b[363])^(a[146] & b[364])^(a[145] & b[365])^(a[144] & b[366])^(a[143] & b[367])^(a[142] & b[368])^(a[141] & b[369])^(a[140] & b[370])^(a[139] & b[371])^(a[138] & b[372])^(a[137] & b[373])^(a[136] & b[374])^(a[135] & b[375])^(a[134] & b[376])^(a[133] & b[377])^(a[132] & b[378])^(a[131] & b[379])^(a[130] & b[380])^(a[129] & b[381])^(a[128] & b[382])^(a[127] & b[383])^(a[126] & b[384])^(a[125] & b[385])^(a[124] & b[386])^(a[123] & b[387])^(a[122] & b[388])^(a[121] & b[389])^(a[120] & b[390])^(a[119] & b[391])^(a[118] & b[392])^(a[117] & b[393])^(a[116] & b[394])^(a[115] & b[395])^(a[114] & b[396])^(a[113] & b[397])^(a[112] & b[398])^(a[111] & b[399])^(a[110] & b[400])^(a[109] & b[401])^(a[108] & b[402])^(a[107] & b[403])^(a[106] & b[404])^(a[105] & b[405])^(a[104] & b[406])^(a[103] & b[407])^(a[102] & b[408]);
assign y[511] = (a[408] & b[103])^(a[407] & b[104])^(a[406] & b[105])^(a[405] & b[106])^(a[404] & b[107])^(a[403] & b[108])^(a[402] & b[109])^(a[401] & b[110])^(a[400] & b[111])^(a[399] & b[112])^(a[398] & b[113])^(a[397] & b[114])^(a[396] & b[115])^(a[395] & b[116])^(a[394] & b[117])^(a[393] & b[118])^(a[392] & b[119])^(a[391] & b[120])^(a[390] & b[121])^(a[389] & b[122])^(a[388] & b[123])^(a[387] & b[124])^(a[386] & b[125])^(a[385] & b[126])^(a[384] & b[127])^(a[383] & b[128])^(a[382] & b[129])^(a[381] & b[130])^(a[380] & b[131])^(a[379] & b[132])^(a[378] & b[133])^(a[377] & b[134])^(a[376] & b[135])^(a[375] & b[136])^(a[374] & b[137])^(a[373] & b[138])^(a[372] & b[139])^(a[371] & b[140])^(a[370] & b[141])^(a[369] & b[142])^(a[368] & b[143])^(a[367] & b[144])^(a[366] & b[145])^(a[365] & b[146])^(a[364] & b[147])^(a[363] & b[148])^(a[362] & b[149])^(a[361] & b[150])^(a[360] & b[151])^(a[359] & b[152])^(a[358] & b[153])^(a[357] & b[154])^(a[356] & b[155])^(a[355] & b[156])^(a[354] & b[157])^(a[353] & b[158])^(a[352] & b[159])^(a[351] & b[160])^(a[350] & b[161])^(a[349] & b[162])^(a[348] & b[163])^(a[347] & b[164])^(a[346] & b[165])^(a[345] & b[166])^(a[344] & b[167])^(a[343] & b[168])^(a[342] & b[169])^(a[341] & b[170])^(a[340] & b[171])^(a[339] & b[172])^(a[338] & b[173])^(a[337] & b[174])^(a[336] & b[175])^(a[335] & b[176])^(a[334] & b[177])^(a[333] & b[178])^(a[332] & b[179])^(a[331] & b[180])^(a[330] & b[181])^(a[329] & b[182])^(a[328] & b[183])^(a[327] & b[184])^(a[326] & b[185])^(a[325] & b[186])^(a[324] & b[187])^(a[323] & b[188])^(a[322] & b[189])^(a[321] & b[190])^(a[320] & b[191])^(a[319] & b[192])^(a[318] & b[193])^(a[317] & b[194])^(a[316] & b[195])^(a[315] & b[196])^(a[314] & b[197])^(a[313] & b[198])^(a[312] & b[199])^(a[311] & b[200])^(a[310] & b[201])^(a[309] & b[202])^(a[308] & b[203])^(a[307] & b[204])^(a[306] & b[205])^(a[305] & b[206])^(a[304] & b[207])^(a[303] & b[208])^(a[302] & b[209])^(a[301] & b[210])^(a[300] & b[211])^(a[299] & b[212])^(a[298] & b[213])^(a[297] & b[214])^(a[296] & b[215])^(a[295] & b[216])^(a[294] & b[217])^(a[293] & b[218])^(a[292] & b[219])^(a[291] & b[220])^(a[290] & b[221])^(a[289] & b[222])^(a[288] & b[223])^(a[287] & b[224])^(a[286] & b[225])^(a[285] & b[226])^(a[284] & b[227])^(a[283] & b[228])^(a[282] & b[229])^(a[281] & b[230])^(a[280] & b[231])^(a[279] & b[232])^(a[278] & b[233])^(a[277] & b[234])^(a[276] & b[235])^(a[275] & b[236])^(a[274] & b[237])^(a[273] & b[238])^(a[272] & b[239])^(a[271] & b[240])^(a[270] & b[241])^(a[269] & b[242])^(a[268] & b[243])^(a[267] & b[244])^(a[266] & b[245])^(a[265] & b[246])^(a[264] & b[247])^(a[263] & b[248])^(a[262] & b[249])^(a[261] & b[250])^(a[260] & b[251])^(a[259] & b[252])^(a[258] & b[253])^(a[257] & b[254])^(a[256] & b[255])^(a[255] & b[256])^(a[254] & b[257])^(a[253] & b[258])^(a[252] & b[259])^(a[251] & b[260])^(a[250] & b[261])^(a[249] & b[262])^(a[248] & b[263])^(a[247] & b[264])^(a[246] & b[265])^(a[245] & b[266])^(a[244] & b[267])^(a[243] & b[268])^(a[242] & b[269])^(a[241] & b[270])^(a[240] & b[271])^(a[239] & b[272])^(a[238] & b[273])^(a[237] & b[274])^(a[236] & b[275])^(a[235] & b[276])^(a[234] & b[277])^(a[233] & b[278])^(a[232] & b[279])^(a[231] & b[280])^(a[230] & b[281])^(a[229] & b[282])^(a[228] & b[283])^(a[227] & b[284])^(a[226] & b[285])^(a[225] & b[286])^(a[224] & b[287])^(a[223] & b[288])^(a[222] & b[289])^(a[221] & b[290])^(a[220] & b[291])^(a[219] & b[292])^(a[218] & b[293])^(a[217] & b[294])^(a[216] & b[295])^(a[215] & b[296])^(a[214] & b[297])^(a[213] & b[298])^(a[212] & b[299])^(a[211] & b[300])^(a[210] & b[301])^(a[209] & b[302])^(a[208] & b[303])^(a[207] & b[304])^(a[206] & b[305])^(a[205] & b[306])^(a[204] & b[307])^(a[203] & b[308])^(a[202] & b[309])^(a[201] & b[310])^(a[200] & b[311])^(a[199] & b[312])^(a[198] & b[313])^(a[197] & b[314])^(a[196] & b[315])^(a[195] & b[316])^(a[194] & b[317])^(a[193] & b[318])^(a[192] & b[319])^(a[191] & b[320])^(a[190] & b[321])^(a[189] & b[322])^(a[188] & b[323])^(a[187] & b[324])^(a[186] & b[325])^(a[185] & b[326])^(a[184] & b[327])^(a[183] & b[328])^(a[182] & b[329])^(a[181] & b[330])^(a[180] & b[331])^(a[179] & b[332])^(a[178] & b[333])^(a[177] & b[334])^(a[176] & b[335])^(a[175] & b[336])^(a[174] & b[337])^(a[173] & b[338])^(a[172] & b[339])^(a[171] & b[340])^(a[170] & b[341])^(a[169] & b[342])^(a[168] & b[343])^(a[167] & b[344])^(a[166] & b[345])^(a[165] & b[346])^(a[164] & b[347])^(a[163] & b[348])^(a[162] & b[349])^(a[161] & b[350])^(a[160] & b[351])^(a[159] & b[352])^(a[158] & b[353])^(a[157] & b[354])^(a[156] & b[355])^(a[155] & b[356])^(a[154] & b[357])^(a[153] & b[358])^(a[152] & b[359])^(a[151] & b[360])^(a[150] & b[361])^(a[149] & b[362])^(a[148] & b[363])^(a[147] & b[364])^(a[146] & b[365])^(a[145] & b[366])^(a[144] & b[367])^(a[143] & b[368])^(a[142] & b[369])^(a[141] & b[370])^(a[140] & b[371])^(a[139] & b[372])^(a[138] & b[373])^(a[137] & b[374])^(a[136] & b[375])^(a[135] & b[376])^(a[134] & b[377])^(a[133] & b[378])^(a[132] & b[379])^(a[131] & b[380])^(a[130] & b[381])^(a[129] & b[382])^(a[128] & b[383])^(a[127] & b[384])^(a[126] & b[385])^(a[125] & b[386])^(a[124] & b[387])^(a[123] & b[388])^(a[122] & b[389])^(a[121] & b[390])^(a[120] & b[391])^(a[119] & b[392])^(a[118] & b[393])^(a[117] & b[394])^(a[116] & b[395])^(a[115] & b[396])^(a[114] & b[397])^(a[113] & b[398])^(a[112] & b[399])^(a[111] & b[400])^(a[110] & b[401])^(a[109] & b[402])^(a[108] & b[403])^(a[107] & b[404])^(a[106] & b[405])^(a[105] & b[406])^(a[104] & b[407])^(a[103] & b[408]);
assign y[512] = (a[408] & b[104])^(a[407] & b[105])^(a[406] & b[106])^(a[405] & b[107])^(a[404] & b[108])^(a[403] & b[109])^(a[402] & b[110])^(a[401] & b[111])^(a[400] & b[112])^(a[399] & b[113])^(a[398] & b[114])^(a[397] & b[115])^(a[396] & b[116])^(a[395] & b[117])^(a[394] & b[118])^(a[393] & b[119])^(a[392] & b[120])^(a[391] & b[121])^(a[390] & b[122])^(a[389] & b[123])^(a[388] & b[124])^(a[387] & b[125])^(a[386] & b[126])^(a[385] & b[127])^(a[384] & b[128])^(a[383] & b[129])^(a[382] & b[130])^(a[381] & b[131])^(a[380] & b[132])^(a[379] & b[133])^(a[378] & b[134])^(a[377] & b[135])^(a[376] & b[136])^(a[375] & b[137])^(a[374] & b[138])^(a[373] & b[139])^(a[372] & b[140])^(a[371] & b[141])^(a[370] & b[142])^(a[369] & b[143])^(a[368] & b[144])^(a[367] & b[145])^(a[366] & b[146])^(a[365] & b[147])^(a[364] & b[148])^(a[363] & b[149])^(a[362] & b[150])^(a[361] & b[151])^(a[360] & b[152])^(a[359] & b[153])^(a[358] & b[154])^(a[357] & b[155])^(a[356] & b[156])^(a[355] & b[157])^(a[354] & b[158])^(a[353] & b[159])^(a[352] & b[160])^(a[351] & b[161])^(a[350] & b[162])^(a[349] & b[163])^(a[348] & b[164])^(a[347] & b[165])^(a[346] & b[166])^(a[345] & b[167])^(a[344] & b[168])^(a[343] & b[169])^(a[342] & b[170])^(a[341] & b[171])^(a[340] & b[172])^(a[339] & b[173])^(a[338] & b[174])^(a[337] & b[175])^(a[336] & b[176])^(a[335] & b[177])^(a[334] & b[178])^(a[333] & b[179])^(a[332] & b[180])^(a[331] & b[181])^(a[330] & b[182])^(a[329] & b[183])^(a[328] & b[184])^(a[327] & b[185])^(a[326] & b[186])^(a[325] & b[187])^(a[324] & b[188])^(a[323] & b[189])^(a[322] & b[190])^(a[321] & b[191])^(a[320] & b[192])^(a[319] & b[193])^(a[318] & b[194])^(a[317] & b[195])^(a[316] & b[196])^(a[315] & b[197])^(a[314] & b[198])^(a[313] & b[199])^(a[312] & b[200])^(a[311] & b[201])^(a[310] & b[202])^(a[309] & b[203])^(a[308] & b[204])^(a[307] & b[205])^(a[306] & b[206])^(a[305] & b[207])^(a[304] & b[208])^(a[303] & b[209])^(a[302] & b[210])^(a[301] & b[211])^(a[300] & b[212])^(a[299] & b[213])^(a[298] & b[214])^(a[297] & b[215])^(a[296] & b[216])^(a[295] & b[217])^(a[294] & b[218])^(a[293] & b[219])^(a[292] & b[220])^(a[291] & b[221])^(a[290] & b[222])^(a[289] & b[223])^(a[288] & b[224])^(a[287] & b[225])^(a[286] & b[226])^(a[285] & b[227])^(a[284] & b[228])^(a[283] & b[229])^(a[282] & b[230])^(a[281] & b[231])^(a[280] & b[232])^(a[279] & b[233])^(a[278] & b[234])^(a[277] & b[235])^(a[276] & b[236])^(a[275] & b[237])^(a[274] & b[238])^(a[273] & b[239])^(a[272] & b[240])^(a[271] & b[241])^(a[270] & b[242])^(a[269] & b[243])^(a[268] & b[244])^(a[267] & b[245])^(a[266] & b[246])^(a[265] & b[247])^(a[264] & b[248])^(a[263] & b[249])^(a[262] & b[250])^(a[261] & b[251])^(a[260] & b[252])^(a[259] & b[253])^(a[258] & b[254])^(a[257] & b[255])^(a[256] & b[256])^(a[255] & b[257])^(a[254] & b[258])^(a[253] & b[259])^(a[252] & b[260])^(a[251] & b[261])^(a[250] & b[262])^(a[249] & b[263])^(a[248] & b[264])^(a[247] & b[265])^(a[246] & b[266])^(a[245] & b[267])^(a[244] & b[268])^(a[243] & b[269])^(a[242] & b[270])^(a[241] & b[271])^(a[240] & b[272])^(a[239] & b[273])^(a[238] & b[274])^(a[237] & b[275])^(a[236] & b[276])^(a[235] & b[277])^(a[234] & b[278])^(a[233] & b[279])^(a[232] & b[280])^(a[231] & b[281])^(a[230] & b[282])^(a[229] & b[283])^(a[228] & b[284])^(a[227] & b[285])^(a[226] & b[286])^(a[225] & b[287])^(a[224] & b[288])^(a[223] & b[289])^(a[222] & b[290])^(a[221] & b[291])^(a[220] & b[292])^(a[219] & b[293])^(a[218] & b[294])^(a[217] & b[295])^(a[216] & b[296])^(a[215] & b[297])^(a[214] & b[298])^(a[213] & b[299])^(a[212] & b[300])^(a[211] & b[301])^(a[210] & b[302])^(a[209] & b[303])^(a[208] & b[304])^(a[207] & b[305])^(a[206] & b[306])^(a[205] & b[307])^(a[204] & b[308])^(a[203] & b[309])^(a[202] & b[310])^(a[201] & b[311])^(a[200] & b[312])^(a[199] & b[313])^(a[198] & b[314])^(a[197] & b[315])^(a[196] & b[316])^(a[195] & b[317])^(a[194] & b[318])^(a[193] & b[319])^(a[192] & b[320])^(a[191] & b[321])^(a[190] & b[322])^(a[189] & b[323])^(a[188] & b[324])^(a[187] & b[325])^(a[186] & b[326])^(a[185] & b[327])^(a[184] & b[328])^(a[183] & b[329])^(a[182] & b[330])^(a[181] & b[331])^(a[180] & b[332])^(a[179] & b[333])^(a[178] & b[334])^(a[177] & b[335])^(a[176] & b[336])^(a[175] & b[337])^(a[174] & b[338])^(a[173] & b[339])^(a[172] & b[340])^(a[171] & b[341])^(a[170] & b[342])^(a[169] & b[343])^(a[168] & b[344])^(a[167] & b[345])^(a[166] & b[346])^(a[165] & b[347])^(a[164] & b[348])^(a[163] & b[349])^(a[162] & b[350])^(a[161] & b[351])^(a[160] & b[352])^(a[159] & b[353])^(a[158] & b[354])^(a[157] & b[355])^(a[156] & b[356])^(a[155] & b[357])^(a[154] & b[358])^(a[153] & b[359])^(a[152] & b[360])^(a[151] & b[361])^(a[150] & b[362])^(a[149] & b[363])^(a[148] & b[364])^(a[147] & b[365])^(a[146] & b[366])^(a[145] & b[367])^(a[144] & b[368])^(a[143] & b[369])^(a[142] & b[370])^(a[141] & b[371])^(a[140] & b[372])^(a[139] & b[373])^(a[138] & b[374])^(a[137] & b[375])^(a[136] & b[376])^(a[135] & b[377])^(a[134] & b[378])^(a[133] & b[379])^(a[132] & b[380])^(a[131] & b[381])^(a[130] & b[382])^(a[129] & b[383])^(a[128] & b[384])^(a[127] & b[385])^(a[126] & b[386])^(a[125] & b[387])^(a[124] & b[388])^(a[123] & b[389])^(a[122] & b[390])^(a[121] & b[391])^(a[120] & b[392])^(a[119] & b[393])^(a[118] & b[394])^(a[117] & b[395])^(a[116] & b[396])^(a[115] & b[397])^(a[114] & b[398])^(a[113] & b[399])^(a[112] & b[400])^(a[111] & b[401])^(a[110] & b[402])^(a[109] & b[403])^(a[108] & b[404])^(a[107] & b[405])^(a[106] & b[406])^(a[105] & b[407])^(a[104] & b[408]);
assign y[513] = (a[408] & b[105])^(a[407] & b[106])^(a[406] & b[107])^(a[405] & b[108])^(a[404] & b[109])^(a[403] & b[110])^(a[402] & b[111])^(a[401] & b[112])^(a[400] & b[113])^(a[399] & b[114])^(a[398] & b[115])^(a[397] & b[116])^(a[396] & b[117])^(a[395] & b[118])^(a[394] & b[119])^(a[393] & b[120])^(a[392] & b[121])^(a[391] & b[122])^(a[390] & b[123])^(a[389] & b[124])^(a[388] & b[125])^(a[387] & b[126])^(a[386] & b[127])^(a[385] & b[128])^(a[384] & b[129])^(a[383] & b[130])^(a[382] & b[131])^(a[381] & b[132])^(a[380] & b[133])^(a[379] & b[134])^(a[378] & b[135])^(a[377] & b[136])^(a[376] & b[137])^(a[375] & b[138])^(a[374] & b[139])^(a[373] & b[140])^(a[372] & b[141])^(a[371] & b[142])^(a[370] & b[143])^(a[369] & b[144])^(a[368] & b[145])^(a[367] & b[146])^(a[366] & b[147])^(a[365] & b[148])^(a[364] & b[149])^(a[363] & b[150])^(a[362] & b[151])^(a[361] & b[152])^(a[360] & b[153])^(a[359] & b[154])^(a[358] & b[155])^(a[357] & b[156])^(a[356] & b[157])^(a[355] & b[158])^(a[354] & b[159])^(a[353] & b[160])^(a[352] & b[161])^(a[351] & b[162])^(a[350] & b[163])^(a[349] & b[164])^(a[348] & b[165])^(a[347] & b[166])^(a[346] & b[167])^(a[345] & b[168])^(a[344] & b[169])^(a[343] & b[170])^(a[342] & b[171])^(a[341] & b[172])^(a[340] & b[173])^(a[339] & b[174])^(a[338] & b[175])^(a[337] & b[176])^(a[336] & b[177])^(a[335] & b[178])^(a[334] & b[179])^(a[333] & b[180])^(a[332] & b[181])^(a[331] & b[182])^(a[330] & b[183])^(a[329] & b[184])^(a[328] & b[185])^(a[327] & b[186])^(a[326] & b[187])^(a[325] & b[188])^(a[324] & b[189])^(a[323] & b[190])^(a[322] & b[191])^(a[321] & b[192])^(a[320] & b[193])^(a[319] & b[194])^(a[318] & b[195])^(a[317] & b[196])^(a[316] & b[197])^(a[315] & b[198])^(a[314] & b[199])^(a[313] & b[200])^(a[312] & b[201])^(a[311] & b[202])^(a[310] & b[203])^(a[309] & b[204])^(a[308] & b[205])^(a[307] & b[206])^(a[306] & b[207])^(a[305] & b[208])^(a[304] & b[209])^(a[303] & b[210])^(a[302] & b[211])^(a[301] & b[212])^(a[300] & b[213])^(a[299] & b[214])^(a[298] & b[215])^(a[297] & b[216])^(a[296] & b[217])^(a[295] & b[218])^(a[294] & b[219])^(a[293] & b[220])^(a[292] & b[221])^(a[291] & b[222])^(a[290] & b[223])^(a[289] & b[224])^(a[288] & b[225])^(a[287] & b[226])^(a[286] & b[227])^(a[285] & b[228])^(a[284] & b[229])^(a[283] & b[230])^(a[282] & b[231])^(a[281] & b[232])^(a[280] & b[233])^(a[279] & b[234])^(a[278] & b[235])^(a[277] & b[236])^(a[276] & b[237])^(a[275] & b[238])^(a[274] & b[239])^(a[273] & b[240])^(a[272] & b[241])^(a[271] & b[242])^(a[270] & b[243])^(a[269] & b[244])^(a[268] & b[245])^(a[267] & b[246])^(a[266] & b[247])^(a[265] & b[248])^(a[264] & b[249])^(a[263] & b[250])^(a[262] & b[251])^(a[261] & b[252])^(a[260] & b[253])^(a[259] & b[254])^(a[258] & b[255])^(a[257] & b[256])^(a[256] & b[257])^(a[255] & b[258])^(a[254] & b[259])^(a[253] & b[260])^(a[252] & b[261])^(a[251] & b[262])^(a[250] & b[263])^(a[249] & b[264])^(a[248] & b[265])^(a[247] & b[266])^(a[246] & b[267])^(a[245] & b[268])^(a[244] & b[269])^(a[243] & b[270])^(a[242] & b[271])^(a[241] & b[272])^(a[240] & b[273])^(a[239] & b[274])^(a[238] & b[275])^(a[237] & b[276])^(a[236] & b[277])^(a[235] & b[278])^(a[234] & b[279])^(a[233] & b[280])^(a[232] & b[281])^(a[231] & b[282])^(a[230] & b[283])^(a[229] & b[284])^(a[228] & b[285])^(a[227] & b[286])^(a[226] & b[287])^(a[225] & b[288])^(a[224] & b[289])^(a[223] & b[290])^(a[222] & b[291])^(a[221] & b[292])^(a[220] & b[293])^(a[219] & b[294])^(a[218] & b[295])^(a[217] & b[296])^(a[216] & b[297])^(a[215] & b[298])^(a[214] & b[299])^(a[213] & b[300])^(a[212] & b[301])^(a[211] & b[302])^(a[210] & b[303])^(a[209] & b[304])^(a[208] & b[305])^(a[207] & b[306])^(a[206] & b[307])^(a[205] & b[308])^(a[204] & b[309])^(a[203] & b[310])^(a[202] & b[311])^(a[201] & b[312])^(a[200] & b[313])^(a[199] & b[314])^(a[198] & b[315])^(a[197] & b[316])^(a[196] & b[317])^(a[195] & b[318])^(a[194] & b[319])^(a[193] & b[320])^(a[192] & b[321])^(a[191] & b[322])^(a[190] & b[323])^(a[189] & b[324])^(a[188] & b[325])^(a[187] & b[326])^(a[186] & b[327])^(a[185] & b[328])^(a[184] & b[329])^(a[183] & b[330])^(a[182] & b[331])^(a[181] & b[332])^(a[180] & b[333])^(a[179] & b[334])^(a[178] & b[335])^(a[177] & b[336])^(a[176] & b[337])^(a[175] & b[338])^(a[174] & b[339])^(a[173] & b[340])^(a[172] & b[341])^(a[171] & b[342])^(a[170] & b[343])^(a[169] & b[344])^(a[168] & b[345])^(a[167] & b[346])^(a[166] & b[347])^(a[165] & b[348])^(a[164] & b[349])^(a[163] & b[350])^(a[162] & b[351])^(a[161] & b[352])^(a[160] & b[353])^(a[159] & b[354])^(a[158] & b[355])^(a[157] & b[356])^(a[156] & b[357])^(a[155] & b[358])^(a[154] & b[359])^(a[153] & b[360])^(a[152] & b[361])^(a[151] & b[362])^(a[150] & b[363])^(a[149] & b[364])^(a[148] & b[365])^(a[147] & b[366])^(a[146] & b[367])^(a[145] & b[368])^(a[144] & b[369])^(a[143] & b[370])^(a[142] & b[371])^(a[141] & b[372])^(a[140] & b[373])^(a[139] & b[374])^(a[138] & b[375])^(a[137] & b[376])^(a[136] & b[377])^(a[135] & b[378])^(a[134] & b[379])^(a[133] & b[380])^(a[132] & b[381])^(a[131] & b[382])^(a[130] & b[383])^(a[129] & b[384])^(a[128] & b[385])^(a[127] & b[386])^(a[126] & b[387])^(a[125] & b[388])^(a[124] & b[389])^(a[123] & b[390])^(a[122] & b[391])^(a[121] & b[392])^(a[120] & b[393])^(a[119] & b[394])^(a[118] & b[395])^(a[117] & b[396])^(a[116] & b[397])^(a[115] & b[398])^(a[114] & b[399])^(a[113] & b[400])^(a[112] & b[401])^(a[111] & b[402])^(a[110] & b[403])^(a[109] & b[404])^(a[108] & b[405])^(a[107] & b[406])^(a[106] & b[407])^(a[105] & b[408]);
assign y[514] = (a[408] & b[106])^(a[407] & b[107])^(a[406] & b[108])^(a[405] & b[109])^(a[404] & b[110])^(a[403] & b[111])^(a[402] & b[112])^(a[401] & b[113])^(a[400] & b[114])^(a[399] & b[115])^(a[398] & b[116])^(a[397] & b[117])^(a[396] & b[118])^(a[395] & b[119])^(a[394] & b[120])^(a[393] & b[121])^(a[392] & b[122])^(a[391] & b[123])^(a[390] & b[124])^(a[389] & b[125])^(a[388] & b[126])^(a[387] & b[127])^(a[386] & b[128])^(a[385] & b[129])^(a[384] & b[130])^(a[383] & b[131])^(a[382] & b[132])^(a[381] & b[133])^(a[380] & b[134])^(a[379] & b[135])^(a[378] & b[136])^(a[377] & b[137])^(a[376] & b[138])^(a[375] & b[139])^(a[374] & b[140])^(a[373] & b[141])^(a[372] & b[142])^(a[371] & b[143])^(a[370] & b[144])^(a[369] & b[145])^(a[368] & b[146])^(a[367] & b[147])^(a[366] & b[148])^(a[365] & b[149])^(a[364] & b[150])^(a[363] & b[151])^(a[362] & b[152])^(a[361] & b[153])^(a[360] & b[154])^(a[359] & b[155])^(a[358] & b[156])^(a[357] & b[157])^(a[356] & b[158])^(a[355] & b[159])^(a[354] & b[160])^(a[353] & b[161])^(a[352] & b[162])^(a[351] & b[163])^(a[350] & b[164])^(a[349] & b[165])^(a[348] & b[166])^(a[347] & b[167])^(a[346] & b[168])^(a[345] & b[169])^(a[344] & b[170])^(a[343] & b[171])^(a[342] & b[172])^(a[341] & b[173])^(a[340] & b[174])^(a[339] & b[175])^(a[338] & b[176])^(a[337] & b[177])^(a[336] & b[178])^(a[335] & b[179])^(a[334] & b[180])^(a[333] & b[181])^(a[332] & b[182])^(a[331] & b[183])^(a[330] & b[184])^(a[329] & b[185])^(a[328] & b[186])^(a[327] & b[187])^(a[326] & b[188])^(a[325] & b[189])^(a[324] & b[190])^(a[323] & b[191])^(a[322] & b[192])^(a[321] & b[193])^(a[320] & b[194])^(a[319] & b[195])^(a[318] & b[196])^(a[317] & b[197])^(a[316] & b[198])^(a[315] & b[199])^(a[314] & b[200])^(a[313] & b[201])^(a[312] & b[202])^(a[311] & b[203])^(a[310] & b[204])^(a[309] & b[205])^(a[308] & b[206])^(a[307] & b[207])^(a[306] & b[208])^(a[305] & b[209])^(a[304] & b[210])^(a[303] & b[211])^(a[302] & b[212])^(a[301] & b[213])^(a[300] & b[214])^(a[299] & b[215])^(a[298] & b[216])^(a[297] & b[217])^(a[296] & b[218])^(a[295] & b[219])^(a[294] & b[220])^(a[293] & b[221])^(a[292] & b[222])^(a[291] & b[223])^(a[290] & b[224])^(a[289] & b[225])^(a[288] & b[226])^(a[287] & b[227])^(a[286] & b[228])^(a[285] & b[229])^(a[284] & b[230])^(a[283] & b[231])^(a[282] & b[232])^(a[281] & b[233])^(a[280] & b[234])^(a[279] & b[235])^(a[278] & b[236])^(a[277] & b[237])^(a[276] & b[238])^(a[275] & b[239])^(a[274] & b[240])^(a[273] & b[241])^(a[272] & b[242])^(a[271] & b[243])^(a[270] & b[244])^(a[269] & b[245])^(a[268] & b[246])^(a[267] & b[247])^(a[266] & b[248])^(a[265] & b[249])^(a[264] & b[250])^(a[263] & b[251])^(a[262] & b[252])^(a[261] & b[253])^(a[260] & b[254])^(a[259] & b[255])^(a[258] & b[256])^(a[257] & b[257])^(a[256] & b[258])^(a[255] & b[259])^(a[254] & b[260])^(a[253] & b[261])^(a[252] & b[262])^(a[251] & b[263])^(a[250] & b[264])^(a[249] & b[265])^(a[248] & b[266])^(a[247] & b[267])^(a[246] & b[268])^(a[245] & b[269])^(a[244] & b[270])^(a[243] & b[271])^(a[242] & b[272])^(a[241] & b[273])^(a[240] & b[274])^(a[239] & b[275])^(a[238] & b[276])^(a[237] & b[277])^(a[236] & b[278])^(a[235] & b[279])^(a[234] & b[280])^(a[233] & b[281])^(a[232] & b[282])^(a[231] & b[283])^(a[230] & b[284])^(a[229] & b[285])^(a[228] & b[286])^(a[227] & b[287])^(a[226] & b[288])^(a[225] & b[289])^(a[224] & b[290])^(a[223] & b[291])^(a[222] & b[292])^(a[221] & b[293])^(a[220] & b[294])^(a[219] & b[295])^(a[218] & b[296])^(a[217] & b[297])^(a[216] & b[298])^(a[215] & b[299])^(a[214] & b[300])^(a[213] & b[301])^(a[212] & b[302])^(a[211] & b[303])^(a[210] & b[304])^(a[209] & b[305])^(a[208] & b[306])^(a[207] & b[307])^(a[206] & b[308])^(a[205] & b[309])^(a[204] & b[310])^(a[203] & b[311])^(a[202] & b[312])^(a[201] & b[313])^(a[200] & b[314])^(a[199] & b[315])^(a[198] & b[316])^(a[197] & b[317])^(a[196] & b[318])^(a[195] & b[319])^(a[194] & b[320])^(a[193] & b[321])^(a[192] & b[322])^(a[191] & b[323])^(a[190] & b[324])^(a[189] & b[325])^(a[188] & b[326])^(a[187] & b[327])^(a[186] & b[328])^(a[185] & b[329])^(a[184] & b[330])^(a[183] & b[331])^(a[182] & b[332])^(a[181] & b[333])^(a[180] & b[334])^(a[179] & b[335])^(a[178] & b[336])^(a[177] & b[337])^(a[176] & b[338])^(a[175] & b[339])^(a[174] & b[340])^(a[173] & b[341])^(a[172] & b[342])^(a[171] & b[343])^(a[170] & b[344])^(a[169] & b[345])^(a[168] & b[346])^(a[167] & b[347])^(a[166] & b[348])^(a[165] & b[349])^(a[164] & b[350])^(a[163] & b[351])^(a[162] & b[352])^(a[161] & b[353])^(a[160] & b[354])^(a[159] & b[355])^(a[158] & b[356])^(a[157] & b[357])^(a[156] & b[358])^(a[155] & b[359])^(a[154] & b[360])^(a[153] & b[361])^(a[152] & b[362])^(a[151] & b[363])^(a[150] & b[364])^(a[149] & b[365])^(a[148] & b[366])^(a[147] & b[367])^(a[146] & b[368])^(a[145] & b[369])^(a[144] & b[370])^(a[143] & b[371])^(a[142] & b[372])^(a[141] & b[373])^(a[140] & b[374])^(a[139] & b[375])^(a[138] & b[376])^(a[137] & b[377])^(a[136] & b[378])^(a[135] & b[379])^(a[134] & b[380])^(a[133] & b[381])^(a[132] & b[382])^(a[131] & b[383])^(a[130] & b[384])^(a[129] & b[385])^(a[128] & b[386])^(a[127] & b[387])^(a[126] & b[388])^(a[125] & b[389])^(a[124] & b[390])^(a[123] & b[391])^(a[122] & b[392])^(a[121] & b[393])^(a[120] & b[394])^(a[119] & b[395])^(a[118] & b[396])^(a[117] & b[397])^(a[116] & b[398])^(a[115] & b[399])^(a[114] & b[400])^(a[113] & b[401])^(a[112] & b[402])^(a[111] & b[403])^(a[110] & b[404])^(a[109] & b[405])^(a[108] & b[406])^(a[107] & b[407])^(a[106] & b[408]);
assign y[515] = (a[408] & b[107])^(a[407] & b[108])^(a[406] & b[109])^(a[405] & b[110])^(a[404] & b[111])^(a[403] & b[112])^(a[402] & b[113])^(a[401] & b[114])^(a[400] & b[115])^(a[399] & b[116])^(a[398] & b[117])^(a[397] & b[118])^(a[396] & b[119])^(a[395] & b[120])^(a[394] & b[121])^(a[393] & b[122])^(a[392] & b[123])^(a[391] & b[124])^(a[390] & b[125])^(a[389] & b[126])^(a[388] & b[127])^(a[387] & b[128])^(a[386] & b[129])^(a[385] & b[130])^(a[384] & b[131])^(a[383] & b[132])^(a[382] & b[133])^(a[381] & b[134])^(a[380] & b[135])^(a[379] & b[136])^(a[378] & b[137])^(a[377] & b[138])^(a[376] & b[139])^(a[375] & b[140])^(a[374] & b[141])^(a[373] & b[142])^(a[372] & b[143])^(a[371] & b[144])^(a[370] & b[145])^(a[369] & b[146])^(a[368] & b[147])^(a[367] & b[148])^(a[366] & b[149])^(a[365] & b[150])^(a[364] & b[151])^(a[363] & b[152])^(a[362] & b[153])^(a[361] & b[154])^(a[360] & b[155])^(a[359] & b[156])^(a[358] & b[157])^(a[357] & b[158])^(a[356] & b[159])^(a[355] & b[160])^(a[354] & b[161])^(a[353] & b[162])^(a[352] & b[163])^(a[351] & b[164])^(a[350] & b[165])^(a[349] & b[166])^(a[348] & b[167])^(a[347] & b[168])^(a[346] & b[169])^(a[345] & b[170])^(a[344] & b[171])^(a[343] & b[172])^(a[342] & b[173])^(a[341] & b[174])^(a[340] & b[175])^(a[339] & b[176])^(a[338] & b[177])^(a[337] & b[178])^(a[336] & b[179])^(a[335] & b[180])^(a[334] & b[181])^(a[333] & b[182])^(a[332] & b[183])^(a[331] & b[184])^(a[330] & b[185])^(a[329] & b[186])^(a[328] & b[187])^(a[327] & b[188])^(a[326] & b[189])^(a[325] & b[190])^(a[324] & b[191])^(a[323] & b[192])^(a[322] & b[193])^(a[321] & b[194])^(a[320] & b[195])^(a[319] & b[196])^(a[318] & b[197])^(a[317] & b[198])^(a[316] & b[199])^(a[315] & b[200])^(a[314] & b[201])^(a[313] & b[202])^(a[312] & b[203])^(a[311] & b[204])^(a[310] & b[205])^(a[309] & b[206])^(a[308] & b[207])^(a[307] & b[208])^(a[306] & b[209])^(a[305] & b[210])^(a[304] & b[211])^(a[303] & b[212])^(a[302] & b[213])^(a[301] & b[214])^(a[300] & b[215])^(a[299] & b[216])^(a[298] & b[217])^(a[297] & b[218])^(a[296] & b[219])^(a[295] & b[220])^(a[294] & b[221])^(a[293] & b[222])^(a[292] & b[223])^(a[291] & b[224])^(a[290] & b[225])^(a[289] & b[226])^(a[288] & b[227])^(a[287] & b[228])^(a[286] & b[229])^(a[285] & b[230])^(a[284] & b[231])^(a[283] & b[232])^(a[282] & b[233])^(a[281] & b[234])^(a[280] & b[235])^(a[279] & b[236])^(a[278] & b[237])^(a[277] & b[238])^(a[276] & b[239])^(a[275] & b[240])^(a[274] & b[241])^(a[273] & b[242])^(a[272] & b[243])^(a[271] & b[244])^(a[270] & b[245])^(a[269] & b[246])^(a[268] & b[247])^(a[267] & b[248])^(a[266] & b[249])^(a[265] & b[250])^(a[264] & b[251])^(a[263] & b[252])^(a[262] & b[253])^(a[261] & b[254])^(a[260] & b[255])^(a[259] & b[256])^(a[258] & b[257])^(a[257] & b[258])^(a[256] & b[259])^(a[255] & b[260])^(a[254] & b[261])^(a[253] & b[262])^(a[252] & b[263])^(a[251] & b[264])^(a[250] & b[265])^(a[249] & b[266])^(a[248] & b[267])^(a[247] & b[268])^(a[246] & b[269])^(a[245] & b[270])^(a[244] & b[271])^(a[243] & b[272])^(a[242] & b[273])^(a[241] & b[274])^(a[240] & b[275])^(a[239] & b[276])^(a[238] & b[277])^(a[237] & b[278])^(a[236] & b[279])^(a[235] & b[280])^(a[234] & b[281])^(a[233] & b[282])^(a[232] & b[283])^(a[231] & b[284])^(a[230] & b[285])^(a[229] & b[286])^(a[228] & b[287])^(a[227] & b[288])^(a[226] & b[289])^(a[225] & b[290])^(a[224] & b[291])^(a[223] & b[292])^(a[222] & b[293])^(a[221] & b[294])^(a[220] & b[295])^(a[219] & b[296])^(a[218] & b[297])^(a[217] & b[298])^(a[216] & b[299])^(a[215] & b[300])^(a[214] & b[301])^(a[213] & b[302])^(a[212] & b[303])^(a[211] & b[304])^(a[210] & b[305])^(a[209] & b[306])^(a[208] & b[307])^(a[207] & b[308])^(a[206] & b[309])^(a[205] & b[310])^(a[204] & b[311])^(a[203] & b[312])^(a[202] & b[313])^(a[201] & b[314])^(a[200] & b[315])^(a[199] & b[316])^(a[198] & b[317])^(a[197] & b[318])^(a[196] & b[319])^(a[195] & b[320])^(a[194] & b[321])^(a[193] & b[322])^(a[192] & b[323])^(a[191] & b[324])^(a[190] & b[325])^(a[189] & b[326])^(a[188] & b[327])^(a[187] & b[328])^(a[186] & b[329])^(a[185] & b[330])^(a[184] & b[331])^(a[183] & b[332])^(a[182] & b[333])^(a[181] & b[334])^(a[180] & b[335])^(a[179] & b[336])^(a[178] & b[337])^(a[177] & b[338])^(a[176] & b[339])^(a[175] & b[340])^(a[174] & b[341])^(a[173] & b[342])^(a[172] & b[343])^(a[171] & b[344])^(a[170] & b[345])^(a[169] & b[346])^(a[168] & b[347])^(a[167] & b[348])^(a[166] & b[349])^(a[165] & b[350])^(a[164] & b[351])^(a[163] & b[352])^(a[162] & b[353])^(a[161] & b[354])^(a[160] & b[355])^(a[159] & b[356])^(a[158] & b[357])^(a[157] & b[358])^(a[156] & b[359])^(a[155] & b[360])^(a[154] & b[361])^(a[153] & b[362])^(a[152] & b[363])^(a[151] & b[364])^(a[150] & b[365])^(a[149] & b[366])^(a[148] & b[367])^(a[147] & b[368])^(a[146] & b[369])^(a[145] & b[370])^(a[144] & b[371])^(a[143] & b[372])^(a[142] & b[373])^(a[141] & b[374])^(a[140] & b[375])^(a[139] & b[376])^(a[138] & b[377])^(a[137] & b[378])^(a[136] & b[379])^(a[135] & b[380])^(a[134] & b[381])^(a[133] & b[382])^(a[132] & b[383])^(a[131] & b[384])^(a[130] & b[385])^(a[129] & b[386])^(a[128] & b[387])^(a[127] & b[388])^(a[126] & b[389])^(a[125] & b[390])^(a[124] & b[391])^(a[123] & b[392])^(a[122] & b[393])^(a[121] & b[394])^(a[120] & b[395])^(a[119] & b[396])^(a[118] & b[397])^(a[117] & b[398])^(a[116] & b[399])^(a[115] & b[400])^(a[114] & b[401])^(a[113] & b[402])^(a[112] & b[403])^(a[111] & b[404])^(a[110] & b[405])^(a[109] & b[406])^(a[108] & b[407])^(a[107] & b[408]);
assign y[516] = (a[408] & b[108])^(a[407] & b[109])^(a[406] & b[110])^(a[405] & b[111])^(a[404] & b[112])^(a[403] & b[113])^(a[402] & b[114])^(a[401] & b[115])^(a[400] & b[116])^(a[399] & b[117])^(a[398] & b[118])^(a[397] & b[119])^(a[396] & b[120])^(a[395] & b[121])^(a[394] & b[122])^(a[393] & b[123])^(a[392] & b[124])^(a[391] & b[125])^(a[390] & b[126])^(a[389] & b[127])^(a[388] & b[128])^(a[387] & b[129])^(a[386] & b[130])^(a[385] & b[131])^(a[384] & b[132])^(a[383] & b[133])^(a[382] & b[134])^(a[381] & b[135])^(a[380] & b[136])^(a[379] & b[137])^(a[378] & b[138])^(a[377] & b[139])^(a[376] & b[140])^(a[375] & b[141])^(a[374] & b[142])^(a[373] & b[143])^(a[372] & b[144])^(a[371] & b[145])^(a[370] & b[146])^(a[369] & b[147])^(a[368] & b[148])^(a[367] & b[149])^(a[366] & b[150])^(a[365] & b[151])^(a[364] & b[152])^(a[363] & b[153])^(a[362] & b[154])^(a[361] & b[155])^(a[360] & b[156])^(a[359] & b[157])^(a[358] & b[158])^(a[357] & b[159])^(a[356] & b[160])^(a[355] & b[161])^(a[354] & b[162])^(a[353] & b[163])^(a[352] & b[164])^(a[351] & b[165])^(a[350] & b[166])^(a[349] & b[167])^(a[348] & b[168])^(a[347] & b[169])^(a[346] & b[170])^(a[345] & b[171])^(a[344] & b[172])^(a[343] & b[173])^(a[342] & b[174])^(a[341] & b[175])^(a[340] & b[176])^(a[339] & b[177])^(a[338] & b[178])^(a[337] & b[179])^(a[336] & b[180])^(a[335] & b[181])^(a[334] & b[182])^(a[333] & b[183])^(a[332] & b[184])^(a[331] & b[185])^(a[330] & b[186])^(a[329] & b[187])^(a[328] & b[188])^(a[327] & b[189])^(a[326] & b[190])^(a[325] & b[191])^(a[324] & b[192])^(a[323] & b[193])^(a[322] & b[194])^(a[321] & b[195])^(a[320] & b[196])^(a[319] & b[197])^(a[318] & b[198])^(a[317] & b[199])^(a[316] & b[200])^(a[315] & b[201])^(a[314] & b[202])^(a[313] & b[203])^(a[312] & b[204])^(a[311] & b[205])^(a[310] & b[206])^(a[309] & b[207])^(a[308] & b[208])^(a[307] & b[209])^(a[306] & b[210])^(a[305] & b[211])^(a[304] & b[212])^(a[303] & b[213])^(a[302] & b[214])^(a[301] & b[215])^(a[300] & b[216])^(a[299] & b[217])^(a[298] & b[218])^(a[297] & b[219])^(a[296] & b[220])^(a[295] & b[221])^(a[294] & b[222])^(a[293] & b[223])^(a[292] & b[224])^(a[291] & b[225])^(a[290] & b[226])^(a[289] & b[227])^(a[288] & b[228])^(a[287] & b[229])^(a[286] & b[230])^(a[285] & b[231])^(a[284] & b[232])^(a[283] & b[233])^(a[282] & b[234])^(a[281] & b[235])^(a[280] & b[236])^(a[279] & b[237])^(a[278] & b[238])^(a[277] & b[239])^(a[276] & b[240])^(a[275] & b[241])^(a[274] & b[242])^(a[273] & b[243])^(a[272] & b[244])^(a[271] & b[245])^(a[270] & b[246])^(a[269] & b[247])^(a[268] & b[248])^(a[267] & b[249])^(a[266] & b[250])^(a[265] & b[251])^(a[264] & b[252])^(a[263] & b[253])^(a[262] & b[254])^(a[261] & b[255])^(a[260] & b[256])^(a[259] & b[257])^(a[258] & b[258])^(a[257] & b[259])^(a[256] & b[260])^(a[255] & b[261])^(a[254] & b[262])^(a[253] & b[263])^(a[252] & b[264])^(a[251] & b[265])^(a[250] & b[266])^(a[249] & b[267])^(a[248] & b[268])^(a[247] & b[269])^(a[246] & b[270])^(a[245] & b[271])^(a[244] & b[272])^(a[243] & b[273])^(a[242] & b[274])^(a[241] & b[275])^(a[240] & b[276])^(a[239] & b[277])^(a[238] & b[278])^(a[237] & b[279])^(a[236] & b[280])^(a[235] & b[281])^(a[234] & b[282])^(a[233] & b[283])^(a[232] & b[284])^(a[231] & b[285])^(a[230] & b[286])^(a[229] & b[287])^(a[228] & b[288])^(a[227] & b[289])^(a[226] & b[290])^(a[225] & b[291])^(a[224] & b[292])^(a[223] & b[293])^(a[222] & b[294])^(a[221] & b[295])^(a[220] & b[296])^(a[219] & b[297])^(a[218] & b[298])^(a[217] & b[299])^(a[216] & b[300])^(a[215] & b[301])^(a[214] & b[302])^(a[213] & b[303])^(a[212] & b[304])^(a[211] & b[305])^(a[210] & b[306])^(a[209] & b[307])^(a[208] & b[308])^(a[207] & b[309])^(a[206] & b[310])^(a[205] & b[311])^(a[204] & b[312])^(a[203] & b[313])^(a[202] & b[314])^(a[201] & b[315])^(a[200] & b[316])^(a[199] & b[317])^(a[198] & b[318])^(a[197] & b[319])^(a[196] & b[320])^(a[195] & b[321])^(a[194] & b[322])^(a[193] & b[323])^(a[192] & b[324])^(a[191] & b[325])^(a[190] & b[326])^(a[189] & b[327])^(a[188] & b[328])^(a[187] & b[329])^(a[186] & b[330])^(a[185] & b[331])^(a[184] & b[332])^(a[183] & b[333])^(a[182] & b[334])^(a[181] & b[335])^(a[180] & b[336])^(a[179] & b[337])^(a[178] & b[338])^(a[177] & b[339])^(a[176] & b[340])^(a[175] & b[341])^(a[174] & b[342])^(a[173] & b[343])^(a[172] & b[344])^(a[171] & b[345])^(a[170] & b[346])^(a[169] & b[347])^(a[168] & b[348])^(a[167] & b[349])^(a[166] & b[350])^(a[165] & b[351])^(a[164] & b[352])^(a[163] & b[353])^(a[162] & b[354])^(a[161] & b[355])^(a[160] & b[356])^(a[159] & b[357])^(a[158] & b[358])^(a[157] & b[359])^(a[156] & b[360])^(a[155] & b[361])^(a[154] & b[362])^(a[153] & b[363])^(a[152] & b[364])^(a[151] & b[365])^(a[150] & b[366])^(a[149] & b[367])^(a[148] & b[368])^(a[147] & b[369])^(a[146] & b[370])^(a[145] & b[371])^(a[144] & b[372])^(a[143] & b[373])^(a[142] & b[374])^(a[141] & b[375])^(a[140] & b[376])^(a[139] & b[377])^(a[138] & b[378])^(a[137] & b[379])^(a[136] & b[380])^(a[135] & b[381])^(a[134] & b[382])^(a[133] & b[383])^(a[132] & b[384])^(a[131] & b[385])^(a[130] & b[386])^(a[129] & b[387])^(a[128] & b[388])^(a[127] & b[389])^(a[126] & b[390])^(a[125] & b[391])^(a[124] & b[392])^(a[123] & b[393])^(a[122] & b[394])^(a[121] & b[395])^(a[120] & b[396])^(a[119] & b[397])^(a[118] & b[398])^(a[117] & b[399])^(a[116] & b[400])^(a[115] & b[401])^(a[114] & b[402])^(a[113] & b[403])^(a[112] & b[404])^(a[111] & b[405])^(a[110] & b[406])^(a[109] & b[407])^(a[108] & b[408]);
assign y[517] = (a[408] & b[109])^(a[407] & b[110])^(a[406] & b[111])^(a[405] & b[112])^(a[404] & b[113])^(a[403] & b[114])^(a[402] & b[115])^(a[401] & b[116])^(a[400] & b[117])^(a[399] & b[118])^(a[398] & b[119])^(a[397] & b[120])^(a[396] & b[121])^(a[395] & b[122])^(a[394] & b[123])^(a[393] & b[124])^(a[392] & b[125])^(a[391] & b[126])^(a[390] & b[127])^(a[389] & b[128])^(a[388] & b[129])^(a[387] & b[130])^(a[386] & b[131])^(a[385] & b[132])^(a[384] & b[133])^(a[383] & b[134])^(a[382] & b[135])^(a[381] & b[136])^(a[380] & b[137])^(a[379] & b[138])^(a[378] & b[139])^(a[377] & b[140])^(a[376] & b[141])^(a[375] & b[142])^(a[374] & b[143])^(a[373] & b[144])^(a[372] & b[145])^(a[371] & b[146])^(a[370] & b[147])^(a[369] & b[148])^(a[368] & b[149])^(a[367] & b[150])^(a[366] & b[151])^(a[365] & b[152])^(a[364] & b[153])^(a[363] & b[154])^(a[362] & b[155])^(a[361] & b[156])^(a[360] & b[157])^(a[359] & b[158])^(a[358] & b[159])^(a[357] & b[160])^(a[356] & b[161])^(a[355] & b[162])^(a[354] & b[163])^(a[353] & b[164])^(a[352] & b[165])^(a[351] & b[166])^(a[350] & b[167])^(a[349] & b[168])^(a[348] & b[169])^(a[347] & b[170])^(a[346] & b[171])^(a[345] & b[172])^(a[344] & b[173])^(a[343] & b[174])^(a[342] & b[175])^(a[341] & b[176])^(a[340] & b[177])^(a[339] & b[178])^(a[338] & b[179])^(a[337] & b[180])^(a[336] & b[181])^(a[335] & b[182])^(a[334] & b[183])^(a[333] & b[184])^(a[332] & b[185])^(a[331] & b[186])^(a[330] & b[187])^(a[329] & b[188])^(a[328] & b[189])^(a[327] & b[190])^(a[326] & b[191])^(a[325] & b[192])^(a[324] & b[193])^(a[323] & b[194])^(a[322] & b[195])^(a[321] & b[196])^(a[320] & b[197])^(a[319] & b[198])^(a[318] & b[199])^(a[317] & b[200])^(a[316] & b[201])^(a[315] & b[202])^(a[314] & b[203])^(a[313] & b[204])^(a[312] & b[205])^(a[311] & b[206])^(a[310] & b[207])^(a[309] & b[208])^(a[308] & b[209])^(a[307] & b[210])^(a[306] & b[211])^(a[305] & b[212])^(a[304] & b[213])^(a[303] & b[214])^(a[302] & b[215])^(a[301] & b[216])^(a[300] & b[217])^(a[299] & b[218])^(a[298] & b[219])^(a[297] & b[220])^(a[296] & b[221])^(a[295] & b[222])^(a[294] & b[223])^(a[293] & b[224])^(a[292] & b[225])^(a[291] & b[226])^(a[290] & b[227])^(a[289] & b[228])^(a[288] & b[229])^(a[287] & b[230])^(a[286] & b[231])^(a[285] & b[232])^(a[284] & b[233])^(a[283] & b[234])^(a[282] & b[235])^(a[281] & b[236])^(a[280] & b[237])^(a[279] & b[238])^(a[278] & b[239])^(a[277] & b[240])^(a[276] & b[241])^(a[275] & b[242])^(a[274] & b[243])^(a[273] & b[244])^(a[272] & b[245])^(a[271] & b[246])^(a[270] & b[247])^(a[269] & b[248])^(a[268] & b[249])^(a[267] & b[250])^(a[266] & b[251])^(a[265] & b[252])^(a[264] & b[253])^(a[263] & b[254])^(a[262] & b[255])^(a[261] & b[256])^(a[260] & b[257])^(a[259] & b[258])^(a[258] & b[259])^(a[257] & b[260])^(a[256] & b[261])^(a[255] & b[262])^(a[254] & b[263])^(a[253] & b[264])^(a[252] & b[265])^(a[251] & b[266])^(a[250] & b[267])^(a[249] & b[268])^(a[248] & b[269])^(a[247] & b[270])^(a[246] & b[271])^(a[245] & b[272])^(a[244] & b[273])^(a[243] & b[274])^(a[242] & b[275])^(a[241] & b[276])^(a[240] & b[277])^(a[239] & b[278])^(a[238] & b[279])^(a[237] & b[280])^(a[236] & b[281])^(a[235] & b[282])^(a[234] & b[283])^(a[233] & b[284])^(a[232] & b[285])^(a[231] & b[286])^(a[230] & b[287])^(a[229] & b[288])^(a[228] & b[289])^(a[227] & b[290])^(a[226] & b[291])^(a[225] & b[292])^(a[224] & b[293])^(a[223] & b[294])^(a[222] & b[295])^(a[221] & b[296])^(a[220] & b[297])^(a[219] & b[298])^(a[218] & b[299])^(a[217] & b[300])^(a[216] & b[301])^(a[215] & b[302])^(a[214] & b[303])^(a[213] & b[304])^(a[212] & b[305])^(a[211] & b[306])^(a[210] & b[307])^(a[209] & b[308])^(a[208] & b[309])^(a[207] & b[310])^(a[206] & b[311])^(a[205] & b[312])^(a[204] & b[313])^(a[203] & b[314])^(a[202] & b[315])^(a[201] & b[316])^(a[200] & b[317])^(a[199] & b[318])^(a[198] & b[319])^(a[197] & b[320])^(a[196] & b[321])^(a[195] & b[322])^(a[194] & b[323])^(a[193] & b[324])^(a[192] & b[325])^(a[191] & b[326])^(a[190] & b[327])^(a[189] & b[328])^(a[188] & b[329])^(a[187] & b[330])^(a[186] & b[331])^(a[185] & b[332])^(a[184] & b[333])^(a[183] & b[334])^(a[182] & b[335])^(a[181] & b[336])^(a[180] & b[337])^(a[179] & b[338])^(a[178] & b[339])^(a[177] & b[340])^(a[176] & b[341])^(a[175] & b[342])^(a[174] & b[343])^(a[173] & b[344])^(a[172] & b[345])^(a[171] & b[346])^(a[170] & b[347])^(a[169] & b[348])^(a[168] & b[349])^(a[167] & b[350])^(a[166] & b[351])^(a[165] & b[352])^(a[164] & b[353])^(a[163] & b[354])^(a[162] & b[355])^(a[161] & b[356])^(a[160] & b[357])^(a[159] & b[358])^(a[158] & b[359])^(a[157] & b[360])^(a[156] & b[361])^(a[155] & b[362])^(a[154] & b[363])^(a[153] & b[364])^(a[152] & b[365])^(a[151] & b[366])^(a[150] & b[367])^(a[149] & b[368])^(a[148] & b[369])^(a[147] & b[370])^(a[146] & b[371])^(a[145] & b[372])^(a[144] & b[373])^(a[143] & b[374])^(a[142] & b[375])^(a[141] & b[376])^(a[140] & b[377])^(a[139] & b[378])^(a[138] & b[379])^(a[137] & b[380])^(a[136] & b[381])^(a[135] & b[382])^(a[134] & b[383])^(a[133] & b[384])^(a[132] & b[385])^(a[131] & b[386])^(a[130] & b[387])^(a[129] & b[388])^(a[128] & b[389])^(a[127] & b[390])^(a[126] & b[391])^(a[125] & b[392])^(a[124] & b[393])^(a[123] & b[394])^(a[122] & b[395])^(a[121] & b[396])^(a[120] & b[397])^(a[119] & b[398])^(a[118] & b[399])^(a[117] & b[400])^(a[116] & b[401])^(a[115] & b[402])^(a[114] & b[403])^(a[113] & b[404])^(a[112] & b[405])^(a[111] & b[406])^(a[110] & b[407])^(a[109] & b[408]);
assign y[518] = (a[408] & b[110])^(a[407] & b[111])^(a[406] & b[112])^(a[405] & b[113])^(a[404] & b[114])^(a[403] & b[115])^(a[402] & b[116])^(a[401] & b[117])^(a[400] & b[118])^(a[399] & b[119])^(a[398] & b[120])^(a[397] & b[121])^(a[396] & b[122])^(a[395] & b[123])^(a[394] & b[124])^(a[393] & b[125])^(a[392] & b[126])^(a[391] & b[127])^(a[390] & b[128])^(a[389] & b[129])^(a[388] & b[130])^(a[387] & b[131])^(a[386] & b[132])^(a[385] & b[133])^(a[384] & b[134])^(a[383] & b[135])^(a[382] & b[136])^(a[381] & b[137])^(a[380] & b[138])^(a[379] & b[139])^(a[378] & b[140])^(a[377] & b[141])^(a[376] & b[142])^(a[375] & b[143])^(a[374] & b[144])^(a[373] & b[145])^(a[372] & b[146])^(a[371] & b[147])^(a[370] & b[148])^(a[369] & b[149])^(a[368] & b[150])^(a[367] & b[151])^(a[366] & b[152])^(a[365] & b[153])^(a[364] & b[154])^(a[363] & b[155])^(a[362] & b[156])^(a[361] & b[157])^(a[360] & b[158])^(a[359] & b[159])^(a[358] & b[160])^(a[357] & b[161])^(a[356] & b[162])^(a[355] & b[163])^(a[354] & b[164])^(a[353] & b[165])^(a[352] & b[166])^(a[351] & b[167])^(a[350] & b[168])^(a[349] & b[169])^(a[348] & b[170])^(a[347] & b[171])^(a[346] & b[172])^(a[345] & b[173])^(a[344] & b[174])^(a[343] & b[175])^(a[342] & b[176])^(a[341] & b[177])^(a[340] & b[178])^(a[339] & b[179])^(a[338] & b[180])^(a[337] & b[181])^(a[336] & b[182])^(a[335] & b[183])^(a[334] & b[184])^(a[333] & b[185])^(a[332] & b[186])^(a[331] & b[187])^(a[330] & b[188])^(a[329] & b[189])^(a[328] & b[190])^(a[327] & b[191])^(a[326] & b[192])^(a[325] & b[193])^(a[324] & b[194])^(a[323] & b[195])^(a[322] & b[196])^(a[321] & b[197])^(a[320] & b[198])^(a[319] & b[199])^(a[318] & b[200])^(a[317] & b[201])^(a[316] & b[202])^(a[315] & b[203])^(a[314] & b[204])^(a[313] & b[205])^(a[312] & b[206])^(a[311] & b[207])^(a[310] & b[208])^(a[309] & b[209])^(a[308] & b[210])^(a[307] & b[211])^(a[306] & b[212])^(a[305] & b[213])^(a[304] & b[214])^(a[303] & b[215])^(a[302] & b[216])^(a[301] & b[217])^(a[300] & b[218])^(a[299] & b[219])^(a[298] & b[220])^(a[297] & b[221])^(a[296] & b[222])^(a[295] & b[223])^(a[294] & b[224])^(a[293] & b[225])^(a[292] & b[226])^(a[291] & b[227])^(a[290] & b[228])^(a[289] & b[229])^(a[288] & b[230])^(a[287] & b[231])^(a[286] & b[232])^(a[285] & b[233])^(a[284] & b[234])^(a[283] & b[235])^(a[282] & b[236])^(a[281] & b[237])^(a[280] & b[238])^(a[279] & b[239])^(a[278] & b[240])^(a[277] & b[241])^(a[276] & b[242])^(a[275] & b[243])^(a[274] & b[244])^(a[273] & b[245])^(a[272] & b[246])^(a[271] & b[247])^(a[270] & b[248])^(a[269] & b[249])^(a[268] & b[250])^(a[267] & b[251])^(a[266] & b[252])^(a[265] & b[253])^(a[264] & b[254])^(a[263] & b[255])^(a[262] & b[256])^(a[261] & b[257])^(a[260] & b[258])^(a[259] & b[259])^(a[258] & b[260])^(a[257] & b[261])^(a[256] & b[262])^(a[255] & b[263])^(a[254] & b[264])^(a[253] & b[265])^(a[252] & b[266])^(a[251] & b[267])^(a[250] & b[268])^(a[249] & b[269])^(a[248] & b[270])^(a[247] & b[271])^(a[246] & b[272])^(a[245] & b[273])^(a[244] & b[274])^(a[243] & b[275])^(a[242] & b[276])^(a[241] & b[277])^(a[240] & b[278])^(a[239] & b[279])^(a[238] & b[280])^(a[237] & b[281])^(a[236] & b[282])^(a[235] & b[283])^(a[234] & b[284])^(a[233] & b[285])^(a[232] & b[286])^(a[231] & b[287])^(a[230] & b[288])^(a[229] & b[289])^(a[228] & b[290])^(a[227] & b[291])^(a[226] & b[292])^(a[225] & b[293])^(a[224] & b[294])^(a[223] & b[295])^(a[222] & b[296])^(a[221] & b[297])^(a[220] & b[298])^(a[219] & b[299])^(a[218] & b[300])^(a[217] & b[301])^(a[216] & b[302])^(a[215] & b[303])^(a[214] & b[304])^(a[213] & b[305])^(a[212] & b[306])^(a[211] & b[307])^(a[210] & b[308])^(a[209] & b[309])^(a[208] & b[310])^(a[207] & b[311])^(a[206] & b[312])^(a[205] & b[313])^(a[204] & b[314])^(a[203] & b[315])^(a[202] & b[316])^(a[201] & b[317])^(a[200] & b[318])^(a[199] & b[319])^(a[198] & b[320])^(a[197] & b[321])^(a[196] & b[322])^(a[195] & b[323])^(a[194] & b[324])^(a[193] & b[325])^(a[192] & b[326])^(a[191] & b[327])^(a[190] & b[328])^(a[189] & b[329])^(a[188] & b[330])^(a[187] & b[331])^(a[186] & b[332])^(a[185] & b[333])^(a[184] & b[334])^(a[183] & b[335])^(a[182] & b[336])^(a[181] & b[337])^(a[180] & b[338])^(a[179] & b[339])^(a[178] & b[340])^(a[177] & b[341])^(a[176] & b[342])^(a[175] & b[343])^(a[174] & b[344])^(a[173] & b[345])^(a[172] & b[346])^(a[171] & b[347])^(a[170] & b[348])^(a[169] & b[349])^(a[168] & b[350])^(a[167] & b[351])^(a[166] & b[352])^(a[165] & b[353])^(a[164] & b[354])^(a[163] & b[355])^(a[162] & b[356])^(a[161] & b[357])^(a[160] & b[358])^(a[159] & b[359])^(a[158] & b[360])^(a[157] & b[361])^(a[156] & b[362])^(a[155] & b[363])^(a[154] & b[364])^(a[153] & b[365])^(a[152] & b[366])^(a[151] & b[367])^(a[150] & b[368])^(a[149] & b[369])^(a[148] & b[370])^(a[147] & b[371])^(a[146] & b[372])^(a[145] & b[373])^(a[144] & b[374])^(a[143] & b[375])^(a[142] & b[376])^(a[141] & b[377])^(a[140] & b[378])^(a[139] & b[379])^(a[138] & b[380])^(a[137] & b[381])^(a[136] & b[382])^(a[135] & b[383])^(a[134] & b[384])^(a[133] & b[385])^(a[132] & b[386])^(a[131] & b[387])^(a[130] & b[388])^(a[129] & b[389])^(a[128] & b[390])^(a[127] & b[391])^(a[126] & b[392])^(a[125] & b[393])^(a[124] & b[394])^(a[123] & b[395])^(a[122] & b[396])^(a[121] & b[397])^(a[120] & b[398])^(a[119] & b[399])^(a[118] & b[400])^(a[117] & b[401])^(a[116] & b[402])^(a[115] & b[403])^(a[114] & b[404])^(a[113] & b[405])^(a[112] & b[406])^(a[111] & b[407])^(a[110] & b[408]);
assign y[519] = (a[408] & b[111])^(a[407] & b[112])^(a[406] & b[113])^(a[405] & b[114])^(a[404] & b[115])^(a[403] & b[116])^(a[402] & b[117])^(a[401] & b[118])^(a[400] & b[119])^(a[399] & b[120])^(a[398] & b[121])^(a[397] & b[122])^(a[396] & b[123])^(a[395] & b[124])^(a[394] & b[125])^(a[393] & b[126])^(a[392] & b[127])^(a[391] & b[128])^(a[390] & b[129])^(a[389] & b[130])^(a[388] & b[131])^(a[387] & b[132])^(a[386] & b[133])^(a[385] & b[134])^(a[384] & b[135])^(a[383] & b[136])^(a[382] & b[137])^(a[381] & b[138])^(a[380] & b[139])^(a[379] & b[140])^(a[378] & b[141])^(a[377] & b[142])^(a[376] & b[143])^(a[375] & b[144])^(a[374] & b[145])^(a[373] & b[146])^(a[372] & b[147])^(a[371] & b[148])^(a[370] & b[149])^(a[369] & b[150])^(a[368] & b[151])^(a[367] & b[152])^(a[366] & b[153])^(a[365] & b[154])^(a[364] & b[155])^(a[363] & b[156])^(a[362] & b[157])^(a[361] & b[158])^(a[360] & b[159])^(a[359] & b[160])^(a[358] & b[161])^(a[357] & b[162])^(a[356] & b[163])^(a[355] & b[164])^(a[354] & b[165])^(a[353] & b[166])^(a[352] & b[167])^(a[351] & b[168])^(a[350] & b[169])^(a[349] & b[170])^(a[348] & b[171])^(a[347] & b[172])^(a[346] & b[173])^(a[345] & b[174])^(a[344] & b[175])^(a[343] & b[176])^(a[342] & b[177])^(a[341] & b[178])^(a[340] & b[179])^(a[339] & b[180])^(a[338] & b[181])^(a[337] & b[182])^(a[336] & b[183])^(a[335] & b[184])^(a[334] & b[185])^(a[333] & b[186])^(a[332] & b[187])^(a[331] & b[188])^(a[330] & b[189])^(a[329] & b[190])^(a[328] & b[191])^(a[327] & b[192])^(a[326] & b[193])^(a[325] & b[194])^(a[324] & b[195])^(a[323] & b[196])^(a[322] & b[197])^(a[321] & b[198])^(a[320] & b[199])^(a[319] & b[200])^(a[318] & b[201])^(a[317] & b[202])^(a[316] & b[203])^(a[315] & b[204])^(a[314] & b[205])^(a[313] & b[206])^(a[312] & b[207])^(a[311] & b[208])^(a[310] & b[209])^(a[309] & b[210])^(a[308] & b[211])^(a[307] & b[212])^(a[306] & b[213])^(a[305] & b[214])^(a[304] & b[215])^(a[303] & b[216])^(a[302] & b[217])^(a[301] & b[218])^(a[300] & b[219])^(a[299] & b[220])^(a[298] & b[221])^(a[297] & b[222])^(a[296] & b[223])^(a[295] & b[224])^(a[294] & b[225])^(a[293] & b[226])^(a[292] & b[227])^(a[291] & b[228])^(a[290] & b[229])^(a[289] & b[230])^(a[288] & b[231])^(a[287] & b[232])^(a[286] & b[233])^(a[285] & b[234])^(a[284] & b[235])^(a[283] & b[236])^(a[282] & b[237])^(a[281] & b[238])^(a[280] & b[239])^(a[279] & b[240])^(a[278] & b[241])^(a[277] & b[242])^(a[276] & b[243])^(a[275] & b[244])^(a[274] & b[245])^(a[273] & b[246])^(a[272] & b[247])^(a[271] & b[248])^(a[270] & b[249])^(a[269] & b[250])^(a[268] & b[251])^(a[267] & b[252])^(a[266] & b[253])^(a[265] & b[254])^(a[264] & b[255])^(a[263] & b[256])^(a[262] & b[257])^(a[261] & b[258])^(a[260] & b[259])^(a[259] & b[260])^(a[258] & b[261])^(a[257] & b[262])^(a[256] & b[263])^(a[255] & b[264])^(a[254] & b[265])^(a[253] & b[266])^(a[252] & b[267])^(a[251] & b[268])^(a[250] & b[269])^(a[249] & b[270])^(a[248] & b[271])^(a[247] & b[272])^(a[246] & b[273])^(a[245] & b[274])^(a[244] & b[275])^(a[243] & b[276])^(a[242] & b[277])^(a[241] & b[278])^(a[240] & b[279])^(a[239] & b[280])^(a[238] & b[281])^(a[237] & b[282])^(a[236] & b[283])^(a[235] & b[284])^(a[234] & b[285])^(a[233] & b[286])^(a[232] & b[287])^(a[231] & b[288])^(a[230] & b[289])^(a[229] & b[290])^(a[228] & b[291])^(a[227] & b[292])^(a[226] & b[293])^(a[225] & b[294])^(a[224] & b[295])^(a[223] & b[296])^(a[222] & b[297])^(a[221] & b[298])^(a[220] & b[299])^(a[219] & b[300])^(a[218] & b[301])^(a[217] & b[302])^(a[216] & b[303])^(a[215] & b[304])^(a[214] & b[305])^(a[213] & b[306])^(a[212] & b[307])^(a[211] & b[308])^(a[210] & b[309])^(a[209] & b[310])^(a[208] & b[311])^(a[207] & b[312])^(a[206] & b[313])^(a[205] & b[314])^(a[204] & b[315])^(a[203] & b[316])^(a[202] & b[317])^(a[201] & b[318])^(a[200] & b[319])^(a[199] & b[320])^(a[198] & b[321])^(a[197] & b[322])^(a[196] & b[323])^(a[195] & b[324])^(a[194] & b[325])^(a[193] & b[326])^(a[192] & b[327])^(a[191] & b[328])^(a[190] & b[329])^(a[189] & b[330])^(a[188] & b[331])^(a[187] & b[332])^(a[186] & b[333])^(a[185] & b[334])^(a[184] & b[335])^(a[183] & b[336])^(a[182] & b[337])^(a[181] & b[338])^(a[180] & b[339])^(a[179] & b[340])^(a[178] & b[341])^(a[177] & b[342])^(a[176] & b[343])^(a[175] & b[344])^(a[174] & b[345])^(a[173] & b[346])^(a[172] & b[347])^(a[171] & b[348])^(a[170] & b[349])^(a[169] & b[350])^(a[168] & b[351])^(a[167] & b[352])^(a[166] & b[353])^(a[165] & b[354])^(a[164] & b[355])^(a[163] & b[356])^(a[162] & b[357])^(a[161] & b[358])^(a[160] & b[359])^(a[159] & b[360])^(a[158] & b[361])^(a[157] & b[362])^(a[156] & b[363])^(a[155] & b[364])^(a[154] & b[365])^(a[153] & b[366])^(a[152] & b[367])^(a[151] & b[368])^(a[150] & b[369])^(a[149] & b[370])^(a[148] & b[371])^(a[147] & b[372])^(a[146] & b[373])^(a[145] & b[374])^(a[144] & b[375])^(a[143] & b[376])^(a[142] & b[377])^(a[141] & b[378])^(a[140] & b[379])^(a[139] & b[380])^(a[138] & b[381])^(a[137] & b[382])^(a[136] & b[383])^(a[135] & b[384])^(a[134] & b[385])^(a[133] & b[386])^(a[132] & b[387])^(a[131] & b[388])^(a[130] & b[389])^(a[129] & b[390])^(a[128] & b[391])^(a[127] & b[392])^(a[126] & b[393])^(a[125] & b[394])^(a[124] & b[395])^(a[123] & b[396])^(a[122] & b[397])^(a[121] & b[398])^(a[120] & b[399])^(a[119] & b[400])^(a[118] & b[401])^(a[117] & b[402])^(a[116] & b[403])^(a[115] & b[404])^(a[114] & b[405])^(a[113] & b[406])^(a[112] & b[407])^(a[111] & b[408]);
assign y[520] = (a[408] & b[112])^(a[407] & b[113])^(a[406] & b[114])^(a[405] & b[115])^(a[404] & b[116])^(a[403] & b[117])^(a[402] & b[118])^(a[401] & b[119])^(a[400] & b[120])^(a[399] & b[121])^(a[398] & b[122])^(a[397] & b[123])^(a[396] & b[124])^(a[395] & b[125])^(a[394] & b[126])^(a[393] & b[127])^(a[392] & b[128])^(a[391] & b[129])^(a[390] & b[130])^(a[389] & b[131])^(a[388] & b[132])^(a[387] & b[133])^(a[386] & b[134])^(a[385] & b[135])^(a[384] & b[136])^(a[383] & b[137])^(a[382] & b[138])^(a[381] & b[139])^(a[380] & b[140])^(a[379] & b[141])^(a[378] & b[142])^(a[377] & b[143])^(a[376] & b[144])^(a[375] & b[145])^(a[374] & b[146])^(a[373] & b[147])^(a[372] & b[148])^(a[371] & b[149])^(a[370] & b[150])^(a[369] & b[151])^(a[368] & b[152])^(a[367] & b[153])^(a[366] & b[154])^(a[365] & b[155])^(a[364] & b[156])^(a[363] & b[157])^(a[362] & b[158])^(a[361] & b[159])^(a[360] & b[160])^(a[359] & b[161])^(a[358] & b[162])^(a[357] & b[163])^(a[356] & b[164])^(a[355] & b[165])^(a[354] & b[166])^(a[353] & b[167])^(a[352] & b[168])^(a[351] & b[169])^(a[350] & b[170])^(a[349] & b[171])^(a[348] & b[172])^(a[347] & b[173])^(a[346] & b[174])^(a[345] & b[175])^(a[344] & b[176])^(a[343] & b[177])^(a[342] & b[178])^(a[341] & b[179])^(a[340] & b[180])^(a[339] & b[181])^(a[338] & b[182])^(a[337] & b[183])^(a[336] & b[184])^(a[335] & b[185])^(a[334] & b[186])^(a[333] & b[187])^(a[332] & b[188])^(a[331] & b[189])^(a[330] & b[190])^(a[329] & b[191])^(a[328] & b[192])^(a[327] & b[193])^(a[326] & b[194])^(a[325] & b[195])^(a[324] & b[196])^(a[323] & b[197])^(a[322] & b[198])^(a[321] & b[199])^(a[320] & b[200])^(a[319] & b[201])^(a[318] & b[202])^(a[317] & b[203])^(a[316] & b[204])^(a[315] & b[205])^(a[314] & b[206])^(a[313] & b[207])^(a[312] & b[208])^(a[311] & b[209])^(a[310] & b[210])^(a[309] & b[211])^(a[308] & b[212])^(a[307] & b[213])^(a[306] & b[214])^(a[305] & b[215])^(a[304] & b[216])^(a[303] & b[217])^(a[302] & b[218])^(a[301] & b[219])^(a[300] & b[220])^(a[299] & b[221])^(a[298] & b[222])^(a[297] & b[223])^(a[296] & b[224])^(a[295] & b[225])^(a[294] & b[226])^(a[293] & b[227])^(a[292] & b[228])^(a[291] & b[229])^(a[290] & b[230])^(a[289] & b[231])^(a[288] & b[232])^(a[287] & b[233])^(a[286] & b[234])^(a[285] & b[235])^(a[284] & b[236])^(a[283] & b[237])^(a[282] & b[238])^(a[281] & b[239])^(a[280] & b[240])^(a[279] & b[241])^(a[278] & b[242])^(a[277] & b[243])^(a[276] & b[244])^(a[275] & b[245])^(a[274] & b[246])^(a[273] & b[247])^(a[272] & b[248])^(a[271] & b[249])^(a[270] & b[250])^(a[269] & b[251])^(a[268] & b[252])^(a[267] & b[253])^(a[266] & b[254])^(a[265] & b[255])^(a[264] & b[256])^(a[263] & b[257])^(a[262] & b[258])^(a[261] & b[259])^(a[260] & b[260])^(a[259] & b[261])^(a[258] & b[262])^(a[257] & b[263])^(a[256] & b[264])^(a[255] & b[265])^(a[254] & b[266])^(a[253] & b[267])^(a[252] & b[268])^(a[251] & b[269])^(a[250] & b[270])^(a[249] & b[271])^(a[248] & b[272])^(a[247] & b[273])^(a[246] & b[274])^(a[245] & b[275])^(a[244] & b[276])^(a[243] & b[277])^(a[242] & b[278])^(a[241] & b[279])^(a[240] & b[280])^(a[239] & b[281])^(a[238] & b[282])^(a[237] & b[283])^(a[236] & b[284])^(a[235] & b[285])^(a[234] & b[286])^(a[233] & b[287])^(a[232] & b[288])^(a[231] & b[289])^(a[230] & b[290])^(a[229] & b[291])^(a[228] & b[292])^(a[227] & b[293])^(a[226] & b[294])^(a[225] & b[295])^(a[224] & b[296])^(a[223] & b[297])^(a[222] & b[298])^(a[221] & b[299])^(a[220] & b[300])^(a[219] & b[301])^(a[218] & b[302])^(a[217] & b[303])^(a[216] & b[304])^(a[215] & b[305])^(a[214] & b[306])^(a[213] & b[307])^(a[212] & b[308])^(a[211] & b[309])^(a[210] & b[310])^(a[209] & b[311])^(a[208] & b[312])^(a[207] & b[313])^(a[206] & b[314])^(a[205] & b[315])^(a[204] & b[316])^(a[203] & b[317])^(a[202] & b[318])^(a[201] & b[319])^(a[200] & b[320])^(a[199] & b[321])^(a[198] & b[322])^(a[197] & b[323])^(a[196] & b[324])^(a[195] & b[325])^(a[194] & b[326])^(a[193] & b[327])^(a[192] & b[328])^(a[191] & b[329])^(a[190] & b[330])^(a[189] & b[331])^(a[188] & b[332])^(a[187] & b[333])^(a[186] & b[334])^(a[185] & b[335])^(a[184] & b[336])^(a[183] & b[337])^(a[182] & b[338])^(a[181] & b[339])^(a[180] & b[340])^(a[179] & b[341])^(a[178] & b[342])^(a[177] & b[343])^(a[176] & b[344])^(a[175] & b[345])^(a[174] & b[346])^(a[173] & b[347])^(a[172] & b[348])^(a[171] & b[349])^(a[170] & b[350])^(a[169] & b[351])^(a[168] & b[352])^(a[167] & b[353])^(a[166] & b[354])^(a[165] & b[355])^(a[164] & b[356])^(a[163] & b[357])^(a[162] & b[358])^(a[161] & b[359])^(a[160] & b[360])^(a[159] & b[361])^(a[158] & b[362])^(a[157] & b[363])^(a[156] & b[364])^(a[155] & b[365])^(a[154] & b[366])^(a[153] & b[367])^(a[152] & b[368])^(a[151] & b[369])^(a[150] & b[370])^(a[149] & b[371])^(a[148] & b[372])^(a[147] & b[373])^(a[146] & b[374])^(a[145] & b[375])^(a[144] & b[376])^(a[143] & b[377])^(a[142] & b[378])^(a[141] & b[379])^(a[140] & b[380])^(a[139] & b[381])^(a[138] & b[382])^(a[137] & b[383])^(a[136] & b[384])^(a[135] & b[385])^(a[134] & b[386])^(a[133] & b[387])^(a[132] & b[388])^(a[131] & b[389])^(a[130] & b[390])^(a[129] & b[391])^(a[128] & b[392])^(a[127] & b[393])^(a[126] & b[394])^(a[125] & b[395])^(a[124] & b[396])^(a[123] & b[397])^(a[122] & b[398])^(a[121] & b[399])^(a[120] & b[400])^(a[119] & b[401])^(a[118] & b[402])^(a[117] & b[403])^(a[116] & b[404])^(a[115] & b[405])^(a[114] & b[406])^(a[113] & b[407])^(a[112] & b[408]);
assign y[521] = (a[408] & b[113])^(a[407] & b[114])^(a[406] & b[115])^(a[405] & b[116])^(a[404] & b[117])^(a[403] & b[118])^(a[402] & b[119])^(a[401] & b[120])^(a[400] & b[121])^(a[399] & b[122])^(a[398] & b[123])^(a[397] & b[124])^(a[396] & b[125])^(a[395] & b[126])^(a[394] & b[127])^(a[393] & b[128])^(a[392] & b[129])^(a[391] & b[130])^(a[390] & b[131])^(a[389] & b[132])^(a[388] & b[133])^(a[387] & b[134])^(a[386] & b[135])^(a[385] & b[136])^(a[384] & b[137])^(a[383] & b[138])^(a[382] & b[139])^(a[381] & b[140])^(a[380] & b[141])^(a[379] & b[142])^(a[378] & b[143])^(a[377] & b[144])^(a[376] & b[145])^(a[375] & b[146])^(a[374] & b[147])^(a[373] & b[148])^(a[372] & b[149])^(a[371] & b[150])^(a[370] & b[151])^(a[369] & b[152])^(a[368] & b[153])^(a[367] & b[154])^(a[366] & b[155])^(a[365] & b[156])^(a[364] & b[157])^(a[363] & b[158])^(a[362] & b[159])^(a[361] & b[160])^(a[360] & b[161])^(a[359] & b[162])^(a[358] & b[163])^(a[357] & b[164])^(a[356] & b[165])^(a[355] & b[166])^(a[354] & b[167])^(a[353] & b[168])^(a[352] & b[169])^(a[351] & b[170])^(a[350] & b[171])^(a[349] & b[172])^(a[348] & b[173])^(a[347] & b[174])^(a[346] & b[175])^(a[345] & b[176])^(a[344] & b[177])^(a[343] & b[178])^(a[342] & b[179])^(a[341] & b[180])^(a[340] & b[181])^(a[339] & b[182])^(a[338] & b[183])^(a[337] & b[184])^(a[336] & b[185])^(a[335] & b[186])^(a[334] & b[187])^(a[333] & b[188])^(a[332] & b[189])^(a[331] & b[190])^(a[330] & b[191])^(a[329] & b[192])^(a[328] & b[193])^(a[327] & b[194])^(a[326] & b[195])^(a[325] & b[196])^(a[324] & b[197])^(a[323] & b[198])^(a[322] & b[199])^(a[321] & b[200])^(a[320] & b[201])^(a[319] & b[202])^(a[318] & b[203])^(a[317] & b[204])^(a[316] & b[205])^(a[315] & b[206])^(a[314] & b[207])^(a[313] & b[208])^(a[312] & b[209])^(a[311] & b[210])^(a[310] & b[211])^(a[309] & b[212])^(a[308] & b[213])^(a[307] & b[214])^(a[306] & b[215])^(a[305] & b[216])^(a[304] & b[217])^(a[303] & b[218])^(a[302] & b[219])^(a[301] & b[220])^(a[300] & b[221])^(a[299] & b[222])^(a[298] & b[223])^(a[297] & b[224])^(a[296] & b[225])^(a[295] & b[226])^(a[294] & b[227])^(a[293] & b[228])^(a[292] & b[229])^(a[291] & b[230])^(a[290] & b[231])^(a[289] & b[232])^(a[288] & b[233])^(a[287] & b[234])^(a[286] & b[235])^(a[285] & b[236])^(a[284] & b[237])^(a[283] & b[238])^(a[282] & b[239])^(a[281] & b[240])^(a[280] & b[241])^(a[279] & b[242])^(a[278] & b[243])^(a[277] & b[244])^(a[276] & b[245])^(a[275] & b[246])^(a[274] & b[247])^(a[273] & b[248])^(a[272] & b[249])^(a[271] & b[250])^(a[270] & b[251])^(a[269] & b[252])^(a[268] & b[253])^(a[267] & b[254])^(a[266] & b[255])^(a[265] & b[256])^(a[264] & b[257])^(a[263] & b[258])^(a[262] & b[259])^(a[261] & b[260])^(a[260] & b[261])^(a[259] & b[262])^(a[258] & b[263])^(a[257] & b[264])^(a[256] & b[265])^(a[255] & b[266])^(a[254] & b[267])^(a[253] & b[268])^(a[252] & b[269])^(a[251] & b[270])^(a[250] & b[271])^(a[249] & b[272])^(a[248] & b[273])^(a[247] & b[274])^(a[246] & b[275])^(a[245] & b[276])^(a[244] & b[277])^(a[243] & b[278])^(a[242] & b[279])^(a[241] & b[280])^(a[240] & b[281])^(a[239] & b[282])^(a[238] & b[283])^(a[237] & b[284])^(a[236] & b[285])^(a[235] & b[286])^(a[234] & b[287])^(a[233] & b[288])^(a[232] & b[289])^(a[231] & b[290])^(a[230] & b[291])^(a[229] & b[292])^(a[228] & b[293])^(a[227] & b[294])^(a[226] & b[295])^(a[225] & b[296])^(a[224] & b[297])^(a[223] & b[298])^(a[222] & b[299])^(a[221] & b[300])^(a[220] & b[301])^(a[219] & b[302])^(a[218] & b[303])^(a[217] & b[304])^(a[216] & b[305])^(a[215] & b[306])^(a[214] & b[307])^(a[213] & b[308])^(a[212] & b[309])^(a[211] & b[310])^(a[210] & b[311])^(a[209] & b[312])^(a[208] & b[313])^(a[207] & b[314])^(a[206] & b[315])^(a[205] & b[316])^(a[204] & b[317])^(a[203] & b[318])^(a[202] & b[319])^(a[201] & b[320])^(a[200] & b[321])^(a[199] & b[322])^(a[198] & b[323])^(a[197] & b[324])^(a[196] & b[325])^(a[195] & b[326])^(a[194] & b[327])^(a[193] & b[328])^(a[192] & b[329])^(a[191] & b[330])^(a[190] & b[331])^(a[189] & b[332])^(a[188] & b[333])^(a[187] & b[334])^(a[186] & b[335])^(a[185] & b[336])^(a[184] & b[337])^(a[183] & b[338])^(a[182] & b[339])^(a[181] & b[340])^(a[180] & b[341])^(a[179] & b[342])^(a[178] & b[343])^(a[177] & b[344])^(a[176] & b[345])^(a[175] & b[346])^(a[174] & b[347])^(a[173] & b[348])^(a[172] & b[349])^(a[171] & b[350])^(a[170] & b[351])^(a[169] & b[352])^(a[168] & b[353])^(a[167] & b[354])^(a[166] & b[355])^(a[165] & b[356])^(a[164] & b[357])^(a[163] & b[358])^(a[162] & b[359])^(a[161] & b[360])^(a[160] & b[361])^(a[159] & b[362])^(a[158] & b[363])^(a[157] & b[364])^(a[156] & b[365])^(a[155] & b[366])^(a[154] & b[367])^(a[153] & b[368])^(a[152] & b[369])^(a[151] & b[370])^(a[150] & b[371])^(a[149] & b[372])^(a[148] & b[373])^(a[147] & b[374])^(a[146] & b[375])^(a[145] & b[376])^(a[144] & b[377])^(a[143] & b[378])^(a[142] & b[379])^(a[141] & b[380])^(a[140] & b[381])^(a[139] & b[382])^(a[138] & b[383])^(a[137] & b[384])^(a[136] & b[385])^(a[135] & b[386])^(a[134] & b[387])^(a[133] & b[388])^(a[132] & b[389])^(a[131] & b[390])^(a[130] & b[391])^(a[129] & b[392])^(a[128] & b[393])^(a[127] & b[394])^(a[126] & b[395])^(a[125] & b[396])^(a[124] & b[397])^(a[123] & b[398])^(a[122] & b[399])^(a[121] & b[400])^(a[120] & b[401])^(a[119] & b[402])^(a[118] & b[403])^(a[117] & b[404])^(a[116] & b[405])^(a[115] & b[406])^(a[114] & b[407])^(a[113] & b[408]);
assign y[522] = (a[408] & b[114])^(a[407] & b[115])^(a[406] & b[116])^(a[405] & b[117])^(a[404] & b[118])^(a[403] & b[119])^(a[402] & b[120])^(a[401] & b[121])^(a[400] & b[122])^(a[399] & b[123])^(a[398] & b[124])^(a[397] & b[125])^(a[396] & b[126])^(a[395] & b[127])^(a[394] & b[128])^(a[393] & b[129])^(a[392] & b[130])^(a[391] & b[131])^(a[390] & b[132])^(a[389] & b[133])^(a[388] & b[134])^(a[387] & b[135])^(a[386] & b[136])^(a[385] & b[137])^(a[384] & b[138])^(a[383] & b[139])^(a[382] & b[140])^(a[381] & b[141])^(a[380] & b[142])^(a[379] & b[143])^(a[378] & b[144])^(a[377] & b[145])^(a[376] & b[146])^(a[375] & b[147])^(a[374] & b[148])^(a[373] & b[149])^(a[372] & b[150])^(a[371] & b[151])^(a[370] & b[152])^(a[369] & b[153])^(a[368] & b[154])^(a[367] & b[155])^(a[366] & b[156])^(a[365] & b[157])^(a[364] & b[158])^(a[363] & b[159])^(a[362] & b[160])^(a[361] & b[161])^(a[360] & b[162])^(a[359] & b[163])^(a[358] & b[164])^(a[357] & b[165])^(a[356] & b[166])^(a[355] & b[167])^(a[354] & b[168])^(a[353] & b[169])^(a[352] & b[170])^(a[351] & b[171])^(a[350] & b[172])^(a[349] & b[173])^(a[348] & b[174])^(a[347] & b[175])^(a[346] & b[176])^(a[345] & b[177])^(a[344] & b[178])^(a[343] & b[179])^(a[342] & b[180])^(a[341] & b[181])^(a[340] & b[182])^(a[339] & b[183])^(a[338] & b[184])^(a[337] & b[185])^(a[336] & b[186])^(a[335] & b[187])^(a[334] & b[188])^(a[333] & b[189])^(a[332] & b[190])^(a[331] & b[191])^(a[330] & b[192])^(a[329] & b[193])^(a[328] & b[194])^(a[327] & b[195])^(a[326] & b[196])^(a[325] & b[197])^(a[324] & b[198])^(a[323] & b[199])^(a[322] & b[200])^(a[321] & b[201])^(a[320] & b[202])^(a[319] & b[203])^(a[318] & b[204])^(a[317] & b[205])^(a[316] & b[206])^(a[315] & b[207])^(a[314] & b[208])^(a[313] & b[209])^(a[312] & b[210])^(a[311] & b[211])^(a[310] & b[212])^(a[309] & b[213])^(a[308] & b[214])^(a[307] & b[215])^(a[306] & b[216])^(a[305] & b[217])^(a[304] & b[218])^(a[303] & b[219])^(a[302] & b[220])^(a[301] & b[221])^(a[300] & b[222])^(a[299] & b[223])^(a[298] & b[224])^(a[297] & b[225])^(a[296] & b[226])^(a[295] & b[227])^(a[294] & b[228])^(a[293] & b[229])^(a[292] & b[230])^(a[291] & b[231])^(a[290] & b[232])^(a[289] & b[233])^(a[288] & b[234])^(a[287] & b[235])^(a[286] & b[236])^(a[285] & b[237])^(a[284] & b[238])^(a[283] & b[239])^(a[282] & b[240])^(a[281] & b[241])^(a[280] & b[242])^(a[279] & b[243])^(a[278] & b[244])^(a[277] & b[245])^(a[276] & b[246])^(a[275] & b[247])^(a[274] & b[248])^(a[273] & b[249])^(a[272] & b[250])^(a[271] & b[251])^(a[270] & b[252])^(a[269] & b[253])^(a[268] & b[254])^(a[267] & b[255])^(a[266] & b[256])^(a[265] & b[257])^(a[264] & b[258])^(a[263] & b[259])^(a[262] & b[260])^(a[261] & b[261])^(a[260] & b[262])^(a[259] & b[263])^(a[258] & b[264])^(a[257] & b[265])^(a[256] & b[266])^(a[255] & b[267])^(a[254] & b[268])^(a[253] & b[269])^(a[252] & b[270])^(a[251] & b[271])^(a[250] & b[272])^(a[249] & b[273])^(a[248] & b[274])^(a[247] & b[275])^(a[246] & b[276])^(a[245] & b[277])^(a[244] & b[278])^(a[243] & b[279])^(a[242] & b[280])^(a[241] & b[281])^(a[240] & b[282])^(a[239] & b[283])^(a[238] & b[284])^(a[237] & b[285])^(a[236] & b[286])^(a[235] & b[287])^(a[234] & b[288])^(a[233] & b[289])^(a[232] & b[290])^(a[231] & b[291])^(a[230] & b[292])^(a[229] & b[293])^(a[228] & b[294])^(a[227] & b[295])^(a[226] & b[296])^(a[225] & b[297])^(a[224] & b[298])^(a[223] & b[299])^(a[222] & b[300])^(a[221] & b[301])^(a[220] & b[302])^(a[219] & b[303])^(a[218] & b[304])^(a[217] & b[305])^(a[216] & b[306])^(a[215] & b[307])^(a[214] & b[308])^(a[213] & b[309])^(a[212] & b[310])^(a[211] & b[311])^(a[210] & b[312])^(a[209] & b[313])^(a[208] & b[314])^(a[207] & b[315])^(a[206] & b[316])^(a[205] & b[317])^(a[204] & b[318])^(a[203] & b[319])^(a[202] & b[320])^(a[201] & b[321])^(a[200] & b[322])^(a[199] & b[323])^(a[198] & b[324])^(a[197] & b[325])^(a[196] & b[326])^(a[195] & b[327])^(a[194] & b[328])^(a[193] & b[329])^(a[192] & b[330])^(a[191] & b[331])^(a[190] & b[332])^(a[189] & b[333])^(a[188] & b[334])^(a[187] & b[335])^(a[186] & b[336])^(a[185] & b[337])^(a[184] & b[338])^(a[183] & b[339])^(a[182] & b[340])^(a[181] & b[341])^(a[180] & b[342])^(a[179] & b[343])^(a[178] & b[344])^(a[177] & b[345])^(a[176] & b[346])^(a[175] & b[347])^(a[174] & b[348])^(a[173] & b[349])^(a[172] & b[350])^(a[171] & b[351])^(a[170] & b[352])^(a[169] & b[353])^(a[168] & b[354])^(a[167] & b[355])^(a[166] & b[356])^(a[165] & b[357])^(a[164] & b[358])^(a[163] & b[359])^(a[162] & b[360])^(a[161] & b[361])^(a[160] & b[362])^(a[159] & b[363])^(a[158] & b[364])^(a[157] & b[365])^(a[156] & b[366])^(a[155] & b[367])^(a[154] & b[368])^(a[153] & b[369])^(a[152] & b[370])^(a[151] & b[371])^(a[150] & b[372])^(a[149] & b[373])^(a[148] & b[374])^(a[147] & b[375])^(a[146] & b[376])^(a[145] & b[377])^(a[144] & b[378])^(a[143] & b[379])^(a[142] & b[380])^(a[141] & b[381])^(a[140] & b[382])^(a[139] & b[383])^(a[138] & b[384])^(a[137] & b[385])^(a[136] & b[386])^(a[135] & b[387])^(a[134] & b[388])^(a[133] & b[389])^(a[132] & b[390])^(a[131] & b[391])^(a[130] & b[392])^(a[129] & b[393])^(a[128] & b[394])^(a[127] & b[395])^(a[126] & b[396])^(a[125] & b[397])^(a[124] & b[398])^(a[123] & b[399])^(a[122] & b[400])^(a[121] & b[401])^(a[120] & b[402])^(a[119] & b[403])^(a[118] & b[404])^(a[117] & b[405])^(a[116] & b[406])^(a[115] & b[407])^(a[114] & b[408]);
assign y[523] = (a[408] & b[115])^(a[407] & b[116])^(a[406] & b[117])^(a[405] & b[118])^(a[404] & b[119])^(a[403] & b[120])^(a[402] & b[121])^(a[401] & b[122])^(a[400] & b[123])^(a[399] & b[124])^(a[398] & b[125])^(a[397] & b[126])^(a[396] & b[127])^(a[395] & b[128])^(a[394] & b[129])^(a[393] & b[130])^(a[392] & b[131])^(a[391] & b[132])^(a[390] & b[133])^(a[389] & b[134])^(a[388] & b[135])^(a[387] & b[136])^(a[386] & b[137])^(a[385] & b[138])^(a[384] & b[139])^(a[383] & b[140])^(a[382] & b[141])^(a[381] & b[142])^(a[380] & b[143])^(a[379] & b[144])^(a[378] & b[145])^(a[377] & b[146])^(a[376] & b[147])^(a[375] & b[148])^(a[374] & b[149])^(a[373] & b[150])^(a[372] & b[151])^(a[371] & b[152])^(a[370] & b[153])^(a[369] & b[154])^(a[368] & b[155])^(a[367] & b[156])^(a[366] & b[157])^(a[365] & b[158])^(a[364] & b[159])^(a[363] & b[160])^(a[362] & b[161])^(a[361] & b[162])^(a[360] & b[163])^(a[359] & b[164])^(a[358] & b[165])^(a[357] & b[166])^(a[356] & b[167])^(a[355] & b[168])^(a[354] & b[169])^(a[353] & b[170])^(a[352] & b[171])^(a[351] & b[172])^(a[350] & b[173])^(a[349] & b[174])^(a[348] & b[175])^(a[347] & b[176])^(a[346] & b[177])^(a[345] & b[178])^(a[344] & b[179])^(a[343] & b[180])^(a[342] & b[181])^(a[341] & b[182])^(a[340] & b[183])^(a[339] & b[184])^(a[338] & b[185])^(a[337] & b[186])^(a[336] & b[187])^(a[335] & b[188])^(a[334] & b[189])^(a[333] & b[190])^(a[332] & b[191])^(a[331] & b[192])^(a[330] & b[193])^(a[329] & b[194])^(a[328] & b[195])^(a[327] & b[196])^(a[326] & b[197])^(a[325] & b[198])^(a[324] & b[199])^(a[323] & b[200])^(a[322] & b[201])^(a[321] & b[202])^(a[320] & b[203])^(a[319] & b[204])^(a[318] & b[205])^(a[317] & b[206])^(a[316] & b[207])^(a[315] & b[208])^(a[314] & b[209])^(a[313] & b[210])^(a[312] & b[211])^(a[311] & b[212])^(a[310] & b[213])^(a[309] & b[214])^(a[308] & b[215])^(a[307] & b[216])^(a[306] & b[217])^(a[305] & b[218])^(a[304] & b[219])^(a[303] & b[220])^(a[302] & b[221])^(a[301] & b[222])^(a[300] & b[223])^(a[299] & b[224])^(a[298] & b[225])^(a[297] & b[226])^(a[296] & b[227])^(a[295] & b[228])^(a[294] & b[229])^(a[293] & b[230])^(a[292] & b[231])^(a[291] & b[232])^(a[290] & b[233])^(a[289] & b[234])^(a[288] & b[235])^(a[287] & b[236])^(a[286] & b[237])^(a[285] & b[238])^(a[284] & b[239])^(a[283] & b[240])^(a[282] & b[241])^(a[281] & b[242])^(a[280] & b[243])^(a[279] & b[244])^(a[278] & b[245])^(a[277] & b[246])^(a[276] & b[247])^(a[275] & b[248])^(a[274] & b[249])^(a[273] & b[250])^(a[272] & b[251])^(a[271] & b[252])^(a[270] & b[253])^(a[269] & b[254])^(a[268] & b[255])^(a[267] & b[256])^(a[266] & b[257])^(a[265] & b[258])^(a[264] & b[259])^(a[263] & b[260])^(a[262] & b[261])^(a[261] & b[262])^(a[260] & b[263])^(a[259] & b[264])^(a[258] & b[265])^(a[257] & b[266])^(a[256] & b[267])^(a[255] & b[268])^(a[254] & b[269])^(a[253] & b[270])^(a[252] & b[271])^(a[251] & b[272])^(a[250] & b[273])^(a[249] & b[274])^(a[248] & b[275])^(a[247] & b[276])^(a[246] & b[277])^(a[245] & b[278])^(a[244] & b[279])^(a[243] & b[280])^(a[242] & b[281])^(a[241] & b[282])^(a[240] & b[283])^(a[239] & b[284])^(a[238] & b[285])^(a[237] & b[286])^(a[236] & b[287])^(a[235] & b[288])^(a[234] & b[289])^(a[233] & b[290])^(a[232] & b[291])^(a[231] & b[292])^(a[230] & b[293])^(a[229] & b[294])^(a[228] & b[295])^(a[227] & b[296])^(a[226] & b[297])^(a[225] & b[298])^(a[224] & b[299])^(a[223] & b[300])^(a[222] & b[301])^(a[221] & b[302])^(a[220] & b[303])^(a[219] & b[304])^(a[218] & b[305])^(a[217] & b[306])^(a[216] & b[307])^(a[215] & b[308])^(a[214] & b[309])^(a[213] & b[310])^(a[212] & b[311])^(a[211] & b[312])^(a[210] & b[313])^(a[209] & b[314])^(a[208] & b[315])^(a[207] & b[316])^(a[206] & b[317])^(a[205] & b[318])^(a[204] & b[319])^(a[203] & b[320])^(a[202] & b[321])^(a[201] & b[322])^(a[200] & b[323])^(a[199] & b[324])^(a[198] & b[325])^(a[197] & b[326])^(a[196] & b[327])^(a[195] & b[328])^(a[194] & b[329])^(a[193] & b[330])^(a[192] & b[331])^(a[191] & b[332])^(a[190] & b[333])^(a[189] & b[334])^(a[188] & b[335])^(a[187] & b[336])^(a[186] & b[337])^(a[185] & b[338])^(a[184] & b[339])^(a[183] & b[340])^(a[182] & b[341])^(a[181] & b[342])^(a[180] & b[343])^(a[179] & b[344])^(a[178] & b[345])^(a[177] & b[346])^(a[176] & b[347])^(a[175] & b[348])^(a[174] & b[349])^(a[173] & b[350])^(a[172] & b[351])^(a[171] & b[352])^(a[170] & b[353])^(a[169] & b[354])^(a[168] & b[355])^(a[167] & b[356])^(a[166] & b[357])^(a[165] & b[358])^(a[164] & b[359])^(a[163] & b[360])^(a[162] & b[361])^(a[161] & b[362])^(a[160] & b[363])^(a[159] & b[364])^(a[158] & b[365])^(a[157] & b[366])^(a[156] & b[367])^(a[155] & b[368])^(a[154] & b[369])^(a[153] & b[370])^(a[152] & b[371])^(a[151] & b[372])^(a[150] & b[373])^(a[149] & b[374])^(a[148] & b[375])^(a[147] & b[376])^(a[146] & b[377])^(a[145] & b[378])^(a[144] & b[379])^(a[143] & b[380])^(a[142] & b[381])^(a[141] & b[382])^(a[140] & b[383])^(a[139] & b[384])^(a[138] & b[385])^(a[137] & b[386])^(a[136] & b[387])^(a[135] & b[388])^(a[134] & b[389])^(a[133] & b[390])^(a[132] & b[391])^(a[131] & b[392])^(a[130] & b[393])^(a[129] & b[394])^(a[128] & b[395])^(a[127] & b[396])^(a[126] & b[397])^(a[125] & b[398])^(a[124] & b[399])^(a[123] & b[400])^(a[122] & b[401])^(a[121] & b[402])^(a[120] & b[403])^(a[119] & b[404])^(a[118] & b[405])^(a[117] & b[406])^(a[116] & b[407])^(a[115] & b[408]);
assign y[524] = (a[408] & b[116])^(a[407] & b[117])^(a[406] & b[118])^(a[405] & b[119])^(a[404] & b[120])^(a[403] & b[121])^(a[402] & b[122])^(a[401] & b[123])^(a[400] & b[124])^(a[399] & b[125])^(a[398] & b[126])^(a[397] & b[127])^(a[396] & b[128])^(a[395] & b[129])^(a[394] & b[130])^(a[393] & b[131])^(a[392] & b[132])^(a[391] & b[133])^(a[390] & b[134])^(a[389] & b[135])^(a[388] & b[136])^(a[387] & b[137])^(a[386] & b[138])^(a[385] & b[139])^(a[384] & b[140])^(a[383] & b[141])^(a[382] & b[142])^(a[381] & b[143])^(a[380] & b[144])^(a[379] & b[145])^(a[378] & b[146])^(a[377] & b[147])^(a[376] & b[148])^(a[375] & b[149])^(a[374] & b[150])^(a[373] & b[151])^(a[372] & b[152])^(a[371] & b[153])^(a[370] & b[154])^(a[369] & b[155])^(a[368] & b[156])^(a[367] & b[157])^(a[366] & b[158])^(a[365] & b[159])^(a[364] & b[160])^(a[363] & b[161])^(a[362] & b[162])^(a[361] & b[163])^(a[360] & b[164])^(a[359] & b[165])^(a[358] & b[166])^(a[357] & b[167])^(a[356] & b[168])^(a[355] & b[169])^(a[354] & b[170])^(a[353] & b[171])^(a[352] & b[172])^(a[351] & b[173])^(a[350] & b[174])^(a[349] & b[175])^(a[348] & b[176])^(a[347] & b[177])^(a[346] & b[178])^(a[345] & b[179])^(a[344] & b[180])^(a[343] & b[181])^(a[342] & b[182])^(a[341] & b[183])^(a[340] & b[184])^(a[339] & b[185])^(a[338] & b[186])^(a[337] & b[187])^(a[336] & b[188])^(a[335] & b[189])^(a[334] & b[190])^(a[333] & b[191])^(a[332] & b[192])^(a[331] & b[193])^(a[330] & b[194])^(a[329] & b[195])^(a[328] & b[196])^(a[327] & b[197])^(a[326] & b[198])^(a[325] & b[199])^(a[324] & b[200])^(a[323] & b[201])^(a[322] & b[202])^(a[321] & b[203])^(a[320] & b[204])^(a[319] & b[205])^(a[318] & b[206])^(a[317] & b[207])^(a[316] & b[208])^(a[315] & b[209])^(a[314] & b[210])^(a[313] & b[211])^(a[312] & b[212])^(a[311] & b[213])^(a[310] & b[214])^(a[309] & b[215])^(a[308] & b[216])^(a[307] & b[217])^(a[306] & b[218])^(a[305] & b[219])^(a[304] & b[220])^(a[303] & b[221])^(a[302] & b[222])^(a[301] & b[223])^(a[300] & b[224])^(a[299] & b[225])^(a[298] & b[226])^(a[297] & b[227])^(a[296] & b[228])^(a[295] & b[229])^(a[294] & b[230])^(a[293] & b[231])^(a[292] & b[232])^(a[291] & b[233])^(a[290] & b[234])^(a[289] & b[235])^(a[288] & b[236])^(a[287] & b[237])^(a[286] & b[238])^(a[285] & b[239])^(a[284] & b[240])^(a[283] & b[241])^(a[282] & b[242])^(a[281] & b[243])^(a[280] & b[244])^(a[279] & b[245])^(a[278] & b[246])^(a[277] & b[247])^(a[276] & b[248])^(a[275] & b[249])^(a[274] & b[250])^(a[273] & b[251])^(a[272] & b[252])^(a[271] & b[253])^(a[270] & b[254])^(a[269] & b[255])^(a[268] & b[256])^(a[267] & b[257])^(a[266] & b[258])^(a[265] & b[259])^(a[264] & b[260])^(a[263] & b[261])^(a[262] & b[262])^(a[261] & b[263])^(a[260] & b[264])^(a[259] & b[265])^(a[258] & b[266])^(a[257] & b[267])^(a[256] & b[268])^(a[255] & b[269])^(a[254] & b[270])^(a[253] & b[271])^(a[252] & b[272])^(a[251] & b[273])^(a[250] & b[274])^(a[249] & b[275])^(a[248] & b[276])^(a[247] & b[277])^(a[246] & b[278])^(a[245] & b[279])^(a[244] & b[280])^(a[243] & b[281])^(a[242] & b[282])^(a[241] & b[283])^(a[240] & b[284])^(a[239] & b[285])^(a[238] & b[286])^(a[237] & b[287])^(a[236] & b[288])^(a[235] & b[289])^(a[234] & b[290])^(a[233] & b[291])^(a[232] & b[292])^(a[231] & b[293])^(a[230] & b[294])^(a[229] & b[295])^(a[228] & b[296])^(a[227] & b[297])^(a[226] & b[298])^(a[225] & b[299])^(a[224] & b[300])^(a[223] & b[301])^(a[222] & b[302])^(a[221] & b[303])^(a[220] & b[304])^(a[219] & b[305])^(a[218] & b[306])^(a[217] & b[307])^(a[216] & b[308])^(a[215] & b[309])^(a[214] & b[310])^(a[213] & b[311])^(a[212] & b[312])^(a[211] & b[313])^(a[210] & b[314])^(a[209] & b[315])^(a[208] & b[316])^(a[207] & b[317])^(a[206] & b[318])^(a[205] & b[319])^(a[204] & b[320])^(a[203] & b[321])^(a[202] & b[322])^(a[201] & b[323])^(a[200] & b[324])^(a[199] & b[325])^(a[198] & b[326])^(a[197] & b[327])^(a[196] & b[328])^(a[195] & b[329])^(a[194] & b[330])^(a[193] & b[331])^(a[192] & b[332])^(a[191] & b[333])^(a[190] & b[334])^(a[189] & b[335])^(a[188] & b[336])^(a[187] & b[337])^(a[186] & b[338])^(a[185] & b[339])^(a[184] & b[340])^(a[183] & b[341])^(a[182] & b[342])^(a[181] & b[343])^(a[180] & b[344])^(a[179] & b[345])^(a[178] & b[346])^(a[177] & b[347])^(a[176] & b[348])^(a[175] & b[349])^(a[174] & b[350])^(a[173] & b[351])^(a[172] & b[352])^(a[171] & b[353])^(a[170] & b[354])^(a[169] & b[355])^(a[168] & b[356])^(a[167] & b[357])^(a[166] & b[358])^(a[165] & b[359])^(a[164] & b[360])^(a[163] & b[361])^(a[162] & b[362])^(a[161] & b[363])^(a[160] & b[364])^(a[159] & b[365])^(a[158] & b[366])^(a[157] & b[367])^(a[156] & b[368])^(a[155] & b[369])^(a[154] & b[370])^(a[153] & b[371])^(a[152] & b[372])^(a[151] & b[373])^(a[150] & b[374])^(a[149] & b[375])^(a[148] & b[376])^(a[147] & b[377])^(a[146] & b[378])^(a[145] & b[379])^(a[144] & b[380])^(a[143] & b[381])^(a[142] & b[382])^(a[141] & b[383])^(a[140] & b[384])^(a[139] & b[385])^(a[138] & b[386])^(a[137] & b[387])^(a[136] & b[388])^(a[135] & b[389])^(a[134] & b[390])^(a[133] & b[391])^(a[132] & b[392])^(a[131] & b[393])^(a[130] & b[394])^(a[129] & b[395])^(a[128] & b[396])^(a[127] & b[397])^(a[126] & b[398])^(a[125] & b[399])^(a[124] & b[400])^(a[123] & b[401])^(a[122] & b[402])^(a[121] & b[403])^(a[120] & b[404])^(a[119] & b[405])^(a[118] & b[406])^(a[117] & b[407])^(a[116] & b[408]);
assign y[525] = (a[408] & b[117])^(a[407] & b[118])^(a[406] & b[119])^(a[405] & b[120])^(a[404] & b[121])^(a[403] & b[122])^(a[402] & b[123])^(a[401] & b[124])^(a[400] & b[125])^(a[399] & b[126])^(a[398] & b[127])^(a[397] & b[128])^(a[396] & b[129])^(a[395] & b[130])^(a[394] & b[131])^(a[393] & b[132])^(a[392] & b[133])^(a[391] & b[134])^(a[390] & b[135])^(a[389] & b[136])^(a[388] & b[137])^(a[387] & b[138])^(a[386] & b[139])^(a[385] & b[140])^(a[384] & b[141])^(a[383] & b[142])^(a[382] & b[143])^(a[381] & b[144])^(a[380] & b[145])^(a[379] & b[146])^(a[378] & b[147])^(a[377] & b[148])^(a[376] & b[149])^(a[375] & b[150])^(a[374] & b[151])^(a[373] & b[152])^(a[372] & b[153])^(a[371] & b[154])^(a[370] & b[155])^(a[369] & b[156])^(a[368] & b[157])^(a[367] & b[158])^(a[366] & b[159])^(a[365] & b[160])^(a[364] & b[161])^(a[363] & b[162])^(a[362] & b[163])^(a[361] & b[164])^(a[360] & b[165])^(a[359] & b[166])^(a[358] & b[167])^(a[357] & b[168])^(a[356] & b[169])^(a[355] & b[170])^(a[354] & b[171])^(a[353] & b[172])^(a[352] & b[173])^(a[351] & b[174])^(a[350] & b[175])^(a[349] & b[176])^(a[348] & b[177])^(a[347] & b[178])^(a[346] & b[179])^(a[345] & b[180])^(a[344] & b[181])^(a[343] & b[182])^(a[342] & b[183])^(a[341] & b[184])^(a[340] & b[185])^(a[339] & b[186])^(a[338] & b[187])^(a[337] & b[188])^(a[336] & b[189])^(a[335] & b[190])^(a[334] & b[191])^(a[333] & b[192])^(a[332] & b[193])^(a[331] & b[194])^(a[330] & b[195])^(a[329] & b[196])^(a[328] & b[197])^(a[327] & b[198])^(a[326] & b[199])^(a[325] & b[200])^(a[324] & b[201])^(a[323] & b[202])^(a[322] & b[203])^(a[321] & b[204])^(a[320] & b[205])^(a[319] & b[206])^(a[318] & b[207])^(a[317] & b[208])^(a[316] & b[209])^(a[315] & b[210])^(a[314] & b[211])^(a[313] & b[212])^(a[312] & b[213])^(a[311] & b[214])^(a[310] & b[215])^(a[309] & b[216])^(a[308] & b[217])^(a[307] & b[218])^(a[306] & b[219])^(a[305] & b[220])^(a[304] & b[221])^(a[303] & b[222])^(a[302] & b[223])^(a[301] & b[224])^(a[300] & b[225])^(a[299] & b[226])^(a[298] & b[227])^(a[297] & b[228])^(a[296] & b[229])^(a[295] & b[230])^(a[294] & b[231])^(a[293] & b[232])^(a[292] & b[233])^(a[291] & b[234])^(a[290] & b[235])^(a[289] & b[236])^(a[288] & b[237])^(a[287] & b[238])^(a[286] & b[239])^(a[285] & b[240])^(a[284] & b[241])^(a[283] & b[242])^(a[282] & b[243])^(a[281] & b[244])^(a[280] & b[245])^(a[279] & b[246])^(a[278] & b[247])^(a[277] & b[248])^(a[276] & b[249])^(a[275] & b[250])^(a[274] & b[251])^(a[273] & b[252])^(a[272] & b[253])^(a[271] & b[254])^(a[270] & b[255])^(a[269] & b[256])^(a[268] & b[257])^(a[267] & b[258])^(a[266] & b[259])^(a[265] & b[260])^(a[264] & b[261])^(a[263] & b[262])^(a[262] & b[263])^(a[261] & b[264])^(a[260] & b[265])^(a[259] & b[266])^(a[258] & b[267])^(a[257] & b[268])^(a[256] & b[269])^(a[255] & b[270])^(a[254] & b[271])^(a[253] & b[272])^(a[252] & b[273])^(a[251] & b[274])^(a[250] & b[275])^(a[249] & b[276])^(a[248] & b[277])^(a[247] & b[278])^(a[246] & b[279])^(a[245] & b[280])^(a[244] & b[281])^(a[243] & b[282])^(a[242] & b[283])^(a[241] & b[284])^(a[240] & b[285])^(a[239] & b[286])^(a[238] & b[287])^(a[237] & b[288])^(a[236] & b[289])^(a[235] & b[290])^(a[234] & b[291])^(a[233] & b[292])^(a[232] & b[293])^(a[231] & b[294])^(a[230] & b[295])^(a[229] & b[296])^(a[228] & b[297])^(a[227] & b[298])^(a[226] & b[299])^(a[225] & b[300])^(a[224] & b[301])^(a[223] & b[302])^(a[222] & b[303])^(a[221] & b[304])^(a[220] & b[305])^(a[219] & b[306])^(a[218] & b[307])^(a[217] & b[308])^(a[216] & b[309])^(a[215] & b[310])^(a[214] & b[311])^(a[213] & b[312])^(a[212] & b[313])^(a[211] & b[314])^(a[210] & b[315])^(a[209] & b[316])^(a[208] & b[317])^(a[207] & b[318])^(a[206] & b[319])^(a[205] & b[320])^(a[204] & b[321])^(a[203] & b[322])^(a[202] & b[323])^(a[201] & b[324])^(a[200] & b[325])^(a[199] & b[326])^(a[198] & b[327])^(a[197] & b[328])^(a[196] & b[329])^(a[195] & b[330])^(a[194] & b[331])^(a[193] & b[332])^(a[192] & b[333])^(a[191] & b[334])^(a[190] & b[335])^(a[189] & b[336])^(a[188] & b[337])^(a[187] & b[338])^(a[186] & b[339])^(a[185] & b[340])^(a[184] & b[341])^(a[183] & b[342])^(a[182] & b[343])^(a[181] & b[344])^(a[180] & b[345])^(a[179] & b[346])^(a[178] & b[347])^(a[177] & b[348])^(a[176] & b[349])^(a[175] & b[350])^(a[174] & b[351])^(a[173] & b[352])^(a[172] & b[353])^(a[171] & b[354])^(a[170] & b[355])^(a[169] & b[356])^(a[168] & b[357])^(a[167] & b[358])^(a[166] & b[359])^(a[165] & b[360])^(a[164] & b[361])^(a[163] & b[362])^(a[162] & b[363])^(a[161] & b[364])^(a[160] & b[365])^(a[159] & b[366])^(a[158] & b[367])^(a[157] & b[368])^(a[156] & b[369])^(a[155] & b[370])^(a[154] & b[371])^(a[153] & b[372])^(a[152] & b[373])^(a[151] & b[374])^(a[150] & b[375])^(a[149] & b[376])^(a[148] & b[377])^(a[147] & b[378])^(a[146] & b[379])^(a[145] & b[380])^(a[144] & b[381])^(a[143] & b[382])^(a[142] & b[383])^(a[141] & b[384])^(a[140] & b[385])^(a[139] & b[386])^(a[138] & b[387])^(a[137] & b[388])^(a[136] & b[389])^(a[135] & b[390])^(a[134] & b[391])^(a[133] & b[392])^(a[132] & b[393])^(a[131] & b[394])^(a[130] & b[395])^(a[129] & b[396])^(a[128] & b[397])^(a[127] & b[398])^(a[126] & b[399])^(a[125] & b[400])^(a[124] & b[401])^(a[123] & b[402])^(a[122] & b[403])^(a[121] & b[404])^(a[120] & b[405])^(a[119] & b[406])^(a[118] & b[407])^(a[117] & b[408]);
assign y[526] = (a[408] & b[118])^(a[407] & b[119])^(a[406] & b[120])^(a[405] & b[121])^(a[404] & b[122])^(a[403] & b[123])^(a[402] & b[124])^(a[401] & b[125])^(a[400] & b[126])^(a[399] & b[127])^(a[398] & b[128])^(a[397] & b[129])^(a[396] & b[130])^(a[395] & b[131])^(a[394] & b[132])^(a[393] & b[133])^(a[392] & b[134])^(a[391] & b[135])^(a[390] & b[136])^(a[389] & b[137])^(a[388] & b[138])^(a[387] & b[139])^(a[386] & b[140])^(a[385] & b[141])^(a[384] & b[142])^(a[383] & b[143])^(a[382] & b[144])^(a[381] & b[145])^(a[380] & b[146])^(a[379] & b[147])^(a[378] & b[148])^(a[377] & b[149])^(a[376] & b[150])^(a[375] & b[151])^(a[374] & b[152])^(a[373] & b[153])^(a[372] & b[154])^(a[371] & b[155])^(a[370] & b[156])^(a[369] & b[157])^(a[368] & b[158])^(a[367] & b[159])^(a[366] & b[160])^(a[365] & b[161])^(a[364] & b[162])^(a[363] & b[163])^(a[362] & b[164])^(a[361] & b[165])^(a[360] & b[166])^(a[359] & b[167])^(a[358] & b[168])^(a[357] & b[169])^(a[356] & b[170])^(a[355] & b[171])^(a[354] & b[172])^(a[353] & b[173])^(a[352] & b[174])^(a[351] & b[175])^(a[350] & b[176])^(a[349] & b[177])^(a[348] & b[178])^(a[347] & b[179])^(a[346] & b[180])^(a[345] & b[181])^(a[344] & b[182])^(a[343] & b[183])^(a[342] & b[184])^(a[341] & b[185])^(a[340] & b[186])^(a[339] & b[187])^(a[338] & b[188])^(a[337] & b[189])^(a[336] & b[190])^(a[335] & b[191])^(a[334] & b[192])^(a[333] & b[193])^(a[332] & b[194])^(a[331] & b[195])^(a[330] & b[196])^(a[329] & b[197])^(a[328] & b[198])^(a[327] & b[199])^(a[326] & b[200])^(a[325] & b[201])^(a[324] & b[202])^(a[323] & b[203])^(a[322] & b[204])^(a[321] & b[205])^(a[320] & b[206])^(a[319] & b[207])^(a[318] & b[208])^(a[317] & b[209])^(a[316] & b[210])^(a[315] & b[211])^(a[314] & b[212])^(a[313] & b[213])^(a[312] & b[214])^(a[311] & b[215])^(a[310] & b[216])^(a[309] & b[217])^(a[308] & b[218])^(a[307] & b[219])^(a[306] & b[220])^(a[305] & b[221])^(a[304] & b[222])^(a[303] & b[223])^(a[302] & b[224])^(a[301] & b[225])^(a[300] & b[226])^(a[299] & b[227])^(a[298] & b[228])^(a[297] & b[229])^(a[296] & b[230])^(a[295] & b[231])^(a[294] & b[232])^(a[293] & b[233])^(a[292] & b[234])^(a[291] & b[235])^(a[290] & b[236])^(a[289] & b[237])^(a[288] & b[238])^(a[287] & b[239])^(a[286] & b[240])^(a[285] & b[241])^(a[284] & b[242])^(a[283] & b[243])^(a[282] & b[244])^(a[281] & b[245])^(a[280] & b[246])^(a[279] & b[247])^(a[278] & b[248])^(a[277] & b[249])^(a[276] & b[250])^(a[275] & b[251])^(a[274] & b[252])^(a[273] & b[253])^(a[272] & b[254])^(a[271] & b[255])^(a[270] & b[256])^(a[269] & b[257])^(a[268] & b[258])^(a[267] & b[259])^(a[266] & b[260])^(a[265] & b[261])^(a[264] & b[262])^(a[263] & b[263])^(a[262] & b[264])^(a[261] & b[265])^(a[260] & b[266])^(a[259] & b[267])^(a[258] & b[268])^(a[257] & b[269])^(a[256] & b[270])^(a[255] & b[271])^(a[254] & b[272])^(a[253] & b[273])^(a[252] & b[274])^(a[251] & b[275])^(a[250] & b[276])^(a[249] & b[277])^(a[248] & b[278])^(a[247] & b[279])^(a[246] & b[280])^(a[245] & b[281])^(a[244] & b[282])^(a[243] & b[283])^(a[242] & b[284])^(a[241] & b[285])^(a[240] & b[286])^(a[239] & b[287])^(a[238] & b[288])^(a[237] & b[289])^(a[236] & b[290])^(a[235] & b[291])^(a[234] & b[292])^(a[233] & b[293])^(a[232] & b[294])^(a[231] & b[295])^(a[230] & b[296])^(a[229] & b[297])^(a[228] & b[298])^(a[227] & b[299])^(a[226] & b[300])^(a[225] & b[301])^(a[224] & b[302])^(a[223] & b[303])^(a[222] & b[304])^(a[221] & b[305])^(a[220] & b[306])^(a[219] & b[307])^(a[218] & b[308])^(a[217] & b[309])^(a[216] & b[310])^(a[215] & b[311])^(a[214] & b[312])^(a[213] & b[313])^(a[212] & b[314])^(a[211] & b[315])^(a[210] & b[316])^(a[209] & b[317])^(a[208] & b[318])^(a[207] & b[319])^(a[206] & b[320])^(a[205] & b[321])^(a[204] & b[322])^(a[203] & b[323])^(a[202] & b[324])^(a[201] & b[325])^(a[200] & b[326])^(a[199] & b[327])^(a[198] & b[328])^(a[197] & b[329])^(a[196] & b[330])^(a[195] & b[331])^(a[194] & b[332])^(a[193] & b[333])^(a[192] & b[334])^(a[191] & b[335])^(a[190] & b[336])^(a[189] & b[337])^(a[188] & b[338])^(a[187] & b[339])^(a[186] & b[340])^(a[185] & b[341])^(a[184] & b[342])^(a[183] & b[343])^(a[182] & b[344])^(a[181] & b[345])^(a[180] & b[346])^(a[179] & b[347])^(a[178] & b[348])^(a[177] & b[349])^(a[176] & b[350])^(a[175] & b[351])^(a[174] & b[352])^(a[173] & b[353])^(a[172] & b[354])^(a[171] & b[355])^(a[170] & b[356])^(a[169] & b[357])^(a[168] & b[358])^(a[167] & b[359])^(a[166] & b[360])^(a[165] & b[361])^(a[164] & b[362])^(a[163] & b[363])^(a[162] & b[364])^(a[161] & b[365])^(a[160] & b[366])^(a[159] & b[367])^(a[158] & b[368])^(a[157] & b[369])^(a[156] & b[370])^(a[155] & b[371])^(a[154] & b[372])^(a[153] & b[373])^(a[152] & b[374])^(a[151] & b[375])^(a[150] & b[376])^(a[149] & b[377])^(a[148] & b[378])^(a[147] & b[379])^(a[146] & b[380])^(a[145] & b[381])^(a[144] & b[382])^(a[143] & b[383])^(a[142] & b[384])^(a[141] & b[385])^(a[140] & b[386])^(a[139] & b[387])^(a[138] & b[388])^(a[137] & b[389])^(a[136] & b[390])^(a[135] & b[391])^(a[134] & b[392])^(a[133] & b[393])^(a[132] & b[394])^(a[131] & b[395])^(a[130] & b[396])^(a[129] & b[397])^(a[128] & b[398])^(a[127] & b[399])^(a[126] & b[400])^(a[125] & b[401])^(a[124] & b[402])^(a[123] & b[403])^(a[122] & b[404])^(a[121] & b[405])^(a[120] & b[406])^(a[119] & b[407])^(a[118] & b[408]);
assign y[527] = (a[408] & b[119])^(a[407] & b[120])^(a[406] & b[121])^(a[405] & b[122])^(a[404] & b[123])^(a[403] & b[124])^(a[402] & b[125])^(a[401] & b[126])^(a[400] & b[127])^(a[399] & b[128])^(a[398] & b[129])^(a[397] & b[130])^(a[396] & b[131])^(a[395] & b[132])^(a[394] & b[133])^(a[393] & b[134])^(a[392] & b[135])^(a[391] & b[136])^(a[390] & b[137])^(a[389] & b[138])^(a[388] & b[139])^(a[387] & b[140])^(a[386] & b[141])^(a[385] & b[142])^(a[384] & b[143])^(a[383] & b[144])^(a[382] & b[145])^(a[381] & b[146])^(a[380] & b[147])^(a[379] & b[148])^(a[378] & b[149])^(a[377] & b[150])^(a[376] & b[151])^(a[375] & b[152])^(a[374] & b[153])^(a[373] & b[154])^(a[372] & b[155])^(a[371] & b[156])^(a[370] & b[157])^(a[369] & b[158])^(a[368] & b[159])^(a[367] & b[160])^(a[366] & b[161])^(a[365] & b[162])^(a[364] & b[163])^(a[363] & b[164])^(a[362] & b[165])^(a[361] & b[166])^(a[360] & b[167])^(a[359] & b[168])^(a[358] & b[169])^(a[357] & b[170])^(a[356] & b[171])^(a[355] & b[172])^(a[354] & b[173])^(a[353] & b[174])^(a[352] & b[175])^(a[351] & b[176])^(a[350] & b[177])^(a[349] & b[178])^(a[348] & b[179])^(a[347] & b[180])^(a[346] & b[181])^(a[345] & b[182])^(a[344] & b[183])^(a[343] & b[184])^(a[342] & b[185])^(a[341] & b[186])^(a[340] & b[187])^(a[339] & b[188])^(a[338] & b[189])^(a[337] & b[190])^(a[336] & b[191])^(a[335] & b[192])^(a[334] & b[193])^(a[333] & b[194])^(a[332] & b[195])^(a[331] & b[196])^(a[330] & b[197])^(a[329] & b[198])^(a[328] & b[199])^(a[327] & b[200])^(a[326] & b[201])^(a[325] & b[202])^(a[324] & b[203])^(a[323] & b[204])^(a[322] & b[205])^(a[321] & b[206])^(a[320] & b[207])^(a[319] & b[208])^(a[318] & b[209])^(a[317] & b[210])^(a[316] & b[211])^(a[315] & b[212])^(a[314] & b[213])^(a[313] & b[214])^(a[312] & b[215])^(a[311] & b[216])^(a[310] & b[217])^(a[309] & b[218])^(a[308] & b[219])^(a[307] & b[220])^(a[306] & b[221])^(a[305] & b[222])^(a[304] & b[223])^(a[303] & b[224])^(a[302] & b[225])^(a[301] & b[226])^(a[300] & b[227])^(a[299] & b[228])^(a[298] & b[229])^(a[297] & b[230])^(a[296] & b[231])^(a[295] & b[232])^(a[294] & b[233])^(a[293] & b[234])^(a[292] & b[235])^(a[291] & b[236])^(a[290] & b[237])^(a[289] & b[238])^(a[288] & b[239])^(a[287] & b[240])^(a[286] & b[241])^(a[285] & b[242])^(a[284] & b[243])^(a[283] & b[244])^(a[282] & b[245])^(a[281] & b[246])^(a[280] & b[247])^(a[279] & b[248])^(a[278] & b[249])^(a[277] & b[250])^(a[276] & b[251])^(a[275] & b[252])^(a[274] & b[253])^(a[273] & b[254])^(a[272] & b[255])^(a[271] & b[256])^(a[270] & b[257])^(a[269] & b[258])^(a[268] & b[259])^(a[267] & b[260])^(a[266] & b[261])^(a[265] & b[262])^(a[264] & b[263])^(a[263] & b[264])^(a[262] & b[265])^(a[261] & b[266])^(a[260] & b[267])^(a[259] & b[268])^(a[258] & b[269])^(a[257] & b[270])^(a[256] & b[271])^(a[255] & b[272])^(a[254] & b[273])^(a[253] & b[274])^(a[252] & b[275])^(a[251] & b[276])^(a[250] & b[277])^(a[249] & b[278])^(a[248] & b[279])^(a[247] & b[280])^(a[246] & b[281])^(a[245] & b[282])^(a[244] & b[283])^(a[243] & b[284])^(a[242] & b[285])^(a[241] & b[286])^(a[240] & b[287])^(a[239] & b[288])^(a[238] & b[289])^(a[237] & b[290])^(a[236] & b[291])^(a[235] & b[292])^(a[234] & b[293])^(a[233] & b[294])^(a[232] & b[295])^(a[231] & b[296])^(a[230] & b[297])^(a[229] & b[298])^(a[228] & b[299])^(a[227] & b[300])^(a[226] & b[301])^(a[225] & b[302])^(a[224] & b[303])^(a[223] & b[304])^(a[222] & b[305])^(a[221] & b[306])^(a[220] & b[307])^(a[219] & b[308])^(a[218] & b[309])^(a[217] & b[310])^(a[216] & b[311])^(a[215] & b[312])^(a[214] & b[313])^(a[213] & b[314])^(a[212] & b[315])^(a[211] & b[316])^(a[210] & b[317])^(a[209] & b[318])^(a[208] & b[319])^(a[207] & b[320])^(a[206] & b[321])^(a[205] & b[322])^(a[204] & b[323])^(a[203] & b[324])^(a[202] & b[325])^(a[201] & b[326])^(a[200] & b[327])^(a[199] & b[328])^(a[198] & b[329])^(a[197] & b[330])^(a[196] & b[331])^(a[195] & b[332])^(a[194] & b[333])^(a[193] & b[334])^(a[192] & b[335])^(a[191] & b[336])^(a[190] & b[337])^(a[189] & b[338])^(a[188] & b[339])^(a[187] & b[340])^(a[186] & b[341])^(a[185] & b[342])^(a[184] & b[343])^(a[183] & b[344])^(a[182] & b[345])^(a[181] & b[346])^(a[180] & b[347])^(a[179] & b[348])^(a[178] & b[349])^(a[177] & b[350])^(a[176] & b[351])^(a[175] & b[352])^(a[174] & b[353])^(a[173] & b[354])^(a[172] & b[355])^(a[171] & b[356])^(a[170] & b[357])^(a[169] & b[358])^(a[168] & b[359])^(a[167] & b[360])^(a[166] & b[361])^(a[165] & b[362])^(a[164] & b[363])^(a[163] & b[364])^(a[162] & b[365])^(a[161] & b[366])^(a[160] & b[367])^(a[159] & b[368])^(a[158] & b[369])^(a[157] & b[370])^(a[156] & b[371])^(a[155] & b[372])^(a[154] & b[373])^(a[153] & b[374])^(a[152] & b[375])^(a[151] & b[376])^(a[150] & b[377])^(a[149] & b[378])^(a[148] & b[379])^(a[147] & b[380])^(a[146] & b[381])^(a[145] & b[382])^(a[144] & b[383])^(a[143] & b[384])^(a[142] & b[385])^(a[141] & b[386])^(a[140] & b[387])^(a[139] & b[388])^(a[138] & b[389])^(a[137] & b[390])^(a[136] & b[391])^(a[135] & b[392])^(a[134] & b[393])^(a[133] & b[394])^(a[132] & b[395])^(a[131] & b[396])^(a[130] & b[397])^(a[129] & b[398])^(a[128] & b[399])^(a[127] & b[400])^(a[126] & b[401])^(a[125] & b[402])^(a[124] & b[403])^(a[123] & b[404])^(a[122] & b[405])^(a[121] & b[406])^(a[120] & b[407])^(a[119] & b[408]);
assign y[528] = (a[408] & b[120])^(a[407] & b[121])^(a[406] & b[122])^(a[405] & b[123])^(a[404] & b[124])^(a[403] & b[125])^(a[402] & b[126])^(a[401] & b[127])^(a[400] & b[128])^(a[399] & b[129])^(a[398] & b[130])^(a[397] & b[131])^(a[396] & b[132])^(a[395] & b[133])^(a[394] & b[134])^(a[393] & b[135])^(a[392] & b[136])^(a[391] & b[137])^(a[390] & b[138])^(a[389] & b[139])^(a[388] & b[140])^(a[387] & b[141])^(a[386] & b[142])^(a[385] & b[143])^(a[384] & b[144])^(a[383] & b[145])^(a[382] & b[146])^(a[381] & b[147])^(a[380] & b[148])^(a[379] & b[149])^(a[378] & b[150])^(a[377] & b[151])^(a[376] & b[152])^(a[375] & b[153])^(a[374] & b[154])^(a[373] & b[155])^(a[372] & b[156])^(a[371] & b[157])^(a[370] & b[158])^(a[369] & b[159])^(a[368] & b[160])^(a[367] & b[161])^(a[366] & b[162])^(a[365] & b[163])^(a[364] & b[164])^(a[363] & b[165])^(a[362] & b[166])^(a[361] & b[167])^(a[360] & b[168])^(a[359] & b[169])^(a[358] & b[170])^(a[357] & b[171])^(a[356] & b[172])^(a[355] & b[173])^(a[354] & b[174])^(a[353] & b[175])^(a[352] & b[176])^(a[351] & b[177])^(a[350] & b[178])^(a[349] & b[179])^(a[348] & b[180])^(a[347] & b[181])^(a[346] & b[182])^(a[345] & b[183])^(a[344] & b[184])^(a[343] & b[185])^(a[342] & b[186])^(a[341] & b[187])^(a[340] & b[188])^(a[339] & b[189])^(a[338] & b[190])^(a[337] & b[191])^(a[336] & b[192])^(a[335] & b[193])^(a[334] & b[194])^(a[333] & b[195])^(a[332] & b[196])^(a[331] & b[197])^(a[330] & b[198])^(a[329] & b[199])^(a[328] & b[200])^(a[327] & b[201])^(a[326] & b[202])^(a[325] & b[203])^(a[324] & b[204])^(a[323] & b[205])^(a[322] & b[206])^(a[321] & b[207])^(a[320] & b[208])^(a[319] & b[209])^(a[318] & b[210])^(a[317] & b[211])^(a[316] & b[212])^(a[315] & b[213])^(a[314] & b[214])^(a[313] & b[215])^(a[312] & b[216])^(a[311] & b[217])^(a[310] & b[218])^(a[309] & b[219])^(a[308] & b[220])^(a[307] & b[221])^(a[306] & b[222])^(a[305] & b[223])^(a[304] & b[224])^(a[303] & b[225])^(a[302] & b[226])^(a[301] & b[227])^(a[300] & b[228])^(a[299] & b[229])^(a[298] & b[230])^(a[297] & b[231])^(a[296] & b[232])^(a[295] & b[233])^(a[294] & b[234])^(a[293] & b[235])^(a[292] & b[236])^(a[291] & b[237])^(a[290] & b[238])^(a[289] & b[239])^(a[288] & b[240])^(a[287] & b[241])^(a[286] & b[242])^(a[285] & b[243])^(a[284] & b[244])^(a[283] & b[245])^(a[282] & b[246])^(a[281] & b[247])^(a[280] & b[248])^(a[279] & b[249])^(a[278] & b[250])^(a[277] & b[251])^(a[276] & b[252])^(a[275] & b[253])^(a[274] & b[254])^(a[273] & b[255])^(a[272] & b[256])^(a[271] & b[257])^(a[270] & b[258])^(a[269] & b[259])^(a[268] & b[260])^(a[267] & b[261])^(a[266] & b[262])^(a[265] & b[263])^(a[264] & b[264])^(a[263] & b[265])^(a[262] & b[266])^(a[261] & b[267])^(a[260] & b[268])^(a[259] & b[269])^(a[258] & b[270])^(a[257] & b[271])^(a[256] & b[272])^(a[255] & b[273])^(a[254] & b[274])^(a[253] & b[275])^(a[252] & b[276])^(a[251] & b[277])^(a[250] & b[278])^(a[249] & b[279])^(a[248] & b[280])^(a[247] & b[281])^(a[246] & b[282])^(a[245] & b[283])^(a[244] & b[284])^(a[243] & b[285])^(a[242] & b[286])^(a[241] & b[287])^(a[240] & b[288])^(a[239] & b[289])^(a[238] & b[290])^(a[237] & b[291])^(a[236] & b[292])^(a[235] & b[293])^(a[234] & b[294])^(a[233] & b[295])^(a[232] & b[296])^(a[231] & b[297])^(a[230] & b[298])^(a[229] & b[299])^(a[228] & b[300])^(a[227] & b[301])^(a[226] & b[302])^(a[225] & b[303])^(a[224] & b[304])^(a[223] & b[305])^(a[222] & b[306])^(a[221] & b[307])^(a[220] & b[308])^(a[219] & b[309])^(a[218] & b[310])^(a[217] & b[311])^(a[216] & b[312])^(a[215] & b[313])^(a[214] & b[314])^(a[213] & b[315])^(a[212] & b[316])^(a[211] & b[317])^(a[210] & b[318])^(a[209] & b[319])^(a[208] & b[320])^(a[207] & b[321])^(a[206] & b[322])^(a[205] & b[323])^(a[204] & b[324])^(a[203] & b[325])^(a[202] & b[326])^(a[201] & b[327])^(a[200] & b[328])^(a[199] & b[329])^(a[198] & b[330])^(a[197] & b[331])^(a[196] & b[332])^(a[195] & b[333])^(a[194] & b[334])^(a[193] & b[335])^(a[192] & b[336])^(a[191] & b[337])^(a[190] & b[338])^(a[189] & b[339])^(a[188] & b[340])^(a[187] & b[341])^(a[186] & b[342])^(a[185] & b[343])^(a[184] & b[344])^(a[183] & b[345])^(a[182] & b[346])^(a[181] & b[347])^(a[180] & b[348])^(a[179] & b[349])^(a[178] & b[350])^(a[177] & b[351])^(a[176] & b[352])^(a[175] & b[353])^(a[174] & b[354])^(a[173] & b[355])^(a[172] & b[356])^(a[171] & b[357])^(a[170] & b[358])^(a[169] & b[359])^(a[168] & b[360])^(a[167] & b[361])^(a[166] & b[362])^(a[165] & b[363])^(a[164] & b[364])^(a[163] & b[365])^(a[162] & b[366])^(a[161] & b[367])^(a[160] & b[368])^(a[159] & b[369])^(a[158] & b[370])^(a[157] & b[371])^(a[156] & b[372])^(a[155] & b[373])^(a[154] & b[374])^(a[153] & b[375])^(a[152] & b[376])^(a[151] & b[377])^(a[150] & b[378])^(a[149] & b[379])^(a[148] & b[380])^(a[147] & b[381])^(a[146] & b[382])^(a[145] & b[383])^(a[144] & b[384])^(a[143] & b[385])^(a[142] & b[386])^(a[141] & b[387])^(a[140] & b[388])^(a[139] & b[389])^(a[138] & b[390])^(a[137] & b[391])^(a[136] & b[392])^(a[135] & b[393])^(a[134] & b[394])^(a[133] & b[395])^(a[132] & b[396])^(a[131] & b[397])^(a[130] & b[398])^(a[129] & b[399])^(a[128] & b[400])^(a[127] & b[401])^(a[126] & b[402])^(a[125] & b[403])^(a[124] & b[404])^(a[123] & b[405])^(a[122] & b[406])^(a[121] & b[407])^(a[120] & b[408]);
assign y[529] = (a[408] & b[121])^(a[407] & b[122])^(a[406] & b[123])^(a[405] & b[124])^(a[404] & b[125])^(a[403] & b[126])^(a[402] & b[127])^(a[401] & b[128])^(a[400] & b[129])^(a[399] & b[130])^(a[398] & b[131])^(a[397] & b[132])^(a[396] & b[133])^(a[395] & b[134])^(a[394] & b[135])^(a[393] & b[136])^(a[392] & b[137])^(a[391] & b[138])^(a[390] & b[139])^(a[389] & b[140])^(a[388] & b[141])^(a[387] & b[142])^(a[386] & b[143])^(a[385] & b[144])^(a[384] & b[145])^(a[383] & b[146])^(a[382] & b[147])^(a[381] & b[148])^(a[380] & b[149])^(a[379] & b[150])^(a[378] & b[151])^(a[377] & b[152])^(a[376] & b[153])^(a[375] & b[154])^(a[374] & b[155])^(a[373] & b[156])^(a[372] & b[157])^(a[371] & b[158])^(a[370] & b[159])^(a[369] & b[160])^(a[368] & b[161])^(a[367] & b[162])^(a[366] & b[163])^(a[365] & b[164])^(a[364] & b[165])^(a[363] & b[166])^(a[362] & b[167])^(a[361] & b[168])^(a[360] & b[169])^(a[359] & b[170])^(a[358] & b[171])^(a[357] & b[172])^(a[356] & b[173])^(a[355] & b[174])^(a[354] & b[175])^(a[353] & b[176])^(a[352] & b[177])^(a[351] & b[178])^(a[350] & b[179])^(a[349] & b[180])^(a[348] & b[181])^(a[347] & b[182])^(a[346] & b[183])^(a[345] & b[184])^(a[344] & b[185])^(a[343] & b[186])^(a[342] & b[187])^(a[341] & b[188])^(a[340] & b[189])^(a[339] & b[190])^(a[338] & b[191])^(a[337] & b[192])^(a[336] & b[193])^(a[335] & b[194])^(a[334] & b[195])^(a[333] & b[196])^(a[332] & b[197])^(a[331] & b[198])^(a[330] & b[199])^(a[329] & b[200])^(a[328] & b[201])^(a[327] & b[202])^(a[326] & b[203])^(a[325] & b[204])^(a[324] & b[205])^(a[323] & b[206])^(a[322] & b[207])^(a[321] & b[208])^(a[320] & b[209])^(a[319] & b[210])^(a[318] & b[211])^(a[317] & b[212])^(a[316] & b[213])^(a[315] & b[214])^(a[314] & b[215])^(a[313] & b[216])^(a[312] & b[217])^(a[311] & b[218])^(a[310] & b[219])^(a[309] & b[220])^(a[308] & b[221])^(a[307] & b[222])^(a[306] & b[223])^(a[305] & b[224])^(a[304] & b[225])^(a[303] & b[226])^(a[302] & b[227])^(a[301] & b[228])^(a[300] & b[229])^(a[299] & b[230])^(a[298] & b[231])^(a[297] & b[232])^(a[296] & b[233])^(a[295] & b[234])^(a[294] & b[235])^(a[293] & b[236])^(a[292] & b[237])^(a[291] & b[238])^(a[290] & b[239])^(a[289] & b[240])^(a[288] & b[241])^(a[287] & b[242])^(a[286] & b[243])^(a[285] & b[244])^(a[284] & b[245])^(a[283] & b[246])^(a[282] & b[247])^(a[281] & b[248])^(a[280] & b[249])^(a[279] & b[250])^(a[278] & b[251])^(a[277] & b[252])^(a[276] & b[253])^(a[275] & b[254])^(a[274] & b[255])^(a[273] & b[256])^(a[272] & b[257])^(a[271] & b[258])^(a[270] & b[259])^(a[269] & b[260])^(a[268] & b[261])^(a[267] & b[262])^(a[266] & b[263])^(a[265] & b[264])^(a[264] & b[265])^(a[263] & b[266])^(a[262] & b[267])^(a[261] & b[268])^(a[260] & b[269])^(a[259] & b[270])^(a[258] & b[271])^(a[257] & b[272])^(a[256] & b[273])^(a[255] & b[274])^(a[254] & b[275])^(a[253] & b[276])^(a[252] & b[277])^(a[251] & b[278])^(a[250] & b[279])^(a[249] & b[280])^(a[248] & b[281])^(a[247] & b[282])^(a[246] & b[283])^(a[245] & b[284])^(a[244] & b[285])^(a[243] & b[286])^(a[242] & b[287])^(a[241] & b[288])^(a[240] & b[289])^(a[239] & b[290])^(a[238] & b[291])^(a[237] & b[292])^(a[236] & b[293])^(a[235] & b[294])^(a[234] & b[295])^(a[233] & b[296])^(a[232] & b[297])^(a[231] & b[298])^(a[230] & b[299])^(a[229] & b[300])^(a[228] & b[301])^(a[227] & b[302])^(a[226] & b[303])^(a[225] & b[304])^(a[224] & b[305])^(a[223] & b[306])^(a[222] & b[307])^(a[221] & b[308])^(a[220] & b[309])^(a[219] & b[310])^(a[218] & b[311])^(a[217] & b[312])^(a[216] & b[313])^(a[215] & b[314])^(a[214] & b[315])^(a[213] & b[316])^(a[212] & b[317])^(a[211] & b[318])^(a[210] & b[319])^(a[209] & b[320])^(a[208] & b[321])^(a[207] & b[322])^(a[206] & b[323])^(a[205] & b[324])^(a[204] & b[325])^(a[203] & b[326])^(a[202] & b[327])^(a[201] & b[328])^(a[200] & b[329])^(a[199] & b[330])^(a[198] & b[331])^(a[197] & b[332])^(a[196] & b[333])^(a[195] & b[334])^(a[194] & b[335])^(a[193] & b[336])^(a[192] & b[337])^(a[191] & b[338])^(a[190] & b[339])^(a[189] & b[340])^(a[188] & b[341])^(a[187] & b[342])^(a[186] & b[343])^(a[185] & b[344])^(a[184] & b[345])^(a[183] & b[346])^(a[182] & b[347])^(a[181] & b[348])^(a[180] & b[349])^(a[179] & b[350])^(a[178] & b[351])^(a[177] & b[352])^(a[176] & b[353])^(a[175] & b[354])^(a[174] & b[355])^(a[173] & b[356])^(a[172] & b[357])^(a[171] & b[358])^(a[170] & b[359])^(a[169] & b[360])^(a[168] & b[361])^(a[167] & b[362])^(a[166] & b[363])^(a[165] & b[364])^(a[164] & b[365])^(a[163] & b[366])^(a[162] & b[367])^(a[161] & b[368])^(a[160] & b[369])^(a[159] & b[370])^(a[158] & b[371])^(a[157] & b[372])^(a[156] & b[373])^(a[155] & b[374])^(a[154] & b[375])^(a[153] & b[376])^(a[152] & b[377])^(a[151] & b[378])^(a[150] & b[379])^(a[149] & b[380])^(a[148] & b[381])^(a[147] & b[382])^(a[146] & b[383])^(a[145] & b[384])^(a[144] & b[385])^(a[143] & b[386])^(a[142] & b[387])^(a[141] & b[388])^(a[140] & b[389])^(a[139] & b[390])^(a[138] & b[391])^(a[137] & b[392])^(a[136] & b[393])^(a[135] & b[394])^(a[134] & b[395])^(a[133] & b[396])^(a[132] & b[397])^(a[131] & b[398])^(a[130] & b[399])^(a[129] & b[400])^(a[128] & b[401])^(a[127] & b[402])^(a[126] & b[403])^(a[125] & b[404])^(a[124] & b[405])^(a[123] & b[406])^(a[122] & b[407])^(a[121] & b[408]);
assign y[530] = (a[408] & b[122])^(a[407] & b[123])^(a[406] & b[124])^(a[405] & b[125])^(a[404] & b[126])^(a[403] & b[127])^(a[402] & b[128])^(a[401] & b[129])^(a[400] & b[130])^(a[399] & b[131])^(a[398] & b[132])^(a[397] & b[133])^(a[396] & b[134])^(a[395] & b[135])^(a[394] & b[136])^(a[393] & b[137])^(a[392] & b[138])^(a[391] & b[139])^(a[390] & b[140])^(a[389] & b[141])^(a[388] & b[142])^(a[387] & b[143])^(a[386] & b[144])^(a[385] & b[145])^(a[384] & b[146])^(a[383] & b[147])^(a[382] & b[148])^(a[381] & b[149])^(a[380] & b[150])^(a[379] & b[151])^(a[378] & b[152])^(a[377] & b[153])^(a[376] & b[154])^(a[375] & b[155])^(a[374] & b[156])^(a[373] & b[157])^(a[372] & b[158])^(a[371] & b[159])^(a[370] & b[160])^(a[369] & b[161])^(a[368] & b[162])^(a[367] & b[163])^(a[366] & b[164])^(a[365] & b[165])^(a[364] & b[166])^(a[363] & b[167])^(a[362] & b[168])^(a[361] & b[169])^(a[360] & b[170])^(a[359] & b[171])^(a[358] & b[172])^(a[357] & b[173])^(a[356] & b[174])^(a[355] & b[175])^(a[354] & b[176])^(a[353] & b[177])^(a[352] & b[178])^(a[351] & b[179])^(a[350] & b[180])^(a[349] & b[181])^(a[348] & b[182])^(a[347] & b[183])^(a[346] & b[184])^(a[345] & b[185])^(a[344] & b[186])^(a[343] & b[187])^(a[342] & b[188])^(a[341] & b[189])^(a[340] & b[190])^(a[339] & b[191])^(a[338] & b[192])^(a[337] & b[193])^(a[336] & b[194])^(a[335] & b[195])^(a[334] & b[196])^(a[333] & b[197])^(a[332] & b[198])^(a[331] & b[199])^(a[330] & b[200])^(a[329] & b[201])^(a[328] & b[202])^(a[327] & b[203])^(a[326] & b[204])^(a[325] & b[205])^(a[324] & b[206])^(a[323] & b[207])^(a[322] & b[208])^(a[321] & b[209])^(a[320] & b[210])^(a[319] & b[211])^(a[318] & b[212])^(a[317] & b[213])^(a[316] & b[214])^(a[315] & b[215])^(a[314] & b[216])^(a[313] & b[217])^(a[312] & b[218])^(a[311] & b[219])^(a[310] & b[220])^(a[309] & b[221])^(a[308] & b[222])^(a[307] & b[223])^(a[306] & b[224])^(a[305] & b[225])^(a[304] & b[226])^(a[303] & b[227])^(a[302] & b[228])^(a[301] & b[229])^(a[300] & b[230])^(a[299] & b[231])^(a[298] & b[232])^(a[297] & b[233])^(a[296] & b[234])^(a[295] & b[235])^(a[294] & b[236])^(a[293] & b[237])^(a[292] & b[238])^(a[291] & b[239])^(a[290] & b[240])^(a[289] & b[241])^(a[288] & b[242])^(a[287] & b[243])^(a[286] & b[244])^(a[285] & b[245])^(a[284] & b[246])^(a[283] & b[247])^(a[282] & b[248])^(a[281] & b[249])^(a[280] & b[250])^(a[279] & b[251])^(a[278] & b[252])^(a[277] & b[253])^(a[276] & b[254])^(a[275] & b[255])^(a[274] & b[256])^(a[273] & b[257])^(a[272] & b[258])^(a[271] & b[259])^(a[270] & b[260])^(a[269] & b[261])^(a[268] & b[262])^(a[267] & b[263])^(a[266] & b[264])^(a[265] & b[265])^(a[264] & b[266])^(a[263] & b[267])^(a[262] & b[268])^(a[261] & b[269])^(a[260] & b[270])^(a[259] & b[271])^(a[258] & b[272])^(a[257] & b[273])^(a[256] & b[274])^(a[255] & b[275])^(a[254] & b[276])^(a[253] & b[277])^(a[252] & b[278])^(a[251] & b[279])^(a[250] & b[280])^(a[249] & b[281])^(a[248] & b[282])^(a[247] & b[283])^(a[246] & b[284])^(a[245] & b[285])^(a[244] & b[286])^(a[243] & b[287])^(a[242] & b[288])^(a[241] & b[289])^(a[240] & b[290])^(a[239] & b[291])^(a[238] & b[292])^(a[237] & b[293])^(a[236] & b[294])^(a[235] & b[295])^(a[234] & b[296])^(a[233] & b[297])^(a[232] & b[298])^(a[231] & b[299])^(a[230] & b[300])^(a[229] & b[301])^(a[228] & b[302])^(a[227] & b[303])^(a[226] & b[304])^(a[225] & b[305])^(a[224] & b[306])^(a[223] & b[307])^(a[222] & b[308])^(a[221] & b[309])^(a[220] & b[310])^(a[219] & b[311])^(a[218] & b[312])^(a[217] & b[313])^(a[216] & b[314])^(a[215] & b[315])^(a[214] & b[316])^(a[213] & b[317])^(a[212] & b[318])^(a[211] & b[319])^(a[210] & b[320])^(a[209] & b[321])^(a[208] & b[322])^(a[207] & b[323])^(a[206] & b[324])^(a[205] & b[325])^(a[204] & b[326])^(a[203] & b[327])^(a[202] & b[328])^(a[201] & b[329])^(a[200] & b[330])^(a[199] & b[331])^(a[198] & b[332])^(a[197] & b[333])^(a[196] & b[334])^(a[195] & b[335])^(a[194] & b[336])^(a[193] & b[337])^(a[192] & b[338])^(a[191] & b[339])^(a[190] & b[340])^(a[189] & b[341])^(a[188] & b[342])^(a[187] & b[343])^(a[186] & b[344])^(a[185] & b[345])^(a[184] & b[346])^(a[183] & b[347])^(a[182] & b[348])^(a[181] & b[349])^(a[180] & b[350])^(a[179] & b[351])^(a[178] & b[352])^(a[177] & b[353])^(a[176] & b[354])^(a[175] & b[355])^(a[174] & b[356])^(a[173] & b[357])^(a[172] & b[358])^(a[171] & b[359])^(a[170] & b[360])^(a[169] & b[361])^(a[168] & b[362])^(a[167] & b[363])^(a[166] & b[364])^(a[165] & b[365])^(a[164] & b[366])^(a[163] & b[367])^(a[162] & b[368])^(a[161] & b[369])^(a[160] & b[370])^(a[159] & b[371])^(a[158] & b[372])^(a[157] & b[373])^(a[156] & b[374])^(a[155] & b[375])^(a[154] & b[376])^(a[153] & b[377])^(a[152] & b[378])^(a[151] & b[379])^(a[150] & b[380])^(a[149] & b[381])^(a[148] & b[382])^(a[147] & b[383])^(a[146] & b[384])^(a[145] & b[385])^(a[144] & b[386])^(a[143] & b[387])^(a[142] & b[388])^(a[141] & b[389])^(a[140] & b[390])^(a[139] & b[391])^(a[138] & b[392])^(a[137] & b[393])^(a[136] & b[394])^(a[135] & b[395])^(a[134] & b[396])^(a[133] & b[397])^(a[132] & b[398])^(a[131] & b[399])^(a[130] & b[400])^(a[129] & b[401])^(a[128] & b[402])^(a[127] & b[403])^(a[126] & b[404])^(a[125] & b[405])^(a[124] & b[406])^(a[123] & b[407])^(a[122] & b[408]);
assign y[531] = (a[408] & b[123])^(a[407] & b[124])^(a[406] & b[125])^(a[405] & b[126])^(a[404] & b[127])^(a[403] & b[128])^(a[402] & b[129])^(a[401] & b[130])^(a[400] & b[131])^(a[399] & b[132])^(a[398] & b[133])^(a[397] & b[134])^(a[396] & b[135])^(a[395] & b[136])^(a[394] & b[137])^(a[393] & b[138])^(a[392] & b[139])^(a[391] & b[140])^(a[390] & b[141])^(a[389] & b[142])^(a[388] & b[143])^(a[387] & b[144])^(a[386] & b[145])^(a[385] & b[146])^(a[384] & b[147])^(a[383] & b[148])^(a[382] & b[149])^(a[381] & b[150])^(a[380] & b[151])^(a[379] & b[152])^(a[378] & b[153])^(a[377] & b[154])^(a[376] & b[155])^(a[375] & b[156])^(a[374] & b[157])^(a[373] & b[158])^(a[372] & b[159])^(a[371] & b[160])^(a[370] & b[161])^(a[369] & b[162])^(a[368] & b[163])^(a[367] & b[164])^(a[366] & b[165])^(a[365] & b[166])^(a[364] & b[167])^(a[363] & b[168])^(a[362] & b[169])^(a[361] & b[170])^(a[360] & b[171])^(a[359] & b[172])^(a[358] & b[173])^(a[357] & b[174])^(a[356] & b[175])^(a[355] & b[176])^(a[354] & b[177])^(a[353] & b[178])^(a[352] & b[179])^(a[351] & b[180])^(a[350] & b[181])^(a[349] & b[182])^(a[348] & b[183])^(a[347] & b[184])^(a[346] & b[185])^(a[345] & b[186])^(a[344] & b[187])^(a[343] & b[188])^(a[342] & b[189])^(a[341] & b[190])^(a[340] & b[191])^(a[339] & b[192])^(a[338] & b[193])^(a[337] & b[194])^(a[336] & b[195])^(a[335] & b[196])^(a[334] & b[197])^(a[333] & b[198])^(a[332] & b[199])^(a[331] & b[200])^(a[330] & b[201])^(a[329] & b[202])^(a[328] & b[203])^(a[327] & b[204])^(a[326] & b[205])^(a[325] & b[206])^(a[324] & b[207])^(a[323] & b[208])^(a[322] & b[209])^(a[321] & b[210])^(a[320] & b[211])^(a[319] & b[212])^(a[318] & b[213])^(a[317] & b[214])^(a[316] & b[215])^(a[315] & b[216])^(a[314] & b[217])^(a[313] & b[218])^(a[312] & b[219])^(a[311] & b[220])^(a[310] & b[221])^(a[309] & b[222])^(a[308] & b[223])^(a[307] & b[224])^(a[306] & b[225])^(a[305] & b[226])^(a[304] & b[227])^(a[303] & b[228])^(a[302] & b[229])^(a[301] & b[230])^(a[300] & b[231])^(a[299] & b[232])^(a[298] & b[233])^(a[297] & b[234])^(a[296] & b[235])^(a[295] & b[236])^(a[294] & b[237])^(a[293] & b[238])^(a[292] & b[239])^(a[291] & b[240])^(a[290] & b[241])^(a[289] & b[242])^(a[288] & b[243])^(a[287] & b[244])^(a[286] & b[245])^(a[285] & b[246])^(a[284] & b[247])^(a[283] & b[248])^(a[282] & b[249])^(a[281] & b[250])^(a[280] & b[251])^(a[279] & b[252])^(a[278] & b[253])^(a[277] & b[254])^(a[276] & b[255])^(a[275] & b[256])^(a[274] & b[257])^(a[273] & b[258])^(a[272] & b[259])^(a[271] & b[260])^(a[270] & b[261])^(a[269] & b[262])^(a[268] & b[263])^(a[267] & b[264])^(a[266] & b[265])^(a[265] & b[266])^(a[264] & b[267])^(a[263] & b[268])^(a[262] & b[269])^(a[261] & b[270])^(a[260] & b[271])^(a[259] & b[272])^(a[258] & b[273])^(a[257] & b[274])^(a[256] & b[275])^(a[255] & b[276])^(a[254] & b[277])^(a[253] & b[278])^(a[252] & b[279])^(a[251] & b[280])^(a[250] & b[281])^(a[249] & b[282])^(a[248] & b[283])^(a[247] & b[284])^(a[246] & b[285])^(a[245] & b[286])^(a[244] & b[287])^(a[243] & b[288])^(a[242] & b[289])^(a[241] & b[290])^(a[240] & b[291])^(a[239] & b[292])^(a[238] & b[293])^(a[237] & b[294])^(a[236] & b[295])^(a[235] & b[296])^(a[234] & b[297])^(a[233] & b[298])^(a[232] & b[299])^(a[231] & b[300])^(a[230] & b[301])^(a[229] & b[302])^(a[228] & b[303])^(a[227] & b[304])^(a[226] & b[305])^(a[225] & b[306])^(a[224] & b[307])^(a[223] & b[308])^(a[222] & b[309])^(a[221] & b[310])^(a[220] & b[311])^(a[219] & b[312])^(a[218] & b[313])^(a[217] & b[314])^(a[216] & b[315])^(a[215] & b[316])^(a[214] & b[317])^(a[213] & b[318])^(a[212] & b[319])^(a[211] & b[320])^(a[210] & b[321])^(a[209] & b[322])^(a[208] & b[323])^(a[207] & b[324])^(a[206] & b[325])^(a[205] & b[326])^(a[204] & b[327])^(a[203] & b[328])^(a[202] & b[329])^(a[201] & b[330])^(a[200] & b[331])^(a[199] & b[332])^(a[198] & b[333])^(a[197] & b[334])^(a[196] & b[335])^(a[195] & b[336])^(a[194] & b[337])^(a[193] & b[338])^(a[192] & b[339])^(a[191] & b[340])^(a[190] & b[341])^(a[189] & b[342])^(a[188] & b[343])^(a[187] & b[344])^(a[186] & b[345])^(a[185] & b[346])^(a[184] & b[347])^(a[183] & b[348])^(a[182] & b[349])^(a[181] & b[350])^(a[180] & b[351])^(a[179] & b[352])^(a[178] & b[353])^(a[177] & b[354])^(a[176] & b[355])^(a[175] & b[356])^(a[174] & b[357])^(a[173] & b[358])^(a[172] & b[359])^(a[171] & b[360])^(a[170] & b[361])^(a[169] & b[362])^(a[168] & b[363])^(a[167] & b[364])^(a[166] & b[365])^(a[165] & b[366])^(a[164] & b[367])^(a[163] & b[368])^(a[162] & b[369])^(a[161] & b[370])^(a[160] & b[371])^(a[159] & b[372])^(a[158] & b[373])^(a[157] & b[374])^(a[156] & b[375])^(a[155] & b[376])^(a[154] & b[377])^(a[153] & b[378])^(a[152] & b[379])^(a[151] & b[380])^(a[150] & b[381])^(a[149] & b[382])^(a[148] & b[383])^(a[147] & b[384])^(a[146] & b[385])^(a[145] & b[386])^(a[144] & b[387])^(a[143] & b[388])^(a[142] & b[389])^(a[141] & b[390])^(a[140] & b[391])^(a[139] & b[392])^(a[138] & b[393])^(a[137] & b[394])^(a[136] & b[395])^(a[135] & b[396])^(a[134] & b[397])^(a[133] & b[398])^(a[132] & b[399])^(a[131] & b[400])^(a[130] & b[401])^(a[129] & b[402])^(a[128] & b[403])^(a[127] & b[404])^(a[126] & b[405])^(a[125] & b[406])^(a[124] & b[407])^(a[123] & b[408]);
assign y[532] = (a[408] & b[124])^(a[407] & b[125])^(a[406] & b[126])^(a[405] & b[127])^(a[404] & b[128])^(a[403] & b[129])^(a[402] & b[130])^(a[401] & b[131])^(a[400] & b[132])^(a[399] & b[133])^(a[398] & b[134])^(a[397] & b[135])^(a[396] & b[136])^(a[395] & b[137])^(a[394] & b[138])^(a[393] & b[139])^(a[392] & b[140])^(a[391] & b[141])^(a[390] & b[142])^(a[389] & b[143])^(a[388] & b[144])^(a[387] & b[145])^(a[386] & b[146])^(a[385] & b[147])^(a[384] & b[148])^(a[383] & b[149])^(a[382] & b[150])^(a[381] & b[151])^(a[380] & b[152])^(a[379] & b[153])^(a[378] & b[154])^(a[377] & b[155])^(a[376] & b[156])^(a[375] & b[157])^(a[374] & b[158])^(a[373] & b[159])^(a[372] & b[160])^(a[371] & b[161])^(a[370] & b[162])^(a[369] & b[163])^(a[368] & b[164])^(a[367] & b[165])^(a[366] & b[166])^(a[365] & b[167])^(a[364] & b[168])^(a[363] & b[169])^(a[362] & b[170])^(a[361] & b[171])^(a[360] & b[172])^(a[359] & b[173])^(a[358] & b[174])^(a[357] & b[175])^(a[356] & b[176])^(a[355] & b[177])^(a[354] & b[178])^(a[353] & b[179])^(a[352] & b[180])^(a[351] & b[181])^(a[350] & b[182])^(a[349] & b[183])^(a[348] & b[184])^(a[347] & b[185])^(a[346] & b[186])^(a[345] & b[187])^(a[344] & b[188])^(a[343] & b[189])^(a[342] & b[190])^(a[341] & b[191])^(a[340] & b[192])^(a[339] & b[193])^(a[338] & b[194])^(a[337] & b[195])^(a[336] & b[196])^(a[335] & b[197])^(a[334] & b[198])^(a[333] & b[199])^(a[332] & b[200])^(a[331] & b[201])^(a[330] & b[202])^(a[329] & b[203])^(a[328] & b[204])^(a[327] & b[205])^(a[326] & b[206])^(a[325] & b[207])^(a[324] & b[208])^(a[323] & b[209])^(a[322] & b[210])^(a[321] & b[211])^(a[320] & b[212])^(a[319] & b[213])^(a[318] & b[214])^(a[317] & b[215])^(a[316] & b[216])^(a[315] & b[217])^(a[314] & b[218])^(a[313] & b[219])^(a[312] & b[220])^(a[311] & b[221])^(a[310] & b[222])^(a[309] & b[223])^(a[308] & b[224])^(a[307] & b[225])^(a[306] & b[226])^(a[305] & b[227])^(a[304] & b[228])^(a[303] & b[229])^(a[302] & b[230])^(a[301] & b[231])^(a[300] & b[232])^(a[299] & b[233])^(a[298] & b[234])^(a[297] & b[235])^(a[296] & b[236])^(a[295] & b[237])^(a[294] & b[238])^(a[293] & b[239])^(a[292] & b[240])^(a[291] & b[241])^(a[290] & b[242])^(a[289] & b[243])^(a[288] & b[244])^(a[287] & b[245])^(a[286] & b[246])^(a[285] & b[247])^(a[284] & b[248])^(a[283] & b[249])^(a[282] & b[250])^(a[281] & b[251])^(a[280] & b[252])^(a[279] & b[253])^(a[278] & b[254])^(a[277] & b[255])^(a[276] & b[256])^(a[275] & b[257])^(a[274] & b[258])^(a[273] & b[259])^(a[272] & b[260])^(a[271] & b[261])^(a[270] & b[262])^(a[269] & b[263])^(a[268] & b[264])^(a[267] & b[265])^(a[266] & b[266])^(a[265] & b[267])^(a[264] & b[268])^(a[263] & b[269])^(a[262] & b[270])^(a[261] & b[271])^(a[260] & b[272])^(a[259] & b[273])^(a[258] & b[274])^(a[257] & b[275])^(a[256] & b[276])^(a[255] & b[277])^(a[254] & b[278])^(a[253] & b[279])^(a[252] & b[280])^(a[251] & b[281])^(a[250] & b[282])^(a[249] & b[283])^(a[248] & b[284])^(a[247] & b[285])^(a[246] & b[286])^(a[245] & b[287])^(a[244] & b[288])^(a[243] & b[289])^(a[242] & b[290])^(a[241] & b[291])^(a[240] & b[292])^(a[239] & b[293])^(a[238] & b[294])^(a[237] & b[295])^(a[236] & b[296])^(a[235] & b[297])^(a[234] & b[298])^(a[233] & b[299])^(a[232] & b[300])^(a[231] & b[301])^(a[230] & b[302])^(a[229] & b[303])^(a[228] & b[304])^(a[227] & b[305])^(a[226] & b[306])^(a[225] & b[307])^(a[224] & b[308])^(a[223] & b[309])^(a[222] & b[310])^(a[221] & b[311])^(a[220] & b[312])^(a[219] & b[313])^(a[218] & b[314])^(a[217] & b[315])^(a[216] & b[316])^(a[215] & b[317])^(a[214] & b[318])^(a[213] & b[319])^(a[212] & b[320])^(a[211] & b[321])^(a[210] & b[322])^(a[209] & b[323])^(a[208] & b[324])^(a[207] & b[325])^(a[206] & b[326])^(a[205] & b[327])^(a[204] & b[328])^(a[203] & b[329])^(a[202] & b[330])^(a[201] & b[331])^(a[200] & b[332])^(a[199] & b[333])^(a[198] & b[334])^(a[197] & b[335])^(a[196] & b[336])^(a[195] & b[337])^(a[194] & b[338])^(a[193] & b[339])^(a[192] & b[340])^(a[191] & b[341])^(a[190] & b[342])^(a[189] & b[343])^(a[188] & b[344])^(a[187] & b[345])^(a[186] & b[346])^(a[185] & b[347])^(a[184] & b[348])^(a[183] & b[349])^(a[182] & b[350])^(a[181] & b[351])^(a[180] & b[352])^(a[179] & b[353])^(a[178] & b[354])^(a[177] & b[355])^(a[176] & b[356])^(a[175] & b[357])^(a[174] & b[358])^(a[173] & b[359])^(a[172] & b[360])^(a[171] & b[361])^(a[170] & b[362])^(a[169] & b[363])^(a[168] & b[364])^(a[167] & b[365])^(a[166] & b[366])^(a[165] & b[367])^(a[164] & b[368])^(a[163] & b[369])^(a[162] & b[370])^(a[161] & b[371])^(a[160] & b[372])^(a[159] & b[373])^(a[158] & b[374])^(a[157] & b[375])^(a[156] & b[376])^(a[155] & b[377])^(a[154] & b[378])^(a[153] & b[379])^(a[152] & b[380])^(a[151] & b[381])^(a[150] & b[382])^(a[149] & b[383])^(a[148] & b[384])^(a[147] & b[385])^(a[146] & b[386])^(a[145] & b[387])^(a[144] & b[388])^(a[143] & b[389])^(a[142] & b[390])^(a[141] & b[391])^(a[140] & b[392])^(a[139] & b[393])^(a[138] & b[394])^(a[137] & b[395])^(a[136] & b[396])^(a[135] & b[397])^(a[134] & b[398])^(a[133] & b[399])^(a[132] & b[400])^(a[131] & b[401])^(a[130] & b[402])^(a[129] & b[403])^(a[128] & b[404])^(a[127] & b[405])^(a[126] & b[406])^(a[125] & b[407])^(a[124] & b[408]);
assign y[533] = (a[408] & b[125])^(a[407] & b[126])^(a[406] & b[127])^(a[405] & b[128])^(a[404] & b[129])^(a[403] & b[130])^(a[402] & b[131])^(a[401] & b[132])^(a[400] & b[133])^(a[399] & b[134])^(a[398] & b[135])^(a[397] & b[136])^(a[396] & b[137])^(a[395] & b[138])^(a[394] & b[139])^(a[393] & b[140])^(a[392] & b[141])^(a[391] & b[142])^(a[390] & b[143])^(a[389] & b[144])^(a[388] & b[145])^(a[387] & b[146])^(a[386] & b[147])^(a[385] & b[148])^(a[384] & b[149])^(a[383] & b[150])^(a[382] & b[151])^(a[381] & b[152])^(a[380] & b[153])^(a[379] & b[154])^(a[378] & b[155])^(a[377] & b[156])^(a[376] & b[157])^(a[375] & b[158])^(a[374] & b[159])^(a[373] & b[160])^(a[372] & b[161])^(a[371] & b[162])^(a[370] & b[163])^(a[369] & b[164])^(a[368] & b[165])^(a[367] & b[166])^(a[366] & b[167])^(a[365] & b[168])^(a[364] & b[169])^(a[363] & b[170])^(a[362] & b[171])^(a[361] & b[172])^(a[360] & b[173])^(a[359] & b[174])^(a[358] & b[175])^(a[357] & b[176])^(a[356] & b[177])^(a[355] & b[178])^(a[354] & b[179])^(a[353] & b[180])^(a[352] & b[181])^(a[351] & b[182])^(a[350] & b[183])^(a[349] & b[184])^(a[348] & b[185])^(a[347] & b[186])^(a[346] & b[187])^(a[345] & b[188])^(a[344] & b[189])^(a[343] & b[190])^(a[342] & b[191])^(a[341] & b[192])^(a[340] & b[193])^(a[339] & b[194])^(a[338] & b[195])^(a[337] & b[196])^(a[336] & b[197])^(a[335] & b[198])^(a[334] & b[199])^(a[333] & b[200])^(a[332] & b[201])^(a[331] & b[202])^(a[330] & b[203])^(a[329] & b[204])^(a[328] & b[205])^(a[327] & b[206])^(a[326] & b[207])^(a[325] & b[208])^(a[324] & b[209])^(a[323] & b[210])^(a[322] & b[211])^(a[321] & b[212])^(a[320] & b[213])^(a[319] & b[214])^(a[318] & b[215])^(a[317] & b[216])^(a[316] & b[217])^(a[315] & b[218])^(a[314] & b[219])^(a[313] & b[220])^(a[312] & b[221])^(a[311] & b[222])^(a[310] & b[223])^(a[309] & b[224])^(a[308] & b[225])^(a[307] & b[226])^(a[306] & b[227])^(a[305] & b[228])^(a[304] & b[229])^(a[303] & b[230])^(a[302] & b[231])^(a[301] & b[232])^(a[300] & b[233])^(a[299] & b[234])^(a[298] & b[235])^(a[297] & b[236])^(a[296] & b[237])^(a[295] & b[238])^(a[294] & b[239])^(a[293] & b[240])^(a[292] & b[241])^(a[291] & b[242])^(a[290] & b[243])^(a[289] & b[244])^(a[288] & b[245])^(a[287] & b[246])^(a[286] & b[247])^(a[285] & b[248])^(a[284] & b[249])^(a[283] & b[250])^(a[282] & b[251])^(a[281] & b[252])^(a[280] & b[253])^(a[279] & b[254])^(a[278] & b[255])^(a[277] & b[256])^(a[276] & b[257])^(a[275] & b[258])^(a[274] & b[259])^(a[273] & b[260])^(a[272] & b[261])^(a[271] & b[262])^(a[270] & b[263])^(a[269] & b[264])^(a[268] & b[265])^(a[267] & b[266])^(a[266] & b[267])^(a[265] & b[268])^(a[264] & b[269])^(a[263] & b[270])^(a[262] & b[271])^(a[261] & b[272])^(a[260] & b[273])^(a[259] & b[274])^(a[258] & b[275])^(a[257] & b[276])^(a[256] & b[277])^(a[255] & b[278])^(a[254] & b[279])^(a[253] & b[280])^(a[252] & b[281])^(a[251] & b[282])^(a[250] & b[283])^(a[249] & b[284])^(a[248] & b[285])^(a[247] & b[286])^(a[246] & b[287])^(a[245] & b[288])^(a[244] & b[289])^(a[243] & b[290])^(a[242] & b[291])^(a[241] & b[292])^(a[240] & b[293])^(a[239] & b[294])^(a[238] & b[295])^(a[237] & b[296])^(a[236] & b[297])^(a[235] & b[298])^(a[234] & b[299])^(a[233] & b[300])^(a[232] & b[301])^(a[231] & b[302])^(a[230] & b[303])^(a[229] & b[304])^(a[228] & b[305])^(a[227] & b[306])^(a[226] & b[307])^(a[225] & b[308])^(a[224] & b[309])^(a[223] & b[310])^(a[222] & b[311])^(a[221] & b[312])^(a[220] & b[313])^(a[219] & b[314])^(a[218] & b[315])^(a[217] & b[316])^(a[216] & b[317])^(a[215] & b[318])^(a[214] & b[319])^(a[213] & b[320])^(a[212] & b[321])^(a[211] & b[322])^(a[210] & b[323])^(a[209] & b[324])^(a[208] & b[325])^(a[207] & b[326])^(a[206] & b[327])^(a[205] & b[328])^(a[204] & b[329])^(a[203] & b[330])^(a[202] & b[331])^(a[201] & b[332])^(a[200] & b[333])^(a[199] & b[334])^(a[198] & b[335])^(a[197] & b[336])^(a[196] & b[337])^(a[195] & b[338])^(a[194] & b[339])^(a[193] & b[340])^(a[192] & b[341])^(a[191] & b[342])^(a[190] & b[343])^(a[189] & b[344])^(a[188] & b[345])^(a[187] & b[346])^(a[186] & b[347])^(a[185] & b[348])^(a[184] & b[349])^(a[183] & b[350])^(a[182] & b[351])^(a[181] & b[352])^(a[180] & b[353])^(a[179] & b[354])^(a[178] & b[355])^(a[177] & b[356])^(a[176] & b[357])^(a[175] & b[358])^(a[174] & b[359])^(a[173] & b[360])^(a[172] & b[361])^(a[171] & b[362])^(a[170] & b[363])^(a[169] & b[364])^(a[168] & b[365])^(a[167] & b[366])^(a[166] & b[367])^(a[165] & b[368])^(a[164] & b[369])^(a[163] & b[370])^(a[162] & b[371])^(a[161] & b[372])^(a[160] & b[373])^(a[159] & b[374])^(a[158] & b[375])^(a[157] & b[376])^(a[156] & b[377])^(a[155] & b[378])^(a[154] & b[379])^(a[153] & b[380])^(a[152] & b[381])^(a[151] & b[382])^(a[150] & b[383])^(a[149] & b[384])^(a[148] & b[385])^(a[147] & b[386])^(a[146] & b[387])^(a[145] & b[388])^(a[144] & b[389])^(a[143] & b[390])^(a[142] & b[391])^(a[141] & b[392])^(a[140] & b[393])^(a[139] & b[394])^(a[138] & b[395])^(a[137] & b[396])^(a[136] & b[397])^(a[135] & b[398])^(a[134] & b[399])^(a[133] & b[400])^(a[132] & b[401])^(a[131] & b[402])^(a[130] & b[403])^(a[129] & b[404])^(a[128] & b[405])^(a[127] & b[406])^(a[126] & b[407])^(a[125] & b[408]);
assign y[534] = (a[408] & b[126])^(a[407] & b[127])^(a[406] & b[128])^(a[405] & b[129])^(a[404] & b[130])^(a[403] & b[131])^(a[402] & b[132])^(a[401] & b[133])^(a[400] & b[134])^(a[399] & b[135])^(a[398] & b[136])^(a[397] & b[137])^(a[396] & b[138])^(a[395] & b[139])^(a[394] & b[140])^(a[393] & b[141])^(a[392] & b[142])^(a[391] & b[143])^(a[390] & b[144])^(a[389] & b[145])^(a[388] & b[146])^(a[387] & b[147])^(a[386] & b[148])^(a[385] & b[149])^(a[384] & b[150])^(a[383] & b[151])^(a[382] & b[152])^(a[381] & b[153])^(a[380] & b[154])^(a[379] & b[155])^(a[378] & b[156])^(a[377] & b[157])^(a[376] & b[158])^(a[375] & b[159])^(a[374] & b[160])^(a[373] & b[161])^(a[372] & b[162])^(a[371] & b[163])^(a[370] & b[164])^(a[369] & b[165])^(a[368] & b[166])^(a[367] & b[167])^(a[366] & b[168])^(a[365] & b[169])^(a[364] & b[170])^(a[363] & b[171])^(a[362] & b[172])^(a[361] & b[173])^(a[360] & b[174])^(a[359] & b[175])^(a[358] & b[176])^(a[357] & b[177])^(a[356] & b[178])^(a[355] & b[179])^(a[354] & b[180])^(a[353] & b[181])^(a[352] & b[182])^(a[351] & b[183])^(a[350] & b[184])^(a[349] & b[185])^(a[348] & b[186])^(a[347] & b[187])^(a[346] & b[188])^(a[345] & b[189])^(a[344] & b[190])^(a[343] & b[191])^(a[342] & b[192])^(a[341] & b[193])^(a[340] & b[194])^(a[339] & b[195])^(a[338] & b[196])^(a[337] & b[197])^(a[336] & b[198])^(a[335] & b[199])^(a[334] & b[200])^(a[333] & b[201])^(a[332] & b[202])^(a[331] & b[203])^(a[330] & b[204])^(a[329] & b[205])^(a[328] & b[206])^(a[327] & b[207])^(a[326] & b[208])^(a[325] & b[209])^(a[324] & b[210])^(a[323] & b[211])^(a[322] & b[212])^(a[321] & b[213])^(a[320] & b[214])^(a[319] & b[215])^(a[318] & b[216])^(a[317] & b[217])^(a[316] & b[218])^(a[315] & b[219])^(a[314] & b[220])^(a[313] & b[221])^(a[312] & b[222])^(a[311] & b[223])^(a[310] & b[224])^(a[309] & b[225])^(a[308] & b[226])^(a[307] & b[227])^(a[306] & b[228])^(a[305] & b[229])^(a[304] & b[230])^(a[303] & b[231])^(a[302] & b[232])^(a[301] & b[233])^(a[300] & b[234])^(a[299] & b[235])^(a[298] & b[236])^(a[297] & b[237])^(a[296] & b[238])^(a[295] & b[239])^(a[294] & b[240])^(a[293] & b[241])^(a[292] & b[242])^(a[291] & b[243])^(a[290] & b[244])^(a[289] & b[245])^(a[288] & b[246])^(a[287] & b[247])^(a[286] & b[248])^(a[285] & b[249])^(a[284] & b[250])^(a[283] & b[251])^(a[282] & b[252])^(a[281] & b[253])^(a[280] & b[254])^(a[279] & b[255])^(a[278] & b[256])^(a[277] & b[257])^(a[276] & b[258])^(a[275] & b[259])^(a[274] & b[260])^(a[273] & b[261])^(a[272] & b[262])^(a[271] & b[263])^(a[270] & b[264])^(a[269] & b[265])^(a[268] & b[266])^(a[267] & b[267])^(a[266] & b[268])^(a[265] & b[269])^(a[264] & b[270])^(a[263] & b[271])^(a[262] & b[272])^(a[261] & b[273])^(a[260] & b[274])^(a[259] & b[275])^(a[258] & b[276])^(a[257] & b[277])^(a[256] & b[278])^(a[255] & b[279])^(a[254] & b[280])^(a[253] & b[281])^(a[252] & b[282])^(a[251] & b[283])^(a[250] & b[284])^(a[249] & b[285])^(a[248] & b[286])^(a[247] & b[287])^(a[246] & b[288])^(a[245] & b[289])^(a[244] & b[290])^(a[243] & b[291])^(a[242] & b[292])^(a[241] & b[293])^(a[240] & b[294])^(a[239] & b[295])^(a[238] & b[296])^(a[237] & b[297])^(a[236] & b[298])^(a[235] & b[299])^(a[234] & b[300])^(a[233] & b[301])^(a[232] & b[302])^(a[231] & b[303])^(a[230] & b[304])^(a[229] & b[305])^(a[228] & b[306])^(a[227] & b[307])^(a[226] & b[308])^(a[225] & b[309])^(a[224] & b[310])^(a[223] & b[311])^(a[222] & b[312])^(a[221] & b[313])^(a[220] & b[314])^(a[219] & b[315])^(a[218] & b[316])^(a[217] & b[317])^(a[216] & b[318])^(a[215] & b[319])^(a[214] & b[320])^(a[213] & b[321])^(a[212] & b[322])^(a[211] & b[323])^(a[210] & b[324])^(a[209] & b[325])^(a[208] & b[326])^(a[207] & b[327])^(a[206] & b[328])^(a[205] & b[329])^(a[204] & b[330])^(a[203] & b[331])^(a[202] & b[332])^(a[201] & b[333])^(a[200] & b[334])^(a[199] & b[335])^(a[198] & b[336])^(a[197] & b[337])^(a[196] & b[338])^(a[195] & b[339])^(a[194] & b[340])^(a[193] & b[341])^(a[192] & b[342])^(a[191] & b[343])^(a[190] & b[344])^(a[189] & b[345])^(a[188] & b[346])^(a[187] & b[347])^(a[186] & b[348])^(a[185] & b[349])^(a[184] & b[350])^(a[183] & b[351])^(a[182] & b[352])^(a[181] & b[353])^(a[180] & b[354])^(a[179] & b[355])^(a[178] & b[356])^(a[177] & b[357])^(a[176] & b[358])^(a[175] & b[359])^(a[174] & b[360])^(a[173] & b[361])^(a[172] & b[362])^(a[171] & b[363])^(a[170] & b[364])^(a[169] & b[365])^(a[168] & b[366])^(a[167] & b[367])^(a[166] & b[368])^(a[165] & b[369])^(a[164] & b[370])^(a[163] & b[371])^(a[162] & b[372])^(a[161] & b[373])^(a[160] & b[374])^(a[159] & b[375])^(a[158] & b[376])^(a[157] & b[377])^(a[156] & b[378])^(a[155] & b[379])^(a[154] & b[380])^(a[153] & b[381])^(a[152] & b[382])^(a[151] & b[383])^(a[150] & b[384])^(a[149] & b[385])^(a[148] & b[386])^(a[147] & b[387])^(a[146] & b[388])^(a[145] & b[389])^(a[144] & b[390])^(a[143] & b[391])^(a[142] & b[392])^(a[141] & b[393])^(a[140] & b[394])^(a[139] & b[395])^(a[138] & b[396])^(a[137] & b[397])^(a[136] & b[398])^(a[135] & b[399])^(a[134] & b[400])^(a[133] & b[401])^(a[132] & b[402])^(a[131] & b[403])^(a[130] & b[404])^(a[129] & b[405])^(a[128] & b[406])^(a[127] & b[407])^(a[126] & b[408]);
assign y[535] = (a[408] & b[127])^(a[407] & b[128])^(a[406] & b[129])^(a[405] & b[130])^(a[404] & b[131])^(a[403] & b[132])^(a[402] & b[133])^(a[401] & b[134])^(a[400] & b[135])^(a[399] & b[136])^(a[398] & b[137])^(a[397] & b[138])^(a[396] & b[139])^(a[395] & b[140])^(a[394] & b[141])^(a[393] & b[142])^(a[392] & b[143])^(a[391] & b[144])^(a[390] & b[145])^(a[389] & b[146])^(a[388] & b[147])^(a[387] & b[148])^(a[386] & b[149])^(a[385] & b[150])^(a[384] & b[151])^(a[383] & b[152])^(a[382] & b[153])^(a[381] & b[154])^(a[380] & b[155])^(a[379] & b[156])^(a[378] & b[157])^(a[377] & b[158])^(a[376] & b[159])^(a[375] & b[160])^(a[374] & b[161])^(a[373] & b[162])^(a[372] & b[163])^(a[371] & b[164])^(a[370] & b[165])^(a[369] & b[166])^(a[368] & b[167])^(a[367] & b[168])^(a[366] & b[169])^(a[365] & b[170])^(a[364] & b[171])^(a[363] & b[172])^(a[362] & b[173])^(a[361] & b[174])^(a[360] & b[175])^(a[359] & b[176])^(a[358] & b[177])^(a[357] & b[178])^(a[356] & b[179])^(a[355] & b[180])^(a[354] & b[181])^(a[353] & b[182])^(a[352] & b[183])^(a[351] & b[184])^(a[350] & b[185])^(a[349] & b[186])^(a[348] & b[187])^(a[347] & b[188])^(a[346] & b[189])^(a[345] & b[190])^(a[344] & b[191])^(a[343] & b[192])^(a[342] & b[193])^(a[341] & b[194])^(a[340] & b[195])^(a[339] & b[196])^(a[338] & b[197])^(a[337] & b[198])^(a[336] & b[199])^(a[335] & b[200])^(a[334] & b[201])^(a[333] & b[202])^(a[332] & b[203])^(a[331] & b[204])^(a[330] & b[205])^(a[329] & b[206])^(a[328] & b[207])^(a[327] & b[208])^(a[326] & b[209])^(a[325] & b[210])^(a[324] & b[211])^(a[323] & b[212])^(a[322] & b[213])^(a[321] & b[214])^(a[320] & b[215])^(a[319] & b[216])^(a[318] & b[217])^(a[317] & b[218])^(a[316] & b[219])^(a[315] & b[220])^(a[314] & b[221])^(a[313] & b[222])^(a[312] & b[223])^(a[311] & b[224])^(a[310] & b[225])^(a[309] & b[226])^(a[308] & b[227])^(a[307] & b[228])^(a[306] & b[229])^(a[305] & b[230])^(a[304] & b[231])^(a[303] & b[232])^(a[302] & b[233])^(a[301] & b[234])^(a[300] & b[235])^(a[299] & b[236])^(a[298] & b[237])^(a[297] & b[238])^(a[296] & b[239])^(a[295] & b[240])^(a[294] & b[241])^(a[293] & b[242])^(a[292] & b[243])^(a[291] & b[244])^(a[290] & b[245])^(a[289] & b[246])^(a[288] & b[247])^(a[287] & b[248])^(a[286] & b[249])^(a[285] & b[250])^(a[284] & b[251])^(a[283] & b[252])^(a[282] & b[253])^(a[281] & b[254])^(a[280] & b[255])^(a[279] & b[256])^(a[278] & b[257])^(a[277] & b[258])^(a[276] & b[259])^(a[275] & b[260])^(a[274] & b[261])^(a[273] & b[262])^(a[272] & b[263])^(a[271] & b[264])^(a[270] & b[265])^(a[269] & b[266])^(a[268] & b[267])^(a[267] & b[268])^(a[266] & b[269])^(a[265] & b[270])^(a[264] & b[271])^(a[263] & b[272])^(a[262] & b[273])^(a[261] & b[274])^(a[260] & b[275])^(a[259] & b[276])^(a[258] & b[277])^(a[257] & b[278])^(a[256] & b[279])^(a[255] & b[280])^(a[254] & b[281])^(a[253] & b[282])^(a[252] & b[283])^(a[251] & b[284])^(a[250] & b[285])^(a[249] & b[286])^(a[248] & b[287])^(a[247] & b[288])^(a[246] & b[289])^(a[245] & b[290])^(a[244] & b[291])^(a[243] & b[292])^(a[242] & b[293])^(a[241] & b[294])^(a[240] & b[295])^(a[239] & b[296])^(a[238] & b[297])^(a[237] & b[298])^(a[236] & b[299])^(a[235] & b[300])^(a[234] & b[301])^(a[233] & b[302])^(a[232] & b[303])^(a[231] & b[304])^(a[230] & b[305])^(a[229] & b[306])^(a[228] & b[307])^(a[227] & b[308])^(a[226] & b[309])^(a[225] & b[310])^(a[224] & b[311])^(a[223] & b[312])^(a[222] & b[313])^(a[221] & b[314])^(a[220] & b[315])^(a[219] & b[316])^(a[218] & b[317])^(a[217] & b[318])^(a[216] & b[319])^(a[215] & b[320])^(a[214] & b[321])^(a[213] & b[322])^(a[212] & b[323])^(a[211] & b[324])^(a[210] & b[325])^(a[209] & b[326])^(a[208] & b[327])^(a[207] & b[328])^(a[206] & b[329])^(a[205] & b[330])^(a[204] & b[331])^(a[203] & b[332])^(a[202] & b[333])^(a[201] & b[334])^(a[200] & b[335])^(a[199] & b[336])^(a[198] & b[337])^(a[197] & b[338])^(a[196] & b[339])^(a[195] & b[340])^(a[194] & b[341])^(a[193] & b[342])^(a[192] & b[343])^(a[191] & b[344])^(a[190] & b[345])^(a[189] & b[346])^(a[188] & b[347])^(a[187] & b[348])^(a[186] & b[349])^(a[185] & b[350])^(a[184] & b[351])^(a[183] & b[352])^(a[182] & b[353])^(a[181] & b[354])^(a[180] & b[355])^(a[179] & b[356])^(a[178] & b[357])^(a[177] & b[358])^(a[176] & b[359])^(a[175] & b[360])^(a[174] & b[361])^(a[173] & b[362])^(a[172] & b[363])^(a[171] & b[364])^(a[170] & b[365])^(a[169] & b[366])^(a[168] & b[367])^(a[167] & b[368])^(a[166] & b[369])^(a[165] & b[370])^(a[164] & b[371])^(a[163] & b[372])^(a[162] & b[373])^(a[161] & b[374])^(a[160] & b[375])^(a[159] & b[376])^(a[158] & b[377])^(a[157] & b[378])^(a[156] & b[379])^(a[155] & b[380])^(a[154] & b[381])^(a[153] & b[382])^(a[152] & b[383])^(a[151] & b[384])^(a[150] & b[385])^(a[149] & b[386])^(a[148] & b[387])^(a[147] & b[388])^(a[146] & b[389])^(a[145] & b[390])^(a[144] & b[391])^(a[143] & b[392])^(a[142] & b[393])^(a[141] & b[394])^(a[140] & b[395])^(a[139] & b[396])^(a[138] & b[397])^(a[137] & b[398])^(a[136] & b[399])^(a[135] & b[400])^(a[134] & b[401])^(a[133] & b[402])^(a[132] & b[403])^(a[131] & b[404])^(a[130] & b[405])^(a[129] & b[406])^(a[128] & b[407])^(a[127] & b[408]);
assign y[536] = (a[408] & b[128])^(a[407] & b[129])^(a[406] & b[130])^(a[405] & b[131])^(a[404] & b[132])^(a[403] & b[133])^(a[402] & b[134])^(a[401] & b[135])^(a[400] & b[136])^(a[399] & b[137])^(a[398] & b[138])^(a[397] & b[139])^(a[396] & b[140])^(a[395] & b[141])^(a[394] & b[142])^(a[393] & b[143])^(a[392] & b[144])^(a[391] & b[145])^(a[390] & b[146])^(a[389] & b[147])^(a[388] & b[148])^(a[387] & b[149])^(a[386] & b[150])^(a[385] & b[151])^(a[384] & b[152])^(a[383] & b[153])^(a[382] & b[154])^(a[381] & b[155])^(a[380] & b[156])^(a[379] & b[157])^(a[378] & b[158])^(a[377] & b[159])^(a[376] & b[160])^(a[375] & b[161])^(a[374] & b[162])^(a[373] & b[163])^(a[372] & b[164])^(a[371] & b[165])^(a[370] & b[166])^(a[369] & b[167])^(a[368] & b[168])^(a[367] & b[169])^(a[366] & b[170])^(a[365] & b[171])^(a[364] & b[172])^(a[363] & b[173])^(a[362] & b[174])^(a[361] & b[175])^(a[360] & b[176])^(a[359] & b[177])^(a[358] & b[178])^(a[357] & b[179])^(a[356] & b[180])^(a[355] & b[181])^(a[354] & b[182])^(a[353] & b[183])^(a[352] & b[184])^(a[351] & b[185])^(a[350] & b[186])^(a[349] & b[187])^(a[348] & b[188])^(a[347] & b[189])^(a[346] & b[190])^(a[345] & b[191])^(a[344] & b[192])^(a[343] & b[193])^(a[342] & b[194])^(a[341] & b[195])^(a[340] & b[196])^(a[339] & b[197])^(a[338] & b[198])^(a[337] & b[199])^(a[336] & b[200])^(a[335] & b[201])^(a[334] & b[202])^(a[333] & b[203])^(a[332] & b[204])^(a[331] & b[205])^(a[330] & b[206])^(a[329] & b[207])^(a[328] & b[208])^(a[327] & b[209])^(a[326] & b[210])^(a[325] & b[211])^(a[324] & b[212])^(a[323] & b[213])^(a[322] & b[214])^(a[321] & b[215])^(a[320] & b[216])^(a[319] & b[217])^(a[318] & b[218])^(a[317] & b[219])^(a[316] & b[220])^(a[315] & b[221])^(a[314] & b[222])^(a[313] & b[223])^(a[312] & b[224])^(a[311] & b[225])^(a[310] & b[226])^(a[309] & b[227])^(a[308] & b[228])^(a[307] & b[229])^(a[306] & b[230])^(a[305] & b[231])^(a[304] & b[232])^(a[303] & b[233])^(a[302] & b[234])^(a[301] & b[235])^(a[300] & b[236])^(a[299] & b[237])^(a[298] & b[238])^(a[297] & b[239])^(a[296] & b[240])^(a[295] & b[241])^(a[294] & b[242])^(a[293] & b[243])^(a[292] & b[244])^(a[291] & b[245])^(a[290] & b[246])^(a[289] & b[247])^(a[288] & b[248])^(a[287] & b[249])^(a[286] & b[250])^(a[285] & b[251])^(a[284] & b[252])^(a[283] & b[253])^(a[282] & b[254])^(a[281] & b[255])^(a[280] & b[256])^(a[279] & b[257])^(a[278] & b[258])^(a[277] & b[259])^(a[276] & b[260])^(a[275] & b[261])^(a[274] & b[262])^(a[273] & b[263])^(a[272] & b[264])^(a[271] & b[265])^(a[270] & b[266])^(a[269] & b[267])^(a[268] & b[268])^(a[267] & b[269])^(a[266] & b[270])^(a[265] & b[271])^(a[264] & b[272])^(a[263] & b[273])^(a[262] & b[274])^(a[261] & b[275])^(a[260] & b[276])^(a[259] & b[277])^(a[258] & b[278])^(a[257] & b[279])^(a[256] & b[280])^(a[255] & b[281])^(a[254] & b[282])^(a[253] & b[283])^(a[252] & b[284])^(a[251] & b[285])^(a[250] & b[286])^(a[249] & b[287])^(a[248] & b[288])^(a[247] & b[289])^(a[246] & b[290])^(a[245] & b[291])^(a[244] & b[292])^(a[243] & b[293])^(a[242] & b[294])^(a[241] & b[295])^(a[240] & b[296])^(a[239] & b[297])^(a[238] & b[298])^(a[237] & b[299])^(a[236] & b[300])^(a[235] & b[301])^(a[234] & b[302])^(a[233] & b[303])^(a[232] & b[304])^(a[231] & b[305])^(a[230] & b[306])^(a[229] & b[307])^(a[228] & b[308])^(a[227] & b[309])^(a[226] & b[310])^(a[225] & b[311])^(a[224] & b[312])^(a[223] & b[313])^(a[222] & b[314])^(a[221] & b[315])^(a[220] & b[316])^(a[219] & b[317])^(a[218] & b[318])^(a[217] & b[319])^(a[216] & b[320])^(a[215] & b[321])^(a[214] & b[322])^(a[213] & b[323])^(a[212] & b[324])^(a[211] & b[325])^(a[210] & b[326])^(a[209] & b[327])^(a[208] & b[328])^(a[207] & b[329])^(a[206] & b[330])^(a[205] & b[331])^(a[204] & b[332])^(a[203] & b[333])^(a[202] & b[334])^(a[201] & b[335])^(a[200] & b[336])^(a[199] & b[337])^(a[198] & b[338])^(a[197] & b[339])^(a[196] & b[340])^(a[195] & b[341])^(a[194] & b[342])^(a[193] & b[343])^(a[192] & b[344])^(a[191] & b[345])^(a[190] & b[346])^(a[189] & b[347])^(a[188] & b[348])^(a[187] & b[349])^(a[186] & b[350])^(a[185] & b[351])^(a[184] & b[352])^(a[183] & b[353])^(a[182] & b[354])^(a[181] & b[355])^(a[180] & b[356])^(a[179] & b[357])^(a[178] & b[358])^(a[177] & b[359])^(a[176] & b[360])^(a[175] & b[361])^(a[174] & b[362])^(a[173] & b[363])^(a[172] & b[364])^(a[171] & b[365])^(a[170] & b[366])^(a[169] & b[367])^(a[168] & b[368])^(a[167] & b[369])^(a[166] & b[370])^(a[165] & b[371])^(a[164] & b[372])^(a[163] & b[373])^(a[162] & b[374])^(a[161] & b[375])^(a[160] & b[376])^(a[159] & b[377])^(a[158] & b[378])^(a[157] & b[379])^(a[156] & b[380])^(a[155] & b[381])^(a[154] & b[382])^(a[153] & b[383])^(a[152] & b[384])^(a[151] & b[385])^(a[150] & b[386])^(a[149] & b[387])^(a[148] & b[388])^(a[147] & b[389])^(a[146] & b[390])^(a[145] & b[391])^(a[144] & b[392])^(a[143] & b[393])^(a[142] & b[394])^(a[141] & b[395])^(a[140] & b[396])^(a[139] & b[397])^(a[138] & b[398])^(a[137] & b[399])^(a[136] & b[400])^(a[135] & b[401])^(a[134] & b[402])^(a[133] & b[403])^(a[132] & b[404])^(a[131] & b[405])^(a[130] & b[406])^(a[129] & b[407])^(a[128] & b[408]);
assign y[537] = (a[408] & b[129])^(a[407] & b[130])^(a[406] & b[131])^(a[405] & b[132])^(a[404] & b[133])^(a[403] & b[134])^(a[402] & b[135])^(a[401] & b[136])^(a[400] & b[137])^(a[399] & b[138])^(a[398] & b[139])^(a[397] & b[140])^(a[396] & b[141])^(a[395] & b[142])^(a[394] & b[143])^(a[393] & b[144])^(a[392] & b[145])^(a[391] & b[146])^(a[390] & b[147])^(a[389] & b[148])^(a[388] & b[149])^(a[387] & b[150])^(a[386] & b[151])^(a[385] & b[152])^(a[384] & b[153])^(a[383] & b[154])^(a[382] & b[155])^(a[381] & b[156])^(a[380] & b[157])^(a[379] & b[158])^(a[378] & b[159])^(a[377] & b[160])^(a[376] & b[161])^(a[375] & b[162])^(a[374] & b[163])^(a[373] & b[164])^(a[372] & b[165])^(a[371] & b[166])^(a[370] & b[167])^(a[369] & b[168])^(a[368] & b[169])^(a[367] & b[170])^(a[366] & b[171])^(a[365] & b[172])^(a[364] & b[173])^(a[363] & b[174])^(a[362] & b[175])^(a[361] & b[176])^(a[360] & b[177])^(a[359] & b[178])^(a[358] & b[179])^(a[357] & b[180])^(a[356] & b[181])^(a[355] & b[182])^(a[354] & b[183])^(a[353] & b[184])^(a[352] & b[185])^(a[351] & b[186])^(a[350] & b[187])^(a[349] & b[188])^(a[348] & b[189])^(a[347] & b[190])^(a[346] & b[191])^(a[345] & b[192])^(a[344] & b[193])^(a[343] & b[194])^(a[342] & b[195])^(a[341] & b[196])^(a[340] & b[197])^(a[339] & b[198])^(a[338] & b[199])^(a[337] & b[200])^(a[336] & b[201])^(a[335] & b[202])^(a[334] & b[203])^(a[333] & b[204])^(a[332] & b[205])^(a[331] & b[206])^(a[330] & b[207])^(a[329] & b[208])^(a[328] & b[209])^(a[327] & b[210])^(a[326] & b[211])^(a[325] & b[212])^(a[324] & b[213])^(a[323] & b[214])^(a[322] & b[215])^(a[321] & b[216])^(a[320] & b[217])^(a[319] & b[218])^(a[318] & b[219])^(a[317] & b[220])^(a[316] & b[221])^(a[315] & b[222])^(a[314] & b[223])^(a[313] & b[224])^(a[312] & b[225])^(a[311] & b[226])^(a[310] & b[227])^(a[309] & b[228])^(a[308] & b[229])^(a[307] & b[230])^(a[306] & b[231])^(a[305] & b[232])^(a[304] & b[233])^(a[303] & b[234])^(a[302] & b[235])^(a[301] & b[236])^(a[300] & b[237])^(a[299] & b[238])^(a[298] & b[239])^(a[297] & b[240])^(a[296] & b[241])^(a[295] & b[242])^(a[294] & b[243])^(a[293] & b[244])^(a[292] & b[245])^(a[291] & b[246])^(a[290] & b[247])^(a[289] & b[248])^(a[288] & b[249])^(a[287] & b[250])^(a[286] & b[251])^(a[285] & b[252])^(a[284] & b[253])^(a[283] & b[254])^(a[282] & b[255])^(a[281] & b[256])^(a[280] & b[257])^(a[279] & b[258])^(a[278] & b[259])^(a[277] & b[260])^(a[276] & b[261])^(a[275] & b[262])^(a[274] & b[263])^(a[273] & b[264])^(a[272] & b[265])^(a[271] & b[266])^(a[270] & b[267])^(a[269] & b[268])^(a[268] & b[269])^(a[267] & b[270])^(a[266] & b[271])^(a[265] & b[272])^(a[264] & b[273])^(a[263] & b[274])^(a[262] & b[275])^(a[261] & b[276])^(a[260] & b[277])^(a[259] & b[278])^(a[258] & b[279])^(a[257] & b[280])^(a[256] & b[281])^(a[255] & b[282])^(a[254] & b[283])^(a[253] & b[284])^(a[252] & b[285])^(a[251] & b[286])^(a[250] & b[287])^(a[249] & b[288])^(a[248] & b[289])^(a[247] & b[290])^(a[246] & b[291])^(a[245] & b[292])^(a[244] & b[293])^(a[243] & b[294])^(a[242] & b[295])^(a[241] & b[296])^(a[240] & b[297])^(a[239] & b[298])^(a[238] & b[299])^(a[237] & b[300])^(a[236] & b[301])^(a[235] & b[302])^(a[234] & b[303])^(a[233] & b[304])^(a[232] & b[305])^(a[231] & b[306])^(a[230] & b[307])^(a[229] & b[308])^(a[228] & b[309])^(a[227] & b[310])^(a[226] & b[311])^(a[225] & b[312])^(a[224] & b[313])^(a[223] & b[314])^(a[222] & b[315])^(a[221] & b[316])^(a[220] & b[317])^(a[219] & b[318])^(a[218] & b[319])^(a[217] & b[320])^(a[216] & b[321])^(a[215] & b[322])^(a[214] & b[323])^(a[213] & b[324])^(a[212] & b[325])^(a[211] & b[326])^(a[210] & b[327])^(a[209] & b[328])^(a[208] & b[329])^(a[207] & b[330])^(a[206] & b[331])^(a[205] & b[332])^(a[204] & b[333])^(a[203] & b[334])^(a[202] & b[335])^(a[201] & b[336])^(a[200] & b[337])^(a[199] & b[338])^(a[198] & b[339])^(a[197] & b[340])^(a[196] & b[341])^(a[195] & b[342])^(a[194] & b[343])^(a[193] & b[344])^(a[192] & b[345])^(a[191] & b[346])^(a[190] & b[347])^(a[189] & b[348])^(a[188] & b[349])^(a[187] & b[350])^(a[186] & b[351])^(a[185] & b[352])^(a[184] & b[353])^(a[183] & b[354])^(a[182] & b[355])^(a[181] & b[356])^(a[180] & b[357])^(a[179] & b[358])^(a[178] & b[359])^(a[177] & b[360])^(a[176] & b[361])^(a[175] & b[362])^(a[174] & b[363])^(a[173] & b[364])^(a[172] & b[365])^(a[171] & b[366])^(a[170] & b[367])^(a[169] & b[368])^(a[168] & b[369])^(a[167] & b[370])^(a[166] & b[371])^(a[165] & b[372])^(a[164] & b[373])^(a[163] & b[374])^(a[162] & b[375])^(a[161] & b[376])^(a[160] & b[377])^(a[159] & b[378])^(a[158] & b[379])^(a[157] & b[380])^(a[156] & b[381])^(a[155] & b[382])^(a[154] & b[383])^(a[153] & b[384])^(a[152] & b[385])^(a[151] & b[386])^(a[150] & b[387])^(a[149] & b[388])^(a[148] & b[389])^(a[147] & b[390])^(a[146] & b[391])^(a[145] & b[392])^(a[144] & b[393])^(a[143] & b[394])^(a[142] & b[395])^(a[141] & b[396])^(a[140] & b[397])^(a[139] & b[398])^(a[138] & b[399])^(a[137] & b[400])^(a[136] & b[401])^(a[135] & b[402])^(a[134] & b[403])^(a[133] & b[404])^(a[132] & b[405])^(a[131] & b[406])^(a[130] & b[407])^(a[129] & b[408]);
assign y[538] = (a[408] & b[130])^(a[407] & b[131])^(a[406] & b[132])^(a[405] & b[133])^(a[404] & b[134])^(a[403] & b[135])^(a[402] & b[136])^(a[401] & b[137])^(a[400] & b[138])^(a[399] & b[139])^(a[398] & b[140])^(a[397] & b[141])^(a[396] & b[142])^(a[395] & b[143])^(a[394] & b[144])^(a[393] & b[145])^(a[392] & b[146])^(a[391] & b[147])^(a[390] & b[148])^(a[389] & b[149])^(a[388] & b[150])^(a[387] & b[151])^(a[386] & b[152])^(a[385] & b[153])^(a[384] & b[154])^(a[383] & b[155])^(a[382] & b[156])^(a[381] & b[157])^(a[380] & b[158])^(a[379] & b[159])^(a[378] & b[160])^(a[377] & b[161])^(a[376] & b[162])^(a[375] & b[163])^(a[374] & b[164])^(a[373] & b[165])^(a[372] & b[166])^(a[371] & b[167])^(a[370] & b[168])^(a[369] & b[169])^(a[368] & b[170])^(a[367] & b[171])^(a[366] & b[172])^(a[365] & b[173])^(a[364] & b[174])^(a[363] & b[175])^(a[362] & b[176])^(a[361] & b[177])^(a[360] & b[178])^(a[359] & b[179])^(a[358] & b[180])^(a[357] & b[181])^(a[356] & b[182])^(a[355] & b[183])^(a[354] & b[184])^(a[353] & b[185])^(a[352] & b[186])^(a[351] & b[187])^(a[350] & b[188])^(a[349] & b[189])^(a[348] & b[190])^(a[347] & b[191])^(a[346] & b[192])^(a[345] & b[193])^(a[344] & b[194])^(a[343] & b[195])^(a[342] & b[196])^(a[341] & b[197])^(a[340] & b[198])^(a[339] & b[199])^(a[338] & b[200])^(a[337] & b[201])^(a[336] & b[202])^(a[335] & b[203])^(a[334] & b[204])^(a[333] & b[205])^(a[332] & b[206])^(a[331] & b[207])^(a[330] & b[208])^(a[329] & b[209])^(a[328] & b[210])^(a[327] & b[211])^(a[326] & b[212])^(a[325] & b[213])^(a[324] & b[214])^(a[323] & b[215])^(a[322] & b[216])^(a[321] & b[217])^(a[320] & b[218])^(a[319] & b[219])^(a[318] & b[220])^(a[317] & b[221])^(a[316] & b[222])^(a[315] & b[223])^(a[314] & b[224])^(a[313] & b[225])^(a[312] & b[226])^(a[311] & b[227])^(a[310] & b[228])^(a[309] & b[229])^(a[308] & b[230])^(a[307] & b[231])^(a[306] & b[232])^(a[305] & b[233])^(a[304] & b[234])^(a[303] & b[235])^(a[302] & b[236])^(a[301] & b[237])^(a[300] & b[238])^(a[299] & b[239])^(a[298] & b[240])^(a[297] & b[241])^(a[296] & b[242])^(a[295] & b[243])^(a[294] & b[244])^(a[293] & b[245])^(a[292] & b[246])^(a[291] & b[247])^(a[290] & b[248])^(a[289] & b[249])^(a[288] & b[250])^(a[287] & b[251])^(a[286] & b[252])^(a[285] & b[253])^(a[284] & b[254])^(a[283] & b[255])^(a[282] & b[256])^(a[281] & b[257])^(a[280] & b[258])^(a[279] & b[259])^(a[278] & b[260])^(a[277] & b[261])^(a[276] & b[262])^(a[275] & b[263])^(a[274] & b[264])^(a[273] & b[265])^(a[272] & b[266])^(a[271] & b[267])^(a[270] & b[268])^(a[269] & b[269])^(a[268] & b[270])^(a[267] & b[271])^(a[266] & b[272])^(a[265] & b[273])^(a[264] & b[274])^(a[263] & b[275])^(a[262] & b[276])^(a[261] & b[277])^(a[260] & b[278])^(a[259] & b[279])^(a[258] & b[280])^(a[257] & b[281])^(a[256] & b[282])^(a[255] & b[283])^(a[254] & b[284])^(a[253] & b[285])^(a[252] & b[286])^(a[251] & b[287])^(a[250] & b[288])^(a[249] & b[289])^(a[248] & b[290])^(a[247] & b[291])^(a[246] & b[292])^(a[245] & b[293])^(a[244] & b[294])^(a[243] & b[295])^(a[242] & b[296])^(a[241] & b[297])^(a[240] & b[298])^(a[239] & b[299])^(a[238] & b[300])^(a[237] & b[301])^(a[236] & b[302])^(a[235] & b[303])^(a[234] & b[304])^(a[233] & b[305])^(a[232] & b[306])^(a[231] & b[307])^(a[230] & b[308])^(a[229] & b[309])^(a[228] & b[310])^(a[227] & b[311])^(a[226] & b[312])^(a[225] & b[313])^(a[224] & b[314])^(a[223] & b[315])^(a[222] & b[316])^(a[221] & b[317])^(a[220] & b[318])^(a[219] & b[319])^(a[218] & b[320])^(a[217] & b[321])^(a[216] & b[322])^(a[215] & b[323])^(a[214] & b[324])^(a[213] & b[325])^(a[212] & b[326])^(a[211] & b[327])^(a[210] & b[328])^(a[209] & b[329])^(a[208] & b[330])^(a[207] & b[331])^(a[206] & b[332])^(a[205] & b[333])^(a[204] & b[334])^(a[203] & b[335])^(a[202] & b[336])^(a[201] & b[337])^(a[200] & b[338])^(a[199] & b[339])^(a[198] & b[340])^(a[197] & b[341])^(a[196] & b[342])^(a[195] & b[343])^(a[194] & b[344])^(a[193] & b[345])^(a[192] & b[346])^(a[191] & b[347])^(a[190] & b[348])^(a[189] & b[349])^(a[188] & b[350])^(a[187] & b[351])^(a[186] & b[352])^(a[185] & b[353])^(a[184] & b[354])^(a[183] & b[355])^(a[182] & b[356])^(a[181] & b[357])^(a[180] & b[358])^(a[179] & b[359])^(a[178] & b[360])^(a[177] & b[361])^(a[176] & b[362])^(a[175] & b[363])^(a[174] & b[364])^(a[173] & b[365])^(a[172] & b[366])^(a[171] & b[367])^(a[170] & b[368])^(a[169] & b[369])^(a[168] & b[370])^(a[167] & b[371])^(a[166] & b[372])^(a[165] & b[373])^(a[164] & b[374])^(a[163] & b[375])^(a[162] & b[376])^(a[161] & b[377])^(a[160] & b[378])^(a[159] & b[379])^(a[158] & b[380])^(a[157] & b[381])^(a[156] & b[382])^(a[155] & b[383])^(a[154] & b[384])^(a[153] & b[385])^(a[152] & b[386])^(a[151] & b[387])^(a[150] & b[388])^(a[149] & b[389])^(a[148] & b[390])^(a[147] & b[391])^(a[146] & b[392])^(a[145] & b[393])^(a[144] & b[394])^(a[143] & b[395])^(a[142] & b[396])^(a[141] & b[397])^(a[140] & b[398])^(a[139] & b[399])^(a[138] & b[400])^(a[137] & b[401])^(a[136] & b[402])^(a[135] & b[403])^(a[134] & b[404])^(a[133] & b[405])^(a[132] & b[406])^(a[131] & b[407])^(a[130] & b[408]);
assign y[539] = (a[408] & b[131])^(a[407] & b[132])^(a[406] & b[133])^(a[405] & b[134])^(a[404] & b[135])^(a[403] & b[136])^(a[402] & b[137])^(a[401] & b[138])^(a[400] & b[139])^(a[399] & b[140])^(a[398] & b[141])^(a[397] & b[142])^(a[396] & b[143])^(a[395] & b[144])^(a[394] & b[145])^(a[393] & b[146])^(a[392] & b[147])^(a[391] & b[148])^(a[390] & b[149])^(a[389] & b[150])^(a[388] & b[151])^(a[387] & b[152])^(a[386] & b[153])^(a[385] & b[154])^(a[384] & b[155])^(a[383] & b[156])^(a[382] & b[157])^(a[381] & b[158])^(a[380] & b[159])^(a[379] & b[160])^(a[378] & b[161])^(a[377] & b[162])^(a[376] & b[163])^(a[375] & b[164])^(a[374] & b[165])^(a[373] & b[166])^(a[372] & b[167])^(a[371] & b[168])^(a[370] & b[169])^(a[369] & b[170])^(a[368] & b[171])^(a[367] & b[172])^(a[366] & b[173])^(a[365] & b[174])^(a[364] & b[175])^(a[363] & b[176])^(a[362] & b[177])^(a[361] & b[178])^(a[360] & b[179])^(a[359] & b[180])^(a[358] & b[181])^(a[357] & b[182])^(a[356] & b[183])^(a[355] & b[184])^(a[354] & b[185])^(a[353] & b[186])^(a[352] & b[187])^(a[351] & b[188])^(a[350] & b[189])^(a[349] & b[190])^(a[348] & b[191])^(a[347] & b[192])^(a[346] & b[193])^(a[345] & b[194])^(a[344] & b[195])^(a[343] & b[196])^(a[342] & b[197])^(a[341] & b[198])^(a[340] & b[199])^(a[339] & b[200])^(a[338] & b[201])^(a[337] & b[202])^(a[336] & b[203])^(a[335] & b[204])^(a[334] & b[205])^(a[333] & b[206])^(a[332] & b[207])^(a[331] & b[208])^(a[330] & b[209])^(a[329] & b[210])^(a[328] & b[211])^(a[327] & b[212])^(a[326] & b[213])^(a[325] & b[214])^(a[324] & b[215])^(a[323] & b[216])^(a[322] & b[217])^(a[321] & b[218])^(a[320] & b[219])^(a[319] & b[220])^(a[318] & b[221])^(a[317] & b[222])^(a[316] & b[223])^(a[315] & b[224])^(a[314] & b[225])^(a[313] & b[226])^(a[312] & b[227])^(a[311] & b[228])^(a[310] & b[229])^(a[309] & b[230])^(a[308] & b[231])^(a[307] & b[232])^(a[306] & b[233])^(a[305] & b[234])^(a[304] & b[235])^(a[303] & b[236])^(a[302] & b[237])^(a[301] & b[238])^(a[300] & b[239])^(a[299] & b[240])^(a[298] & b[241])^(a[297] & b[242])^(a[296] & b[243])^(a[295] & b[244])^(a[294] & b[245])^(a[293] & b[246])^(a[292] & b[247])^(a[291] & b[248])^(a[290] & b[249])^(a[289] & b[250])^(a[288] & b[251])^(a[287] & b[252])^(a[286] & b[253])^(a[285] & b[254])^(a[284] & b[255])^(a[283] & b[256])^(a[282] & b[257])^(a[281] & b[258])^(a[280] & b[259])^(a[279] & b[260])^(a[278] & b[261])^(a[277] & b[262])^(a[276] & b[263])^(a[275] & b[264])^(a[274] & b[265])^(a[273] & b[266])^(a[272] & b[267])^(a[271] & b[268])^(a[270] & b[269])^(a[269] & b[270])^(a[268] & b[271])^(a[267] & b[272])^(a[266] & b[273])^(a[265] & b[274])^(a[264] & b[275])^(a[263] & b[276])^(a[262] & b[277])^(a[261] & b[278])^(a[260] & b[279])^(a[259] & b[280])^(a[258] & b[281])^(a[257] & b[282])^(a[256] & b[283])^(a[255] & b[284])^(a[254] & b[285])^(a[253] & b[286])^(a[252] & b[287])^(a[251] & b[288])^(a[250] & b[289])^(a[249] & b[290])^(a[248] & b[291])^(a[247] & b[292])^(a[246] & b[293])^(a[245] & b[294])^(a[244] & b[295])^(a[243] & b[296])^(a[242] & b[297])^(a[241] & b[298])^(a[240] & b[299])^(a[239] & b[300])^(a[238] & b[301])^(a[237] & b[302])^(a[236] & b[303])^(a[235] & b[304])^(a[234] & b[305])^(a[233] & b[306])^(a[232] & b[307])^(a[231] & b[308])^(a[230] & b[309])^(a[229] & b[310])^(a[228] & b[311])^(a[227] & b[312])^(a[226] & b[313])^(a[225] & b[314])^(a[224] & b[315])^(a[223] & b[316])^(a[222] & b[317])^(a[221] & b[318])^(a[220] & b[319])^(a[219] & b[320])^(a[218] & b[321])^(a[217] & b[322])^(a[216] & b[323])^(a[215] & b[324])^(a[214] & b[325])^(a[213] & b[326])^(a[212] & b[327])^(a[211] & b[328])^(a[210] & b[329])^(a[209] & b[330])^(a[208] & b[331])^(a[207] & b[332])^(a[206] & b[333])^(a[205] & b[334])^(a[204] & b[335])^(a[203] & b[336])^(a[202] & b[337])^(a[201] & b[338])^(a[200] & b[339])^(a[199] & b[340])^(a[198] & b[341])^(a[197] & b[342])^(a[196] & b[343])^(a[195] & b[344])^(a[194] & b[345])^(a[193] & b[346])^(a[192] & b[347])^(a[191] & b[348])^(a[190] & b[349])^(a[189] & b[350])^(a[188] & b[351])^(a[187] & b[352])^(a[186] & b[353])^(a[185] & b[354])^(a[184] & b[355])^(a[183] & b[356])^(a[182] & b[357])^(a[181] & b[358])^(a[180] & b[359])^(a[179] & b[360])^(a[178] & b[361])^(a[177] & b[362])^(a[176] & b[363])^(a[175] & b[364])^(a[174] & b[365])^(a[173] & b[366])^(a[172] & b[367])^(a[171] & b[368])^(a[170] & b[369])^(a[169] & b[370])^(a[168] & b[371])^(a[167] & b[372])^(a[166] & b[373])^(a[165] & b[374])^(a[164] & b[375])^(a[163] & b[376])^(a[162] & b[377])^(a[161] & b[378])^(a[160] & b[379])^(a[159] & b[380])^(a[158] & b[381])^(a[157] & b[382])^(a[156] & b[383])^(a[155] & b[384])^(a[154] & b[385])^(a[153] & b[386])^(a[152] & b[387])^(a[151] & b[388])^(a[150] & b[389])^(a[149] & b[390])^(a[148] & b[391])^(a[147] & b[392])^(a[146] & b[393])^(a[145] & b[394])^(a[144] & b[395])^(a[143] & b[396])^(a[142] & b[397])^(a[141] & b[398])^(a[140] & b[399])^(a[139] & b[400])^(a[138] & b[401])^(a[137] & b[402])^(a[136] & b[403])^(a[135] & b[404])^(a[134] & b[405])^(a[133] & b[406])^(a[132] & b[407])^(a[131] & b[408]);
assign y[540] = (a[408] & b[132])^(a[407] & b[133])^(a[406] & b[134])^(a[405] & b[135])^(a[404] & b[136])^(a[403] & b[137])^(a[402] & b[138])^(a[401] & b[139])^(a[400] & b[140])^(a[399] & b[141])^(a[398] & b[142])^(a[397] & b[143])^(a[396] & b[144])^(a[395] & b[145])^(a[394] & b[146])^(a[393] & b[147])^(a[392] & b[148])^(a[391] & b[149])^(a[390] & b[150])^(a[389] & b[151])^(a[388] & b[152])^(a[387] & b[153])^(a[386] & b[154])^(a[385] & b[155])^(a[384] & b[156])^(a[383] & b[157])^(a[382] & b[158])^(a[381] & b[159])^(a[380] & b[160])^(a[379] & b[161])^(a[378] & b[162])^(a[377] & b[163])^(a[376] & b[164])^(a[375] & b[165])^(a[374] & b[166])^(a[373] & b[167])^(a[372] & b[168])^(a[371] & b[169])^(a[370] & b[170])^(a[369] & b[171])^(a[368] & b[172])^(a[367] & b[173])^(a[366] & b[174])^(a[365] & b[175])^(a[364] & b[176])^(a[363] & b[177])^(a[362] & b[178])^(a[361] & b[179])^(a[360] & b[180])^(a[359] & b[181])^(a[358] & b[182])^(a[357] & b[183])^(a[356] & b[184])^(a[355] & b[185])^(a[354] & b[186])^(a[353] & b[187])^(a[352] & b[188])^(a[351] & b[189])^(a[350] & b[190])^(a[349] & b[191])^(a[348] & b[192])^(a[347] & b[193])^(a[346] & b[194])^(a[345] & b[195])^(a[344] & b[196])^(a[343] & b[197])^(a[342] & b[198])^(a[341] & b[199])^(a[340] & b[200])^(a[339] & b[201])^(a[338] & b[202])^(a[337] & b[203])^(a[336] & b[204])^(a[335] & b[205])^(a[334] & b[206])^(a[333] & b[207])^(a[332] & b[208])^(a[331] & b[209])^(a[330] & b[210])^(a[329] & b[211])^(a[328] & b[212])^(a[327] & b[213])^(a[326] & b[214])^(a[325] & b[215])^(a[324] & b[216])^(a[323] & b[217])^(a[322] & b[218])^(a[321] & b[219])^(a[320] & b[220])^(a[319] & b[221])^(a[318] & b[222])^(a[317] & b[223])^(a[316] & b[224])^(a[315] & b[225])^(a[314] & b[226])^(a[313] & b[227])^(a[312] & b[228])^(a[311] & b[229])^(a[310] & b[230])^(a[309] & b[231])^(a[308] & b[232])^(a[307] & b[233])^(a[306] & b[234])^(a[305] & b[235])^(a[304] & b[236])^(a[303] & b[237])^(a[302] & b[238])^(a[301] & b[239])^(a[300] & b[240])^(a[299] & b[241])^(a[298] & b[242])^(a[297] & b[243])^(a[296] & b[244])^(a[295] & b[245])^(a[294] & b[246])^(a[293] & b[247])^(a[292] & b[248])^(a[291] & b[249])^(a[290] & b[250])^(a[289] & b[251])^(a[288] & b[252])^(a[287] & b[253])^(a[286] & b[254])^(a[285] & b[255])^(a[284] & b[256])^(a[283] & b[257])^(a[282] & b[258])^(a[281] & b[259])^(a[280] & b[260])^(a[279] & b[261])^(a[278] & b[262])^(a[277] & b[263])^(a[276] & b[264])^(a[275] & b[265])^(a[274] & b[266])^(a[273] & b[267])^(a[272] & b[268])^(a[271] & b[269])^(a[270] & b[270])^(a[269] & b[271])^(a[268] & b[272])^(a[267] & b[273])^(a[266] & b[274])^(a[265] & b[275])^(a[264] & b[276])^(a[263] & b[277])^(a[262] & b[278])^(a[261] & b[279])^(a[260] & b[280])^(a[259] & b[281])^(a[258] & b[282])^(a[257] & b[283])^(a[256] & b[284])^(a[255] & b[285])^(a[254] & b[286])^(a[253] & b[287])^(a[252] & b[288])^(a[251] & b[289])^(a[250] & b[290])^(a[249] & b[291])^(a[248] & b[292])^(a[247] & b[293])^(a[246] & b[294])^(a[245] & b[295])^(a[244] & b[296])^(a[243] & b[297])^(a[242] & b[298])^(a[241] & b[299])^(a[240] & b[300])^(a[239] & b[301])^(a[238] & b[302])^(a[237] & b[303])^(a[236] & b[304])^(a[235] & b[305])^(a[234] & b[306])^(a[233] & b[307])^(a[232] & b[308])^(a[231] & b[309])^(a[230] & b[310])^(a[229] & b[311])^(a[228] & b[312])^(a[227] & b[313])^(a[226] & b[314])^(a[225] & b[315])^(a[224] & b[316])^(a[223] & b[317])^(a[222] & b[318])^(a[221] & b[319])^(a[220] & b[320])^(a[219] & b[321])^(a[218] & b[322])^(a[217] & b[323])^(a[216] & b[324])^(a[215] & b[325])^(a[214] & b[326])^(a[213] & b[327])^(a[212] & b[328])^(a[211] & b[329])^(a[210] & b[330])^(a[209] & b[331])^(a[208] & b[332])^(a[207] & b[333])^(a[206] & b[334])^(a[205] & b[335])^(a[204] & b[336])^(a[203] & b[337])^(a[202] & b[338])^(a[201] & b[339])^(a[200] & b[340])^(a[199] & b[341])^(a[198] & b[342])^(a[197] & b[343])^(a[196] & b[344])^(a[195] & b[345])^(a[194] & b[346])^(a[193] & b[347])^(a[192] & b[348])^(a[191] & b[349])^(a[190] & b[350])^(a[189] & b[351])^(a[188] & b[352])^(a[187] & b[353])^(a[186] & b[354])^(a[185] & b[355])^(a[184] & b[356])^(a[183] & b[357])^(a[182] & b[358])^(a[181] & b[359])^(a[180] & b[360])^(a[179] & b[361])^(a[178] & b[362])^(a[177] & b[363])^(a[176] & b[364])^(a[175] & b[365])^(a[174] & b[366])^(a[173] & b[367])^(a[172] & b[368])^(a[171] & b[369])^(a[170] & b[370])^(a[169] & b[371])^(a[168] & b[372])^(a[167] & b[373])^(a[166] & b[374])^(a[165] & b[375])^(a[164] & b[376])^(a[163] & b[377])^(a[162] & b[378])^(a[161] & b[379])^(a[160] & b[380])^(a[159] & b[381])^(a[158] & b[382])^(a[157] & b[383])^(a[156] & b[384])^(a[155] & b[385])^(a[154] & b[386])^(a[153] & b[387])^(a[152] & b[388])^(a[151] & b[389])^(a[150] & b[390])^(a[149] & b[391])^(a[148] & b[392])^(a[147] & b[393])^(a[146] & b[394])^(a[145] & b[395])^(a[144] & b[396])^(a[143] & b[397])^(a[142] & b[398])^(a[141] & b[399])^(a[140] & b[400])^(a[139] & b[401])^(a[138] & b[402])^(a[137] & b[403])^(a[136] & b[404])^(a[135] & b[405])^(a[134] & b[406])^(a[133] & b[407])^(a[132] & b[408]);
assign y[541] = (a[408] & b[133])^(a[407] & b[134])^(a[406] & b[135])^(a[405] & b[136])^(a[404] & b[137])^(a[403] & b[138])^(a[402] & b[139])^(a[401] & b[140])^(a[400] & b[141])^(a[399] & b[142])^(a[398] & b[143])^(a[397] & b[144])^(a[396] & b[145])^(a[395] & b[146])^(a[394] & b[147])^(a[393] & b[148])^(a[392] & b[149])^(a[391] & b[150])^(a[390] & b[151])^(a[389] & b[152])^(a[388] & b[153])^(a[387] & b[154])^(a[386] & b[155])^(a[385] & b[156])^(a[384] & b[157])^(a[383] & b[158])^(a[382] & b[159])^(a[381] & b[160])^(a[380] & b[161])^(a[379] & b[162])^(a[378] & b[163])^(a[377] & b[164])^(a[376] & b[165])^(a[375] & b[166])^(a[374] & b[167])^(a[373] & b[168])^(a[372] & b[169])^(a[371] & b[170])^(a[370] & b[171])^(a[369] & b[172])^(a[368] & b[173])^(a[367] & b[174])^(a[366] & b[175])^(a[365] & b[176])^(a[364] & b[177])^(a[363] & b[178])^(a[362] & b[179])^(a[361] & b[180])^(a[360] & b[181])^(a[359] & b[182])^(a[358] & b[183])^(a[357] & b[184])^(a[356] & b[185])^(a[355] & b[186])^(a[354] & b[187])^(a[353] & b[188])^(a[352] & b[189])^(a[351] & b[190])^(a[350] & b[191])^(a[349] & b[192])^(a[348] & b[193])^(a[347] & b[194])^(a[346] & b[195])^(a[345] & b[196])^(a[344] & b[197])^(a[343] & b[198])^(a[342] & b[199])^(a[341] & b[200])^(a[340] & b[201])^(a[339] & b[202])^(a[338] & b[203])^(a[337] & b[204])^(a[336] & b[205])^(a[335] & b[206])^(a[334] & b[207])^(a[333] & b[208])^(a[332] & b[209])^(a[331] & b[210])^(a[330] & b[211])^(a[329] & b[212])^(a[328] & b[213])^(a[327] & b[214])^(a[326] & b[215])^(a[325] & b[216])^(a[324] & b[217])^(a[323] & b[218])^(a[322] & b[219])^(a[321] & b[220])^(a[320] & b[221])^(a[319] & b[222])^(a[318] & b[223])^(a[317] & b[224])^(a[316] & b[225])^(a[315] & b[226])^(a[314] & b[227])^(a[313] & b[228])^(a[312] & b[229])^(a[311] & b[230])^(a[310] & b[231])^(a[309] & b[232])^(a[308] & b[233])^(a[307] & b[234])^(a[306] & b[235])^(a[305] & b[236])^(a[304] & b[237])^(a[303] & b[238])^(a[302] & b[239])^(a[301] & b[240])^(a[300] & b[241])^(a[299] & b[242])^(a[298] & b[243])^(a[297] & b[244])^(a[296] & b[245])^(a[295] & b[246])^(a[294] & b[247])^(a[293] & b[248])^(a[292] & b[249])^(a[291] & b[250])^(a[290] & b[251])^(a[289] & b[252])^(a[288] & b[253])^(a[287] & b[254])^(a[286] & b[255])^(a[285] & b[256])^(a[284] & b[257])^(a[283] & b[258])^(a[282] & b[259])^(a[281] & b[260])^(a[280] & b[261])^(a[279] & b[262])^(a[278] & b[263])^(a[277] & b[264])^(a[276] & b[265])^(a[275] & b[266])^(a[274] & b[267])^(a[273] & b[268])^(a[272] & b[269])^(a[271] & b[270])^(a[270] & b[271])^(a[269] & b[272])^(a[268] & b[273])^(a[267] & b[274])^(a[266] & b[275])^(a[265] & b[276])^(a[264] & b[277])^(a[263] & b[278])^(a[262] & b[279])^(a[261] & b[280])^(a[260] & b[281])^(a[259] & b[282])^(a[258] & b[283])^(a[257] & b[284])^(a[256] & b[285])^(a[255] & b[286])^(a[254] & b[287])^(a[253] & b[288])^(a[252] & b[289])^(a[251] & b[290])^(a[250] & b[291])^(a[249] & b[292])^(a[248] & b[293])^(a[247] & b[294])^(a[246] & b[295])^(a[245] & b[296])^(a[244] & b[297])^(a[243] & b[298])^(a[242] & b[299])^(a[241] & b[300])^(a[240] & b[301])^(a[239] & b[302])^(a[238] & b[303])^(a[237] & b[304])^(a[236] & b[305])^(a[235] & b[306])^(a[234] & b[307])^(a[233] & b[308])^(a[232] & b[309])^(a[231] & b[310])^(a[230] & b[311])^(a[229] & b[312])^(a[228] & b[313])^(a[227] & b[314])^(a[226] & b[315])^(a[225] & b[316])^(a[224] & b[317])^(a[223] & b[318])^(a[222] & b[319])^(a[221] & b[320])^(a[220] & b[321])^(a[219] & b[322])^(a[218] & b[323])^(a[217] & b[324])^(a[216] & b[325])^(a[215] & b[326])^(a[214] & b[327])^(a[213] & b[328])^(a[212] & b[329])^(a[211] & b[330])^(a[210] & b[331])^(a[209] & b[332])^(a[208] & b[333])^(a[207] & b[334])^(a[206] & b[335])^(a[205] & b[336])^(a[204] & b[337])^(a[203] & b[338])^(a[202] & b[339])^(a[201] & b[340])^(a[200] & b[341])^(a[199] & b[342])^(a[198] & b[343])^(a[197] & b[344])^(a[196] & b[345])^(a[195] & b[346])^(a[194] & b[347])^(a[193] & b[348])^(a[192] & b[349])^(a[191] & b[350])^(a[190] & b[351])^(a[189] & b[352])^(a[188] & b[353])^(a[187] & b[354])^(a[186] & b[355])^(a[185] & b[356])^(a[184] & b[357])^(a[183] & b[358])^(a[182] & b[359])^(a[181] & b[360])^(a[180] & b[361])^(a[179] & b[362])^(a[178] & b[363])^(a[177] & b[364])^(a[176] & b[365])^(a[175] & b[366])^(a[174] & b[367])^(a[173] & b[368])^(a[172] & b[369])^(a[171] & b[370])^(a[170] & b[371])^(a[169] & b[372])^(a[168] & b[373])^(a[167] & b[374])^(a[166] & b[375])^(a[165] & b[376])^(a[164] & b[377])^(a[163] & b[378])^(a[162] & b[379])^(a[161] & b[380])^(a[160] & b[381])^(a[159] & b[382])^(a[158] & b[383])^(a[157] & b[384])^(a[156] & b[385])^(a[155] & b[386])^(a[154] & b[387])^(a[153] & b[388])^(a[152] & b[389])^(a[151] & b[390])^(a[150] & b[391])^(a[149] & b[392])^(a[148] & b[393])^(a[147] & b[394])^(a[146] & b[395])^(a[145] & b[396])^(a[144] & b[397])^(a[143] & b[398])^(a[142] & b[399])^(a[141] & b[400])^(a[140] & b[401])^(a[139] & b[402])^(a[138] & b[403])^(a[137] & b[404])^(a[136] & b[405])^(a[135] & b[406])^(a[134] & b[407])^(a[133] & b[408]);
assign y[542] = (a[408] & b[134])^(a[407] & b[135])^(a[406] & b[136])^(a[405] & b[137])^(a[404] & b[138])^(a[403] & b[139])^(a[402] & b[140])^(a[401] & b[141])^(a[400] & b[142])^(a[399] & b[143])^(a[398] & b[144])^(a[397] & b[145])^(a[396] & b[146])^(a[395] & b[147])^(a[394] & b[148])^(a[393] & b[149])^(a[392] & b[150])^(a[391] & b[151])^(a[390] & b[152])^(a[389] & b[153])^(a[388] & b[154])^(a[387] & b[155])^(a[386] & b[156])^(a[385] & b[157])^(a[384] & b[158])^(a[383] & b[159])^(a[382] & b[160])^(a[381] & b[161])^(a[380] & b[162])^(a[379] & b[163])^(a[378] & b[164])^(a[377] & b[165])^(a[376] & b[166])^(a[375] & b[167])^(a[374] & b[168])^(a[373] & b[169])^(a[372] & b[170])^(a[371] & b[171])^(a[370] & b[172])^(a[369] & b[173])^(a[368] & b[174])^(a[367] & b[175])^(a[366] & b[176])^(a[365] & b[177])^(a[364] & b[178])^(a[363] & b[179])^(a[362] & b[180])^(a[361] & b[181])^(a[360] & b[182])^(a[359] & b[183])^(a[358] & b[184])^(a[357] & b[185])^(a[356] & b[186])^(a[355] & b[187])^(a[354] & b[188])^(a[353] & b[189])^(a[352] & b[190])^(a[351] & b[191])^(a[350] & b[192])^(a[349] & b[193])^(a[348] & b[194])^(a[347] & b[195])^(a[346] & b[196])^(a[345] & b[197])^(a[344] & b[198])^(a[343] & b[199])^(a[342] & b[200])^(a[341] & b[201])^(a[340] & b[202])^(a[339] & b[203])^(a[338] & b[204])^(a[337] & b[205])^(a[336] & b[206])^(a[335] & b[207])^(a[334] & b[208])^(a[333] & b[209])^(a[332] & b[210])^(a[331] & b[211])^(a[330] & b[212])^(a[329] & b[213])^(a[328] & b[214])^(a[327] & b[215])^(a[326] & b[216])^(a[325] & b[217])^(a[324] & b[218])^(a[323] & b[219])^(a[322] & b[220])^(a[321] & b[221])^(a[320] & b[222])^(a[319] & b[223])^(a[318] & b[224])^(a[317] & b[225])^(a[316] & b[226])^(a[315] & b[227])^(a[314] & b[228])^(a[313] & b[229])^(a[312] & b[230])^(a[311] & b[231])^(a[310] & b[232])^(a[309] & b[233])^(a[308] & b[234])^(a[307] & b[235])^(a[306] & b[236])^(a[305] & b[237])^(a[304] & b[238])^(a[303] & b[239])^(a[302] & b[240])^(a[301] & b[241])^(a[300] & b[242])^(a[299] & b[243])^(a[298] & b[244])^(a[297] & b[245])^(a[296] & b[246])^(a[295] & b[247])^(a[294] & b[248])^(a[293] & b[249])^(a[292] & b[250])^(a[291] & b[251])^(a[290] & b[252])^(a[289] & b[253])^(a[288] & b[254])^(a[287] & b[255])^(a[286] & b[256])^(a[285] & b[257])^(a[284] & b[258])^(a[283] & b[259])^(a[282] & b[260])^(a[281] & b[261])^(a[280] & b[262])^(a[279] & b[263])^(a[278] & b[264])^(a[277] & b[265])^(a[276] & b[266])^(a[275] & b[267])^(a[274] & b[268])^(a[273] & b[269])^(a[272] & b[270])^(a[271] & b[271])^(a[270] & b[272])^(a[269] & b[273])^(a[268] & b[274])^(a[267] & b[275])^(a[266] & b[276])^(a[265] & b[277])^(a[264] & b[278])^(a[263] & b[279])^(a[262] & b[280])^(a[261] & b[281])^(a[260] & b[282])^(a[259] & b[283])^(a[258] & b[284])^(a[257] & b[285])^(a[256] & b[286])^(a[255] & b[287])^(a[254] & b[288])^(a[253] & b[289])^(a[252] & b[290])^(a[251] & b[291])^(a[250] & b[292])^(a[249] & b[293])^(a[248] & b[294])^(a[247] & b[295])^(a[246] & b[296])^(a[245] & b[297])^(a[244] & b[298])^(a[243] & b[299])^(a[242] & b[300])^(a[241] & b[301])^(a[240] & b[302])^(a[239] & b[303])^(a[238] & b[304])^(a[237] & b[305])^(a[236] & b[306])^(a[235] & b[307])^(a[234] & b[308])^(a[233] & b[309])^(a[232] & b[310])^(a[231] & b[311])^(a[230] & b[312])^(a[229] & b[313])^(a[228] & b[314])^(a[227] & b[315])^(a[226] & b[316])^(a[225] & b[317])^(a[224] & b[318])^(a[223] & b[319])^(a[222] & b[320])^(a[221] & b[321])^(a[220] & b[322])^(a[219] & b[323])^(a[218] & b[324])^(a[217] & b[325])^(a[216] & b[326])^(a[215] & b[327])^(a[214] & b[328])^(a[213] & b[329])^(a[212] & b[330])^(a[211] & b[331])^(a[210] & b[332])^(a[209] & b[333])^(a[208] & b[334])^(a[207] & b[335])^(a[206] & b[336])^(a[205] & b[337])^(a[204] & b[338])^(a[203] & b[339])^(a[202] & b[340])^(a[201] & b[341])^(a[200] & b[342])^(a[199] & b[343])^(a[198] & b[344])^(a[197] & b[345])^(a[196] & b[346])^(a[195] & b[347])^(a[194] & b[348])^(a[193] & b[349])^(a[192] & b[350])^(a[191] & b[351])^(a[190] & b[352])^(a[189] & b[353])^(a[188] & b[354])^(a[187] & b[355])^(a[186] & b[356])^(a[185] & b[357])^(a[184] & b[358])^(a[183] & b[359])^(a[182] & b[360])^(a[181] & b[361])^(a[180] & b[362])^(a[179] & b[363])^(a[178] & b[364])^(a[177] & b[365])^(a[176] & b[366])^(a[175] & b[367])^(a[174] & b[368])^(a[173] & b[369])^(a[172] & b[370])^(a[171] & b[371])^(a[170] & b[372])^(a[169] & b[373])^(a[168] & b[374])^(a[167] & b[375])^(a[166] & b[376])^(a[165] & b[377])^(a[164] & b[378])^(a[163] & b[379])^(a[162] & b[380])^(a[161] & b[381])^(a[160] & b[382])^(a[159] & b[383])^(a[158] & b[384])^(a[157] & b[385])^(a[156] & b[386])^(a[155] & b[387])^(a[154] & b[388])^(a[153] & b[389])^(a[152] & b[390])^(a[151] & b[391])^(a[150] & b[392])^(a[149] & b[393])^(a[148] & b[394])^(a[147] & b[395])^(a[146] & b[396])^(a[145] & b[397])^(a[144] & b[398])^(a[143] & b[399])^(a[142] & b[400])^(a[141] & b[401])^(a[140] & b[402])^(a[139] & b[403])^(a[138] & b[404])^(a[137] & b[405])^(a[136] & b[406])^(a[135] & b[407])^(a[134] & b[408]);
assign y[543] = (a[408] & b[135])^(a[407] & b[136])^(a[406] & b[137])^(a[405] & b[138])^(a[404] & b[139])^(a[403] & b[140])^(a[402] & b[141])^(a[401] & b[142])^(a[400] & b[143])^(a[399] & b[144])^(a[398] & b[145])^(a[397] & b[146])^(a[396] & b[147])^(a[395] & b[148])^(a[394] & b[149])^(a[393] & b[150])^(a[392] & b[151])^(a[391] & b[152])^(a[390] & b[153])^(a[389] & b[154])^(a[388] & b[155])^(a[387] & b[156])^(a[386] & b[157])^(a[385] & b[158])^(a[384] & b[159])^(a[383] & b[160])^(a[382] & b[161])^(a[381] & b[162])^(a[380] & b[163])^(a[379] & b[164])^(a[378] & b[165])^(a[377] & b[166])^(a[376] & b[167])^(a[375] & b[168])^(a[374] & b[169])^(a[373] & b[170])^(a[372] & b[171])^(a[371] & b[172])^(a[370] & b[173])^(a[369] & b[174])^(a[368] & b[175])^(a[367] & b[176])^(a[366] & b[177])^(a[365] & b[178])^(a[364] & b[179])^(a[363] & b[180])^(a[362] & b[181])^(a[361] & b[182])^(a[360] & b[183])^(a[359] & b[184])^(a[358] & b[185])^(a[357] & b[186])^(a[356] & b[187])^(a[355] & b[188])^(a[354] & b[189])^(a[353] & b[190])^(a[352] & b[191])^(a[351] & b[192])^(a[350] & b[193])^(a[349] & b[194])^(a[348] & b[195])^(a[347] & b[196])^(a[346] & b[197])^(a[345] & b[198])^(a[344] & b[199])^(a[343] & b[200])^(a[342] & b[201])^(a[341] & b[202])^(a[340] & b[203])^(a[339] & b[204])^(a[338] & b[205])^(a[337] & b[206])^(a[336] & b[207])^(a[335] & b[208])^(a[334] & b[209])^(a[333] & b[210])^(a[332] & b[211])^(a[331] & b[212])^(a[330] & b[213])^(a[329] & b[214])^(a[328] & b[215])^(a[327] & b[216])^(a[326] & b[217])^(a[325] & b[218])^(a[324] & b[219])^(a[323] & b[220])^(a[322] & b[221])^(a[321] & b[222])^(a[320] & b[223])^(a[319] & b[224])^(a[318] & b[225])^(a[317] & b[226])^(a[316] & b[227])^(a[315] & b[228])^(a[314] & b[229])^(a[313] & b[230])^(a[312] & b[231])^(a[311] & b[232])^(a[310] & b[233])^(a[309] & b[234])^(a[308] & b[235])^(a[307] & b[236])^(a[306] & b[237])^(a[305] & b[238])^(a[304] & b[239])^(a[303] & b[240])^(a[302] & b[241])^(a[301] & b[242])^(a[300] & b[243])^(a[299] & b[244])^(a[298] & b[245])^(a[297] & b[246])^(a[296] & b[247])^(a[295] & b[248])^(a[294] & b[249])^(a[293] & b[250])^(a[292] & b[251])^(a[291] & b[252])^(a[290] & b[253])^(a[289] & b[254])^(a[288] & b[255])^(a[287] & b[256])^(a[286] & b[257])^(a[285] & b[258])^(a[284] & b[259])^(a[283] & b[260])^(a[282] & b[261])^(a[281] & b[262])^(a[280] & b[263])^(a[279] & b[264])^(a[278] & b[265])^(a[277] & b[266])^(a[276] & b[267])^(a[275] & b[268])^(a[274] & b[269])^(a[273] & b[270])^(a[272] & b[271])^(a[271] & b[272])^(a[270] & b[273])^(a[269] & b[274])^(a[268] & b[275])^(a[267] & b[276])^(a[266] & b[277])^(a[265] & b[278])^(a[264] & b[279])^(a[263] & b[280])^(a[262] & b[281])^(a[261] & b[282])^(a[260] & b[283])^(a[259] & b[284])^(a[258] & b[285])^(a[257] & b[286])^(a[256] & b[287])^(a[255] & b[288])^(a[254] & b[289])^(a[253] & b[290])^(a[252] & b[291])^(a[251] & b[292])^(a[250] & b[293])^(a[249] & b[294])^(a[248] & b[295])^(a[247] & b[296])^(a[246] & b[297])^(a[245] & b[298])^(a[244] & b[299])^(a[243] & b[300])^(a[242] & b[301])^(a[241] & b[302])^(a[240] & b[303])^(a[239] & b[304])^(a[238] & b[305])^(a[237] & b[306])^(a[236] & b[307])^(a[235] & b[308])^(a[234] & b[309])^(a[233] & b[310])^(a[232] & b[311])^(a[231] & b[312])^(a[230] & b[313])^(a[229] & b[314])^(a[228] & b[315])^(a[227] & b[316])^(a[226] & b[317])^(a[225] & b[318])^(a[224] & b[319])^(a[223] & b[320])^(a[222] & b[321])^(a[221] & b[322])^(a[220] & b[323])^(a[219] & b[324])^(a[218] & b[325])^(a[217] & b[326])^(a[216] & b[327])^(a[215] & b[328])^(a[214] & b[329])^(a[213] & b[330])^(a[212] & b[331])^(a[211] & b[332])^(a[210] & b[333])^(a[209] & b[334])^(a[208] & b[335])^(a[207] & b[336])^(a[206] & b[337])^(a[205] & b[338])^(a[204] & b[339])^(a[203] & b[340])^(a[202] & b[341])^(a[201] & b[342])^(a[200] & b[343])^(a[199] & b[344])^(a[198] & b[345])^(a[197] & b[346])^(a[196] & b[347])^(a[195] & b[348])^(a[194] & b[349])^(a[193] & b[350])^(a[192] & b[351])^(a[191] & b[352])^(a[190] & b[353])^(a[189] & b[354])^(a[188] & b[355])^(a[187] & b[356])^(a[186] & b[357])^(a[185] & b[358])^(a[184] & b[359])^(a[183] & b[360])^(a[182] & b[361])^(a[181] & b[362])^(a[180] & b[363])^(a[179] & b[364])^(a[178] & b[365])^(a[177] & b[366])^(a[176] & b[367])^(a[175] & b[368])^(a[174] & b[369])^(a[173] & b[370])^(a[172] & b[371])^(a[171] & b[372])^(a[170] & b[373])^(a[169] & b[374])^(a[168] & b[375])^(a[167] & b[376])^(a[166] & b[377])^(a[165] & b[378])^(a[164] & b[379])^(a[163] & b[380])^(a[162] & b[381])^(a[161] & b[382])^(a[160] & b[383])^(a[159] & b[384])^(a[158] & b[385])^(a[157] & b[386])^(a[156] & b[387])^(a[155] & b[388])^(a[154] & b[389])^(a[153] & b[390])^(a[152] & b[391])^(a[151] & b[392])^(a[150] & b[393])^(a[149] & b[394])^(a[148] & b[395])^(a[147] & b[396])^(a[146] & b[397])^(a[145] & b[398])^(a[144] & b[399])^(a[143] & b[400])^(a[142] & b[401])^(a[141] & b[402])^(a[140] & b[403])^(a[139] & b[404])^(a[138] & b[405])^(a[137] & b[406])^(a[136] & b[407])^(a[135] & b[408]);
assign y[544] = (a[408] & b[136])^(a[407] & b[137])^(a[406] & b[138])^(a[405] & b[139])^(a[404] & b[140])^(a[403] & b[141])^(a[402] & b[142])^(a[401] & b[143])^(a[400] & b[144])^(a[399] & b[145])^(a[398] & b[146])^(a[397] & b[147])^(a[396] & b[148])^(a[395] & b[149])^(a[394] & b[150])^(a[393] & b[151])^(a[392] & b[152])^(a[391] & b[153])^(a[390] & b[154])^(a[389] & b[155])^(a[388] & b[156])^(a[387] & b[157])^(a[386] & b[158])^(a[385] & b[159])^(a[384] & b[160])^(a[383] & b[161])^(a[382] & b[162])^(a[381] & b[163])^(a[380] & b[164])^(a[379] & b[165])^(a[378] & b[166])^(a[377] & b[167])^(a[376] & b[168])^(a[375] & b[169])^(a[374] & b[170])^(a[373] & b[171])^(a[372] & b[172])^(a[371] & b[173])^(a[370] & b[174])^(a[369] & b[175])^(a[368] & b[176])^(a[367] & b[177])^(a[366] & b[178])^(a[365] & b[179])^(a[364] & b[180])^(a[363] & b[181])^(a[362] & b[182])^(a[361] & b[183])^(a[360] & b[184])^(a[359] & b[185])^(a[358] & b[186])^(a[357] & b[187])^(a[356] & b[188])^(a[355] & b[189])^(a[354] & b[190])^(a[353] & b[191])^(a[352] & b[192])^(a[351] & b[193])^(a[350] & b[194])^(a[349] & b[195])^(a[348] & b[196])^(a[347] & b[197])^(a[346] & b[198])^(a[345] & b[199])^(a[344] & b[200])^(a[343] & b[201])^(a[342] & b[202])^(a[341] & b[203])^(a[340] & b[204])^(a[339] & b[205])^(a[338] & b[206])^(a[337] & b[207])^(a[336] & b[208])^(a[335] & b[209])^(a[334] & b[210])^(a[333] & b[211])^(a[332] & b[212])^(a[331] & b[213])^(a[330] & b[214])^(a[329] & b[215])^(a[328] & b[216])^(a[327] & b[217])^(a[326] & b[218])^(a[325] & b[219])^(a[324] & b[220])^(a[323] & b[221])^(a[322] & b[222])^(a[321] & b[223])^(a[320] & b[224])^(a[319] & b[225])^(a[318] & b[226])^(a[317] & b[227])^(a[316] & b[228])^(a[315] & b[229])^(a[314] & b[230])^(a[313] & b[231])^(a[312] & b[232])^(a[311] & b[233])^(a[310] & b[234])^(a[309] & b[235])^(a[308] & b[236])^(a[307] & b[237])^(a[306] & b[238])^(a[305] & b[239])^(a[304] & b[240])^(a[303] & b[241])^(a[302] & b[242])^(a[301] & b[243])^(a[300] & b[244])^(a[299] & b[245])^(a[298] & b[246])^(a[297] & b[247])^(a[296] & b[248])^(a[295] & b[249])^(a[294] & b[250])^(a[293] & b[251])^(a[292] & b[252])^(a[291] & b[253])^(a[290] & b[254])^(a[289] & b[255])^(a[288] & b[256])^(a[287] & b[257])^(a[286] & b[258])^(a[285] & b[259])^(a[284] & b[260])^(a[283] & b[261])^(a[282] & b[262])^(a[281] & b[263])^(a[280] & b[264])^(a[279] & b[265])^(a[278] & b[266])^(a[277] & b[267])^(a[276] & b[268])^(a[275] & b[269])^(a[274] & b[270])^(a[273] & b[271])^(a[272] & b[272])^(a[271] & b[273])^(a[270] & b[274])^(a[269] & b[275])^(a[268] & b[276])^(a[267] & b[277])^(a[266] & b[278])^(a[265] & b[279])^(a[264] & b[280])^(a[263] & b[281])^(a[262] & b[282])^(a[261] & b[283])^(a[260] & b[284])^(a[259] & b[285])^(a[258] & b[286])^(a[257] & b[287])^(a[256] & b[288])^(a[255] & b[289])^(a[254] & b[290])^(a[253] & b[291])^(a[252] & b[292])^(a[251] & b[293])^(a[250] & b[294])^(a[249] & b[295])^(a[248] & b[296])^(a[247] & b[297])^(a[246] & b[298])^(a[245] & b[299])^(a[244] & b[300])^(a[243] & b[301])^(a[242] & b[302])^(a[241] & b[303])^(a[240] & b[304])^(a[239] & b[305])^(a[238] & b[306])^(a[237] & b[307])^(a[236] & b[308])^(a[235] & b[309])^(a[234] & b[310])^(a[233] & b[311])^(a[232] & b[312])^(a[231] & b[313])^(a[230] & b[314])^(a[229] & b[315])^(a[228] & b[316])^(a[227] & b[317])^(a[226] & b[318])^(a[225] & b[319])^(a[224] & b[320])^(a[223] & b[321])^(a[222] & b[322])^(a[221] & b[323])^(a[220] & b[324])^(a[219] & b[325])^(a[218] & b[326])^(a[217] & b[327])^(a[216] & b[328])^(a[215] & b[329])^(a[214] & b[330])^(a[213] & b[331])^(a[212] & b[332])^(a[211] & b[333])^(a[210] & b[334])^(a[209] & b[335])^(a[208] & b[336])^(a[207] & b[337])^(a[206] & b[338])^(a[205] & b[339])^(a[204] & b[340])^(a[203] & b[341])^(a[202] & b[342])^(a[201] & b[343])^(a[200] & b[344])^(a[199] & b[345])^(a[198] & b[346])^(a[197] & b[347])^(a[196] & b[348])^(a[195] & b[349])^(a[194] & b[350])^(a[193] & b[351])^(a[192] & b[352])^(a[191] & b[353])^(a[190] & b[354])^(a[189] & b[355])^(a[188] & b[356])^(a[187] & b[357])^(a[186] & b[358])^(a[185] & b[359])^(a[184] & b[360])^(a[183] & b[361])^(a[182] & b[362])^(a[181] & b[363])^(a[180] & b[364])^(a[179] & b[365])^(a[178] & b[366])^(a[177] & b[367])^(a[176] & b[368])^(a[175] & b[369])^(a[174] & b[370])^(a[173] & b[371])^(a[172] & b[372])^(a[171] & b[373])^(a[170] & b[374])^(a[169] & b[375])^(a[168] & b[376])^(a[167] & b[377])^(a[166] & b[378])^(a[165] & b[379])^(a[164] & b[380])^(a[163] & b[381])^(a[162] & b[382])^(a[161] & b[383])^(a[160] & b[384])^(a[159] & b[385])^(a[158] & b[386])^(a[157] & b[387])^(a[156] & b[388])^(a[155] & b[389])^(a[154] & b[390])^(a[153] & b[391])^(a[152] & b[392])^(a[151] & b[393])^(a[150] & b[394])^(a[149] & b[395])^(a[148] & b[396])^(a[147] & b[397])^(a[146] & b[398])^(a[145] & b[399])^(a[144] & b[400])^(a[143] & b[401])^(a[142] & b[402])^(a[141] & b[403])^(a[140] & b[404])^(a[139] & b[405])^(a[138] & b[406])^(a[137] & b[407])^(a[136] & b[408]);
assign y[545] = (a[408] & b[137])^(a[407] & b[138])^(a[406] & b[139])^(a[405] & b[140])^(a[404] & b[141])^(a[403] & b[142])^(a[402] & b[143])^(a[401] & b[144])^(a[400] & b[145])^(a[399] & b[146])^(a[398] & b[147])^(a[397] & b[148])^(a[396] & b[149])^(a[395] & b[150])^(a[394] & b[151])^(a[393] & b[152])^(a[392] & b[153])^(a[391] & b[154])^(a[390] & b[155])^(a[389] & b[156])^(a[388] & b[157])^(a[387] & b[158])^(a[386] & b[159])^(a[385] & b[160])^(a[384] & b[161])^(a[383] & b[162])^(a[382] & b[163])^(a[381] & b[164])^(a[380] & b[165])^(a[379] & b[166])^(a[378] & b[167])^(a[377] & b[168])^(a[376] & b[169])^(a[375] & b[170])^(a[374] & b[171])^(a[373] & b[172])^(a[372] & b[173])^(a[371] & b[174])^(a[370] & b[175])^(a[369] & b[176])^(a[368] & b[177])^(a[367] & b[178])^(a[366] & b[179])^(a[365] & b[180])^(a[364] & b[181])^(a[363] & b[182])^(a[362] & b[183])^(a[361] & b[184])^(a[360] & b[185])^(a[359] & b[186])^(a[358] & b[187])^(a[357] & b[188])^(a[356] & b[189])^(a[355] & b[190])^(a[354] & b[191])^(a[353] & b[192])^(a[352] & b[193])^(a[351] & b[194])^(a[350] & b[195])^(a[349] & b[196])^(a[348] & b[197])^(a[347] & b[198])^(a[346] & b[199])^(a[345] & b[200])^(a[344] & b[201])^(a[343] & b[202])^(a[342] & b[203])^(a[341] & b[204])^(a[340] & b[205])^(a[339] & b[206])^(a[338] & b[207])^(a[337] & b[208])^(a[336] & b[209])^(a[335] & b[210])^(a[334] & b[211])^(a[333] & b[212])^(a[332] & b[213])^(a[331] & b[214])^(a[330] & b[215])^(a[329] & b[216])^(a[328] & b[217])^(a[327] & b[218])^(a[326] & b[219])^(a[325] & b[220])^(a[324] & b[221])^(a[323] & b[222])^(a[322] & b[223])^(a[321] & b[224])^(a[320] & b[225])^(a[319] & b[226])^(a[318] & b[227])^(a[317] & b[228])^(a[316] & b[229])^(a[315] & b[230])^(a[314] & b[231])^(a[313] & b[232])^(a[312] & b[233])^(a[311] & b[234])^(a[310] & b[235])^(a[309] & b[236])^(a[308] & b[237])^(a[307] & b[238])^(a[306] & b[239])^(a[305] & b[240])^(a[304] & b[241])^(a[303] & b[242])^(a[302] & b[243])^(a[301] & b[244])^(a[300] & b[245])^(a[299] & b[246])^(a[298] & b[247])^(a[297] & b[248])^(a[296] & b[249])^(a[295] & b[250])^(a[294] & b[251])^(a[293] & b[252])^(a[292] & b[253])^(a[291] & b[254])^(a[290] & b[255])^(a[289] & b[256])^(a[288] & b[257])^(a[287] & b[258])^(a[286] & b[259])^(a[285] & b[260])^(a[284] & b[261])^(a[283] & b[262])^(a[282] & b[263])^(a[281] & b[264])^(a[280] & b[265])^(a[279] & b[266])^(a[278] & b[267])^(a[277] & b[268])^(a[276] & b[269])^(a[275] & b[270])^(a[274] & b[271])^(a[273] & b[272])^(a[272] & b[273])^(a[271] & b[274])^(a[270] & b[275])^(a[269] & b[276])^(a[268] & b[277])^(a[267] & b[278])^(a[266] & b[279])^(a[265] & b[280])^(a[264] & b[281])^(a[263] & b[282])^(a[262] & b[283])^(a[261] & b[284])^(a[260] & b[285])^(a[259] & b[286])^(a[258] & b[287])^(a[257] & b[288])^(a[256] & b[289])^(a[255] & b[290])^(a[254] & b[291])^(a[253] & b[292])^(a[252] & b[293])^(a[251] & b[294])^(a[250] & b[295])^(a[249] & b[296])^(a[248] & b[297])^(a[247] & b[298])^(a[246] & b[299])^(a[245] & b[300])^(a[244] & b[301])^(a[243] & b[302])^(a[242] & b[303])^(a[241] & b[304])^(a[240] & b[305])^(a[239] & b[306])^(a[238] & b[307])^(a[237] & b[308])^(a[236] & b[309])^(a[235] & b[310])^(a[234] & b[311])^(a[233] & b[312])^(a[232] & b[313])^(a[231] & b[314])^(a[230] & b[315])^(a[229] & b[316])^(a[228] & b[317])^(a[227] & b[318])^(a[226] & b[319])^(a[225] & b[320])^(a[224] & b[321])^(a[223] & b[322])^(a[222] & b[323])^(a[221] & b[324])^(a[220] & b[325])^(a[219] & b[326])^(a[218] & b[327])^(a[217] & b[328])^(a[216] & b[329])^(a[215] & b[330])^(a[214] & b[331])^(a[213] & b[332])^(a[212] & b[333])^(a[211] & b[334])^(a[210] & b[335])^(a[209] & b[336])^(a[208] & b[337])^(a[207] & b[338])^(a[206] & b[339])^(a[205] & b[340])^(a[204] & b[341])^(a[203] & b[342])^(a[202] & b[343])^(a[201] & b[344])^(a[200] & b[345])^(a[199] & b[346])^(a[198] & b[347])^(a[197] & b[348])^(a[196] & b[349])^(a[195] & b[350])^(a[194] & b[351])^(a[193] & b[352])^(a[192] & b[353])^(a[191] & b[354])^(a[190] & b[355])^(a[189] & b[356])^(a[188] & b[357])^(a[187] & b[358])^(a[186] & b[359])^(a[185] & b[360])^(a[184] & b[361])^(a[183] & b[362])^(a[182] & b[363])^(a[181] & b[364])^(a[180] & b[365])^(a[179] & b[366])^(a[178] & b[367])^(a[177] & b[368])^(a[176] & b[369])^(a[175] & b[370])^(a[174] & b[371])^(a[173] & b[372])^(a[172] & b[373])^(a[171] & b[374])^(a[170] & b[375])^(a[169] & b[376])^(a[168] & b[377])^(a[167] & b[378])^(a[166] & b[379])^(a[165] & b[380])^(a[164] & b[381])^(a[163] & b[382])^(a[162] & b[383])^(a[161] & b[384])^(a[160] & b[385])^(a[159] & b[386])^(a[158] & b[387])^(a[157] & b[388])^(a[156] & b[389])^(a[155] & b[390])^(a[154] & b[391])^(a[153] & b[392])^(a[152] & b[393])^(a[151] & b[394])^(a[150] & b[395])^(a[149] & b[396])^(a[148] & b[397])^(a[147] & b[398])^(a[146] & b[399])^(a[145] & b[400])^(a[144] & b[401])^(a[143] & b[402])^(a[142] & b[403])^(a[141] & b[404])^(a[140] & b[405])^(a[139] & b[406])^(a[138] & b[407])^(a[137] & b[408]);
assign y[546] = (a[408] & b[138])^(a[407] & b[139])^(a[406] & b[140])^(a[405] & b[141])^(a[404] & b[142])^(a[403] & b[143])^(a[402] & b[144])^(a[401] & b[145])^(a[400] & b[146])^(a[399] & b[147])^(a[398] & b[148])^(a[397] & b[149])^(a[396] & b[150])^(a[395] & b[151])^(a[394] & b[152])^(a[393] & b[153])^(a[392] & b[154])^(a[391] & b[155])^(a[390] & b[156])^(a[389] & b[157])^(a[388] & b[158])^(a[387] & b[159])^(a[386] & b[160])^(a[385] & b[161])^(a[384] & b[162])^(a[383] & b[163])^(a[382] & b[164])^(a[381] & b[165])^(a[380] & b[166])^(a[379] & b[167])^(a[378] & b[168])^(a[377] & b[169])^(a[376] & b[170])^(a[375] & b[171])^(a[374] & b[172])^(a[373] & b[173])^(a[372] & b[174])^(a[371] & b[175])^(a[370] & b[176])^(a[369] & b[177])^(a[368] & b[178])^(a[367] & b[179])^(a[366] & b[180])^(a[365] & b[181])^(a[364] & b[182])^(a[363] & b[183])^(a[362] & b[184])^(a[361] & b[185])^(a[360] & b[186])^(a[359] & b[187])^(a[358] & b[188])^(a[357] & b[189])^(a[356] & b[190])^(a[355] & b[191])^(a[354] & b[192])^(a[353] & b[193])^(a[352] & b[194])^(a[351] & b[195])^(a[350] & b[196])^(a[349] & b[197])^(a[348] & b[198])^(a[347] & b[199])^(a[346] & b[200])^(a[345] & b[201])^(a[344] & b[202])^(a[343] & b[203])^(a[342] & b[204])^(a[341] & b[205])^(a[340] & b[206])^(a[339] & b[207])^(a[338] & b[208])^(a[337] & b[209])^(a[336] & b[210])^(a[335] & b[211])^(a[334] & b[212])^(a[333] & b[213])^(a[332] & b[214])^(a[331] & b[215])^(a[330] & b[216])^(a[329] & b[217])^(a[328] & b[218])^(a[327] & b[219])^(a[326] & b[220])^(a[325] & b[221])^(a[324] & b[222])^(a[323] & b[223])^(a[322] & b[224])^(a[321] & b[225])^(a[320] & b[226])^(a[319] & b[227])^(a[318] & b[228])^(a[317] & b[229])^(a[316] & b[230])^(a[315] & b[231])^(a[314] & b[232])^(a[313] & b[233])^(a[312] & b[234])^(a[311] & b[235])^(a[310] & b[236])^(a[309] & b[237])^(a[308] & b[238])^(a[307] & b[239])^(a[306] & b[240])^(a[305] & b[241])^(a[304] & b[242])^(a[303] & b[243])^(a[302] & b[244])^(a[301] & b[245])^(a[300] & b[246])^(a[299] & b[247])^(a[298] & b[248])^(a[297] & b[249])^(a[296] & b[250])^(a[295] & b[251])^(a[294] & b[252])^(a[293] & b[253])^(a[292] & b[254])^(a[291] & b[255])^(a[290] & b[256])^(a[289] & b[257])^(a[288] & b[258])^(a[287] & b[259])^(a[286] & b[260])^(a[285] & b[261])^(a[284] & b[262])^(a[283] & b[263])^(a[282] & b[264])^(a[281] & b[265])^(a[280] & b[266])^(a[279] & b[267])^(a[278] & b[268])^(a[277] & b[269])^(a[276] & b[270])^(a[275] & b[271])^(a[274] & b[272])^(a[273] & b[273])^(a[272] & b[274])^(a[271] & b[275])^(a[270] & b[276])^(a[269] & b[277])^(a[268] & b[278])^(a[267] & b[279])^(a[266] & b[280])^(a[265] & b[281])^(a[264] & b[282])^(a[263] & b[283])^(a[262] & b[284])^(a[261] & b[285])^(a[260] & b[286])^(a[259] & b[287])^(a[258] & b[288])^(a[257] & b[289])^(a[256] & b[290])^(a[255] & b[291])^(a[254] & b[292])^(a[253] & b[293])^(a[252] & b[294])^(a[251] & b[295])^(a[250] & b[296])^(a[249] & b[297])^(a[248] & b[298])^(a[247] & b[299])^(a[246] & b[300])^(a[245] & b[301])^(a[244] & b[302])^(a[243] & b[303])^(a[242] & b[304])^(a[241] & b[305])^(a[240] & b[306])^(a[239] & b[307])^(a[238] & b[308])^(a[237] & b[309])^(a[236] & b[310])^(a[235] & b[311])^(a[234] & b[312])^(a[233] & b[313])^(a[232] & b[314])^(a[231] & b[315])^(a[230] & b[316])^(a[229] & b[317])^(a[228] & b[318])^(a[227] & b[319])^(a[226] & b[320])^(a[225] & b[321])^(a[224] & b[322])^(a[223] & b[323])^(a[222] & b[324])^(a[221] & b[325])^(a[220] & b[326])^(a[219] & b[327])^(a[218] & b[328])^(a[217] & b[329])^(a[216] & b[330])^(a[215] & b[331])^(a[214] & b[332])^(a[213] & b[333])^(a[212] & b[334])^(a[211] & b[335])^(a[210] & b[336])^(a[209] & b[337])^(a[208] & b[338])^(a[207] & b[339])^(a[206] & b[340])^(a[205] & b[341])^(a[204] & b[342])^(a[203] & b[343])^(a[202] & b[344])^(a[201] & b[345])^(a[200] & b[346])^(a[199] & b[347])^(a[198] & b[348])^(a[197] & b[349])^(a[196] & b[350])^(a[195] & b[351])^(a[194] & b[352])^(a[193] & b[353])^(a[192] & b[354])^(a[191] & b[355])^(a[190] & b[356])^(a[189] & b[357])^(a[188] & b[358])^(a[187] & b[359])^(a[186] & b[360])^(a[185] & b[361])^(a[184] & b[362])^(a[183] & b[363])^(a[182] & b[364])^(a[181] & b[365])^(a[180] & b[366])^(a[179] & b[367])^(a[178] & b[368])^(a[177] & b[369])^(a[176] & b[370])^(a[175] & b[371])^(a[174] & b[372])^(a[173] & b[373])^(a[172] & b[374])^(a[171] & b[375])^(a[170] & b[376])^(a[169] & b[377])^(a[168] & b[378])^(a[167] & b[379])^(a[166] & b[380])^(a[165] & b[381])^(a[164] & b[382])^(a[163] & b[383])^(a[162] & b[384])^(a[161] & b[385])^(a[160] & b[386])^(a[159] & b[387])^(a[158] & b[388])^(a[157] & b[389])^(a[156] & b[390])^(a[155] & b[391])^(a[154] & b[392])^(a[153] & b[393])^(a[152] & b[394])^(a[151] & b[395])^(a[150] & b[396])^(a[149] & b[397])^(a[148] & b[398])^(a[147] & b[399])^(a[146] & b[400])^(a[145] & b[401])^(a[144] & b[402])^(a[143] & b[403])^(a[142] & b[404])^(a[141] & b[405])^(a[140] & b[406])^(a[139] & b[407])^(a[138] & b[408]);
assign y[547] = (a[408] & b[139])^(a[407] & b[140])^(a[406] & b[141])^(a[405] & b[142])^(a[404] & b[143])^(a[403] & b[144])^(a[402] & b[145])^(a[401] & b[146])^(a[400] & b[147])^(a[399] & b[148])^(a[398] & b[149])^(a[397] & b[150])^(a[396] & b[151])^(a[395] & b[152])^(a[394] & b[153])^(a[393] & b[154])^(a[392] & b[155])^(a[391] & b[156])^(a[390] & b[157])^(a[389] & b[158])^(a[388] & b[159])^(a[387] & b[160])^(a[386] & b[161])^(a[385] & b[162])^(a[384] & b[163])^(a[383] & b[164])^(a[382] & b[165])^(a[381] & b[166])^(a[380] & b[167])^(a[379] & b[168])^(a[378] & b[169])^(a[377] & b[170])^(a[376] & b[171])^(a[375] & b[172])^(a[374] & b[173])^(a[373] & b[174])^(a[372] & b[175])^(a[371] & b[176])^(a[370] & b[177])^(a[369] & b[178])^(a[368] & b[179])^(a[367] & b[180])^(a[366] & b[181])^(a[365] & b[182])^(a[364] & b[183])^(a[363] & b[184])^(a[362] & b[185])^(a[361] & b[186])^(a[360] & b[187])^(a[359] & b[188])^(a[358] & b[189])^(a[357] & b[190])^(a[356] & b[191])^(a[355] & b[192])^(a[354] & b[193])^(a[353] & b[194])^(a[352] & b[195])^(a[351] & b[196])^(a[350] & b[197])^(a[349] & b[198])^(a[348] & b[199])^(a[347] & b[200])^(a[346] & b[201])^(a[345] & b[202])^(a[344] & b[203])^(a[343] & b[204])^(a[342] & b[205])^(a[341] & b[206])^(a[340] & b[207])^(a[339] & b[208])^(a[338] & b[209])^(a[337] & b[210])^(a[336] & b[211])^(a[335] & b[212])^(a[334] & b[213])^(a[333] & b[214])^(a[332] & b[215])^(a[331] & b[216])^(a[330] & b[217])^(a[329] & b[218])^(a[328] & b[219])^(a[327] & b[220])^(a[326] & b[221])^(a[325] & b[222])^(a[324] & b[223])^(a[323] & b[224])^(a[322] & b[225])^(a[321] & b[226])^(a[320] & b[227])^(a[319] & b[228])^(a[318] & b[229])^(a[317] & b[230])^(a[316] & b[231])^(a[315] & b[232])^(a[314] & b[233])^(a[313] & b[234])^(a[312] & b[235])^(a[311] & b[236])^(a[310] & b[237])^(a[309] & b[238])^(a[308] & b[239])^(a[307] & b[240])^(a[306] & b[241])^(a[305] & b[242])^(a[304] & b[243])^(a[303] & b[244])^(a[302] & b[245])^(a[301] & b[246])^(a[300] & b[247])^(a[299] & b[248])^(a[298] & b[249])^(a[297] & b[250])^(a[296] & b[251])^(a[295] & b[252])^(a[294] & b[253])^(a[293] & b[254])^(a[292] & b[255])^(a[291] & b[256])^(a[290] & b[257])^(a[289] & b[258])^(a[288] & b[259])^(a[287] & b[260])^(a[286] & b[261])^(a[285] & b[262])^(a[284] & b[263])^(a[283] & b[264])^(a[282] & b[265])^(a[281] & b[266])^(a[280] & b[267])^(a[279] & b[268])^(a[278] & b[269])^(a[277] & b[270])^(a[276] & b[271])^(a[275] & b[272])^(a[274] & b[273])^(a[273] & b[274])^(a[272] & b[275])^(a[271] & b[276])^(a[270] & b[277])^(a[269] & b[278])^(a[268] & b[279])^(a[267] & b[280])^(a[266] & b[281])^(a[265] & b[282])^(a[264] & b[283])^(a[263] & b[284])^(a[262] & b[285])^(a[261] & b[286])^(a[260] & b[287])^(a[259] & b[288])^(a[258] & b[289])^(a[257] & b[290])^(a[256] & b[291])^(a[255] & b[292])^(a[254] & b[293])^(a[253] & b[294])^(a[252] & b[295])^(a[251] & b[296])^(a[250] & b[297])^(a[249] & b[298])^(a[248] & b[299])^(a[247] & b[300])^(a[246] & b[301])^(a[245] & b[302])^(a[244] & b[303])^(a[243] & b[304])^(a[242] & b[305])^(a[241] & b[306])^(a[240] & b[307])^(a[239] & b[308])^(a[238] & b[309])^(a[237] & b[310])^(a[236] & b[311])^(a[235] & b[312])^(a[234] & b[313])^(a[233] & b[314])^(a[232] & b[315])^(a[231] & b[316])^(a[230] & b[317])^(a[229] & b[318])^(a[228] & b[319])^(a[227] & b[320])^(a[226] & b[321])^(a[225] & b[322])^(a[224] & b[323])^(a[223] & b[324])^(a[222] & b[325])^(a[221] & b[326])^(a[220] & b[327])^(a[219] & b[328])^(a[218] & b[329])^(a[217] & b[330])^(a[216] & b[331])^(a[215] & b[332])^(a[214] & b[333])^(a[213] & b[334])^(a[212] & b[335])^(a[211] & b[336])^(a[210] & b[337])^(a[209] & b[338])^(a[208] & b[339])^(a[207] & b[340])^(a[206] & b[341])^(a[205] & b[342])^(a[204] & b[343])^(a[203] & b[344])^(a[202] & b[345])^(a[201] & b[346])^(a[200] & b[347])^(a[199] & b[348])^(a[198] & b[349])^(a[197] & b[350])^(a[196] & b[351])^(a[195] & b[352])^(a[194] & b[353])^(a[193] & b[354])^(a[192] & b[355])^(a[191] & b[356])^(a[190] & b[357])^(a[189] & b[358])^(a[188] & b[359])^(a[187] & b[360])^(a[186] & b[361])^(a[185] & b[362])^(a[184] & b[363])^(a[183] & b[364])^(a[182] & b[365])^(a[181] & b[366])^(a[180] & b[367])^(a[179] & b[368])^(a[178] & b[369])^(a[177] & b[370])^(a[176] & b[371])^(a[175] & b[372])^(a[174] & b[373])^(a[173] & b[374])^(a[172] & b[375])^(a[171] & b[376])^(a[170] & b[377])^(a[169] & b[378])^(a[168] & b[379])^(a[167] & b[380])^(a[166] & b[381])^(a[165] & b[382])^(a[164] & b[383])^(a[163] & b[384])^(a[162] & b[385])^(a[161] & b[386])^(a[160] & b[387])^(a[159] & b[388])^(a[158] & b[389])^(a[157] & b[390])^(a[156] & b[391])^(a[155] & b[392])^(a[154] & b[393])^(a[153] & b[394])^(a[152] & b[395])^(a[151] & b[396])^(a[150] & b[397])^(a[149] & b[398])^(a[148] & b[399])^(a[147] & b[400])^(a[146] & b[401])^(a[145] & b[402])^(a[144] & b[403])^(a[143] & b[404])^(a[142] & b[405])^(a[141] & b[406])^(a[140] & b[407])^(a[139] & b[408]);
assign y[548] = (a[408] & b[140])^(a[407] & b[141])^(a[406] & b[142])^(a[405] & b[143])^(a[404] & b[144])^(a[403] & b[145])^(a[402] & b[146])^(a[401] & b[147])^(a[400] & b[148])^(a[399] & b[149])^(a[398] & b[150])^(a[397] & b[151])^(a[396] & b[152])^(a[395] & b[153])^(a[394] & b[154])^(a[393] & b[155])^(a[392] & b[156])^(a[391] & b[157])^(a[390] & b[158])^(a[389] & b[159])^(a[388] & b[160])^(a[387] & b[161])^(a[386] & b[162])^(a[385] & b[163])^(a[384] & b[164])^(a[383] & b[165])^(a[382] & b[166])^(a[381] & b[167])^(a[380] & b[168])^(a[379] & b[169])^(a[378] & b[170])^(a[377] & b[171])^(a[376] & b[172])^(a[375] & b[173])^(a[374] & b[174])^(a[373] & b[175])^(a[372] & b[176])^(a[371] & b[177])^(a[370] & b[178])^(a[369] & b[179])^(a[368] & b[180])^(a[367] & b[181])^(a[366] & b[182])^(a[365] & b[183])^(a[364] & b[184])^(a[363] & b[185])^(a[362] & b[186])^(a[361] & b[187])^(a[360] & b[188])^(a[359] & b[189])^(a[358] & b[190])^(a[357] & b[191])^(a[356] & b[192])^(a[355] & b[193])^(a[354] & b[194])^(a[353] & b[195])^(a[352] & b[196])^(a[351] & b[197])^(a[350] & b[198])^(a[349] & b[199])^(a[348] & b[200])^(a[347] & b[201])^(a[346] & b[202])^(a[345] & b[203])^(a[344] & b[204])^(a[343] & b[205])^(a[342] & b[206])^(a[341] & b[207])^(a[340] & b[208])^(a[339] & b[209])^(a[338] & b[210])^(a[337] & b[211])^(a[336] & b[212])^(a[335] & b[213])^(a[334] & b[214])^(a[333] & b[215])^(a[332] & b[216])^(a[331] & b[217])^(a[330] & b[218])^(a[329] & b[219])^(a[328] & b[220])^(a[327] & b[221])^(a[326] & b[222])^(a[325] & b[223])^(a[324] & b[224])^(a[323] & b[225])^(a[322] & b[226])^(a[321] & b[227])^(a[320] & b[228])^(a[319] & b[229])^(a[318] & b[230])^(a[317] & b[231])^(a[316] & b[232])^(a[315] & b[233])^(a[314] & b[234])^(a[313] & b[235])^(a[312] & b[236])^(a[311] & b[237])^(a[310] & b[238])^(a[309] & b[239])^(a[308] & b[240])^(a[307] & b[241])^(a[306] & b[242])^(a[305] & b[243])^(a[304] & b[244])^(a[303] & b[245])^(a[302] & b[246])^(a[301] & b[247])^(a[300] & b[248])^(a[299] & b[249])^(a[298] & b[250])^(a[297] & b[251])^(a[296] & b[252])^(a[295] & b[253])^(a[294] & b[254])^(a[293] & b[255])^(a[292] & b[256])^(a[291] & b[257])^(a[290] & b[258])^(a[289] & b[259])^(a[288] & b[260])^(a[287] & b[261])^(a[286] & b[262])^(a[285] & b[263])^(a[284] & b[264])^(a[283] & b[265])^(a[282] & b[266])^(a[281] & b[267])^(a[280] & b[268])^(a[279] & b[269])^(a[278] & b[270])^(a[277] & b[271])^(a[276] & b[272])^(a[275] & b[273])^(a[274] & b[274])^(a[273] & b[275])^(a[272] & b[276])^(a[271] & b[277])^(a[270] & b[278])^(a[269] & b[279])^(a[268] & b[280])^(a[267] & b[281])^(a[266] & b[282])^(a[265] & b[283])^(a[264] & b[284])^(a[263] & b[285])^(a[262] & b[286])^(a[261] & b[287])^(a[260] & b[288])^(a[259] & b[289])^(a[258] & b[290])^(a[257] & b[291])^(a[256] & b[292])^(a[255] & b[293])^(a[254] & b[294])^(a[253] & b[295])^(a[252] & b[296])^(a[251] & b[297])^(a[250] & b[298])^(a[249] & b[299])^(a[248] & b[300])^(a[247] & b[301])^(a[246] & b[302])^(a[245] & b[303])^(a[244] & b[304])^(a[243] & b[305])^(a[242] & b[306])^(a[241] & b[307])^(a[240] & b[308])^(a[239] & b[309])^(a[238] & b[310])^(a[237] & b[311])^(a[236] & b[312])^(a[235] & b[313])^(a[234] & b[314])^(a[233] & b[315])^(a[232] & b[316])^(a[231] & b[317])^(a[230] & b[318])^(a[229] & b[319])^(a[228] & b[320])^(a[227] & b[321])^(a[226] & b[322])^(a[225] & b[323])^(a[224] & b[324])^(a[223] & b[325])^(a[222] & b[326])^(a[221] & b[327])^(a[220] & b[328])^(a[219] & b[329])^(a[218] & b[330])^(a[217] & b[331])^(a[216] & b[332])^(a[215] & b[333])^(a[214] & b[334])^(a[213] & b[335])^(a[212] & b[336])^(a[211] & b[337])^(a[210] & b[338])^(a[209] & b[339])^(a[208] & b[340])^(a[207] & b[341])^(a[206] & b[342])^(a[205] & b[343])^(a[204] & b[344])^(a[203] & b[345])^(a[202] & b[346])^(a[201] & b[347])^(a[200] & b[348])^(a[199] & b[349])^(a[198] & b[350])^(a[197] & b[351])^(a[196] & b[352])^(a[195] & b[353])^(a[194] & b[354])^(a[193] & b[355])^(a[192] & b[356])^(a[191] & b[357])^(a[190] & b[358])^(a[189] & b[359])^(a[188] & b[360])^(a[187] & b[361])^(a[186] & b[362])^(a[185] & b[363])^(a[184] & b[364])^(a[183] & b[365])^(a[182] & b[366])^(a[181] & b[367])^(a[180] & b[368])^(a[179] & b[369])^(a[178] & b[370])^(a[177] & b[371])^(a[176] & b[372])^(a[175] & b[373])^(a[174] & b[374])^(a[173] & b[375])^(a[172] & b[376])^(a[171] & b[377])^(a[170] & b[378])^(a[169] & b[379])^(a[168] & b[380])^(a[167] & b[381])^(a[166] & b[382])^(a[165] & b[383])^(a[164] & b[384])^(a[163] & b[385])^(a[162] & b[386])^(a[161] & b[387])^(a[160] & b[388])^(a[159] & b[389])^(a[158] & b[390])^(a[157] & b[391])^(a[156] & b[392])^(a[155] & b[393])^(a[154] & b[394])^(a[153] & b[395])^(a[152] & b[396])^(a[151] & b[397])^(a[150] & b[398])^(a[149] & b[399])^(a[148] & b[400])^(a[147] & b[401])^(a[146] & b[402])^(a[145] & b[403])^(a[144] & b[404])^(a[143] & b[405])^(a[142] & b[406])^(a[141] & b[407])^(a[140] & b[408]);
assign y[549] = (a[408] & b[141])^(a[407] & b[142])^(a[406] & b[143])^(a[405] & b[144])^(a[404] & b[145])^(a[403] & b[146])^(a[402] & b[147])^(a[401] & b[148])^(a[400] & b[149])^(a[399] & b[150])^(a[398] & b[151])^(a[397] & b[152])^(a[396] & b[153])^(a[395] & b[154])^(a[394] & b[155])^(a[393] & b[156])^(a[392] & b[157])^(a[391] & b[158])^(a[390] & b[159])^(a[389] & b[160])^(a[388] & b[161])^(a[387] & b[162])^(a[386] & b[163])^(a[385] & b[164])^(a[384] & b[165])^(a[383] & b[166])^(a[382] & b[167])^(a[381] & b[168])^(a[380] & b[169])^(a[379] & b[170])^(a[378] & b[171])^(a[377] & b[172])^(a[376] & b[173])^(a[375] & b[174])^(a[374] & b[175])^(a[373] & b[176])^(a[372] & b[177])^(a[371] & b[178])^(a[370] & b[179])^(a[369] & b[180])^(a[368] & b[181])^(a[367] & b[182])^(a[366] & b[183])^(a[365] & b[184])^(a[364] & b[185])^(a[363] & b[186])^(a[362] & b[187])^(a[361] & b[188])^(a[360] & b[189])^(a[359] & b[190])^(a[358] & b[191])^(a[357] & b[192])^(a[356] & b[193])^(a[355] & b[194])^(a[354] & b[195])^(a[353] & b[196])^(a[352] & b[197])^(a[351] & b[198])^(a[350] & b[199])^(a[349] & b[200])^(a[348] & b[201])^(a[347] & b[202])^(a[346] & b[203])^(a[345] & b[204])^(a[344] & b[205])^(a[343] & b[206])^(a[342] & b[207])^(a[341] & b[208])^(a[340] & b[209])^(a[339] & b[210])^(a[338] & b[211])^(a[337] & b[212])^(a[336] & b[213])^(a[335] & b[214])^(a[334] & b[215])^(a[333] & b[216])^(a[332] & b[217])^(a[331] & b[218])^(a[330] & b[219])^(a[329] & b[220])^(a[328] & b[221])^(a[327] & b[222])^(a[326] & b[223])^(a[325] & b[224])^(a[324] & b[225])^(a[323] & b[226])^(a[322] & b[227])^(a[321] & b[228])^(a[320] & b[229])^(a[319] & b[230])^(a[318] & b[231])^(a[317] & b[232])^(a[316] & b[233])^(a[315] & b[234])^(a[314] & b[235])^(a[313] & b[236])^(a[312] & b[237])^(a[311] & b[238])^(a[310] & b[239])^(a[309] & b[240])^(a[308] & b[241])^(a[307] & b[242])^(a[306] & b[243])^(a[305] & b[244])^(a[304] & b[245])^(a[303] & b[246])^(a[302] & b[247])^(a[301] & b[248])^(a[300] & b[249])^(a[299] & b[250])^(a[298] & b[251])^(a[297] & b[252])^(a[296] & b[253])^(a[295] & b[254])^(a[294] & b[255])^(a[293] & b[256])^(a[292] & b[257])^(a[291] & b[258])^(a[290] & b[259])^(a[289] & b[260])^(a[288] & b[261])^(a[287] & b[262])^(a[286] & b[263])^(a[285] & b[264])^(a[284] & b[265])^(a[283] & b[266])^(a[282] & b[267])^(a[281] & b[268])^(a[280] & b[269])^(a[279] & b[270])^(a[278] & b[271])^(a[277] & b[272])^(a[276] & b[273])^(a[275] & b[274])^(a[274] & b[275])^(a[273] & b[276])^(a[272] & b[277])^(a[271] & b[278])^(a[270] & b[279])^(a[269] & b[280])^(a[268] & b[281])^(a[267] & b[282])^(a[266] & b[283])^(a[265] & b[284])^(a[264] & b[285])^(a[263] & b[286])^(a[262] & b[287])^(a[261] & b[288])^(a[260] & b[289])^(a[259] & b[290])^(a[258] & b[291])^(a[257] & b[292])^(a[256] & b[293])^(a[255] & b[294])^(a[254] & b[295])^(a[253] & b[296])^(a[252] & b[297])^(a[251] & b[298])^(a[250] & b[299])^(a[249] & b[300])^(a[248] & b[301])^(a[247] & b[302])^(a[246] & b[303])^(a[245] & b[304])^(a[244] & b[305])^(a[243] & b[306])^(a[242] & b[307])^(a[241] & b[308])^(a[240] & b[309])^(a[239] & b[310])^(a[238] & b[311])^(a[237] & b[312])^(a[236] & b[313])^(a[235] & b[314])^(a[234] & b[315])^(a[233] & b[316])^(a[232] & b[317])^(a[231] & b[318])^(a[230] & b[319])^(a[229] & b[320])^(a[228] & b[321])^(a[227] & b[322])^(a[226] & b[323])^(a[225] & b[324])^(a[224] & b[325])^(a[223] & b[326])^(a[222] & b[327])^(a[221] & b[328])^(a[220] & b[329])^(a[219] & b[330])^(a[218] & b[331])^(a[217] & b[332])^(a[216] & b[333])^(a[215] & b[334])^(a[214] & b[335])^(a[213] & b[336])^(a[212] & b[337])^(a[211] & b[338])^(a[210] & b[339])^(a[209] & b[340])^(a[208] & b[341])^(a[207] & b[342])^(a[206] & b[343])^(a[205] & b[344])^(a[204] & b[345])^(a[203] & b[346])^(a[202] & b[347])^(a[201] & b[348])^(a[200] & b[349])^(a[199] & b[350])^(a[198] & b[351])^(a[197] & b[352])^(a[196] & b[353])^(a[195] & b[354])^(a[194] & b[355])^(a[193] & b[356])^(a[192] & b[357])^(a[191] & b[358])^(a[190] & b[359])^(a[189] & b[360])^(a[188] & b[361])^(a[187] & b[362])^(a[186] & b[363])^(a[185] & b[364])^(a[184] & b[365])^(a[183] & b[366])^(a[182] & b[367])^(a[181] & b[368])^(a[180] & b[369])^(a[179] & b[370])^(a[178] & b[371])^(a[177] & b[372])^(a[176] & b[373])^(a[175] & b[374])^(a[174] & b[375])^(a[173] & b[376])^(a[172] & b[377])^(a[171] & b[378])^(a[170] & b[379])^(a[169] & b[380])^(a[168] & b[381])^(a[167] & b[382])^(a[166] & b[383])^(a[165] & b[384])^(a[164] & b[385])^(a[163] & b[386])^(a[162] & b[387])^(a[161] & b[388])^(a[160] & b[389])^(a[159] & b[390])^(a[158] & b[391])^(a[157] & b[392])^(a[156] & b[393])^(a[155] & b[394])^(a[154] & b[395])^(a[153] & b[396])^(a[152] & b[397])^(a[151] & b[398])^(a[150] & b[399])^(a[149] & b[400])^(a[148] & b[401])^(a[147] & b[402])^(a[146] & b[403])^(a[145] & b[404])^(a[144] & b[405])^(a[143] & b[406])^(a[142] & b[407])^(a[141] & b[408]);
assign y[550] = (a[408] & b[142])^(a[407] & b[143])^(a[406] & b[144])^(a[405] & b[145])^(a[404] & b[146])^(a[403] & b[147])^(a[402] & b[148])^(a[401] & b[149])^(a[400] & b[150])^(a[399] & b[151])^(a[398] & b[152])^(a[397] & b[153])^(a[396] & b[154])^(a[395] & b[155])^(a[394] & b[156])^(a[393] & b[157])^(a[392] & b[158])^(a[391] & b[159])^(a[390] & b[160])^(a[389] & b[161])^(a[388] & b[162])^(a[387] & b[163])^(a[386] & b[164])^(a[385] & b[165])^(a[384] & b[166])^(a[383] & b[167])^(a[382] & b[168])^(a[381] & b[169])^(a[380] & b[170])^(a[379] & b[171])^(a[378] & b[172])^(a[377] & b[173])^(a[376] & b[174])^(a[375] & b[175])^(a[374] & b[176])^(a[373] & b[177])^(a[372] & b[178])^(a[371] & b[179])^(a[370] & b[180])^(a[369] & b[181])^(a[368] & b[182])^(a[367] & b[183])^(a[366] & b[184])^(a[365] & b[185])^(a[364] & b[186])^(a[363] & b[187])^(a[362] & b[188])^(a[361] & b[189])^(a[360] & b[190])^(a[359] & b[191])^(a[358] & b[192])^(a[357] & b[193])^(a[356] & b[194])^(a[355] & b[195])^(a[354] & b[196])^(a[353] & b[197])^(a[352] & b[198])^(a[351] & b[199])^(a[350] & b[200])^(a[349] & b[201])^(a[348] & b[202])^(a[347] & b[203])^(a[346] & b[204])^(a[345] & b[205])^(a[344] & b[206])^(a[343] & b[207])^(a[342] & b[208])^(a[341] & b[209])^(a[340] & b[210])^(a[339] & b[211])^(a[338] & b[212])^(a[337] & b[213])^(a[336] & b[214])^(a[335] & b[215])^(a[334] & b[216])^(a[333] & b[217])^(a[332] & b[218])^(a[331] & b[219])^(a[330] & b[220])^(a[329] & b[221])^(a[328] & b[222])^(a[327] & b[223])^(a[326] & b[224])^(a[325] & b[225])^(a[324] & b[226])^(a[323] & b[227])^(a[322] & b[228])^(a[321] & b[229])^(a[320] & b[230])^(a[319] & b[231])^(a[318] & b[232])^(a[317] & b[233])^(a[316] & b[234])^(a[315] & b[235])^(a[314] & b[236])^(a[313] & b[237])^(a[312] & b[238])^(a[311] & b[239])^(a[310] & b[240])^(a[309] & b[241])^(a[308] & b[242])^(a[307] & b[243])^(a[306] & b[244])^(a[305] & b[245])^(a[304] & b[246])^(a[303] & b[247])^(a[302] & b[248])^(a[301] & b[249])^(a[300] & b[250])^(a[299] & b[251])^(a[298] & b[252])^(a[297] & b[253])^(a[296] & b[254])^(a[295] & b[255])^(a[294] & b[256])^(a[293] & b[257])^(a[292] & b[258])^(a[291] & b[259])^(a[290] & b[260])^(a[289] & b[261])^(a[288] & b[262])^(a[287] & b[263])^(a[286] & b[264])^(a[285] & b[265])^(a[284] & b[266])^(a[283] & b[267])^(a[282] & b[268])^(a[281] & b[269])^(a[280] & b[270])^(a[279] & b[271])^(a[278] & b[272])^(a[277] & b[273])^(a[276] & b[274])^(a[275] & b[275])^(a[274] & b[276])^(a[273] & b[277])^(a[272] & b[278])^(a[271] & b[279])^(a[270] & b[280])^(a[269] & b[281])^(a[268] & b[282])^(a[267] & b[283])^(a[266] & b[284])^(a[265] & b[285])^(a[264] & b[286])^(a[263] & b[287])^(a[262] & b[288])^(a[261] & b[289])^(a[260] & b[290])^(a[259] & b[291])^(a[258] & b[292])^(a[257] & b[293])^(a[256] & b[294])^(a[255] & b[295])^(a[254] & b[296])^(a[253] & b[297])^(a[252] & b[298])^(a[251] & b[299])^(a[250] & b[300])^(a[249] & b[301])^(a[248] & b[302])^(a[247] & b[303])^(a[246] & b[304])^(a[245] & b[305])^(a[244] & b[306])^(a[243] & b[307])^(a[242] & b[308])^(a[241] & b[309])^(a[240] & b[310])^(a[239] & b[311])^(a[238] & b[312])^(a[237] & b[313])^(a[236] & b[314])^(a[235] & b[315])^(a[234] & b[316])^(a[233] & b[317])^(a[232] & b[318])^(a[231] & b[319])^(a[230] & b[320])^(a[229] & b[321])^(a[228] & b[322])^(a[227] & b[323])^(a[226] & b[324])^(a[225] & b[325])^(a[224] & b[326])^(a[223] & b[327])^(a[222] & b[328])^(a[221] & b[329])^(a[220] & b[330])^(a[219] & b[331])^(a[218] & b[332])^(a[217] & b[333])^(a[216] & b[334])^(a[215] & b[335])^(a[214] & b[336])^(a[213] & b[337])^(a[212] & b[338])^(a[211] & b[339])^(a[210] & b[340])^(a[209] & b[341])^(a[208] & b[342])^(a[207] & b[343])^(a[206] & b[344])^(a[205] & b[345])^(a[204] & b[346])^(a[203] & b[347])^(a[202] & b[348])^(a[201] & b[349])^(a[200] & b[350])^(a[199] & b[351])^(a[198] & b[352])^(a[197] & b[353])^(a[196] & b[354])^(a[195] & b[355])^(a[194] & b[356])^(a[193] & b[357])^(a[192] & b[358])^(a[191] & b[359])^(a[190] & b[360])^(a[189] & b[361])^(a[188] & b[362])^(a[187] & b[363])^(a[186] & b[364])^(a[185] & b[365])^(a[184] & b[366])^(a[183] & b[367])^(a[182] & b[368])^(a[181] & b[369])^(a[180] & b[370])^(a[179] & b[371])^(a[178] & b[372])^(a[177] & b[373])^(a[176] & b[374])^(a[175] & b[375])^(a[174] & b[376])^(a[173] & b[377])^(a[172] & b[378])^(a[171] & b[379])^(a[170] & b[380])^(a[169] & b[381])^(a[168] & b[382])^(a[167] & b[383])^(a[166] & b[384])^(a[165] & b[385])^(a[164] & b[386])^(a[163] & b[387])^(a[162] & b[388])^(a[161] & b[389])^(a[160] & b[390])^(a[159] & b[391])^(a[158] & b[392])^(a[157] & b[393])^(a[156] & b[394])^(a[155] & b[395])^(a[154] & b[396])^(a[153] & b[397])^(a[152] & b[398])^(a[151] & b[399])^(a[150] & b[400])^(a[149] & b[401])^(a[148] & b[402])^(a[147] & b[403])^(a[146] & b[404])^(a[145] & b[405])^(a[144] & b[406])^(a[143] & b[407])^(a[142] & b[408]);
assign y[551] = (a[408] & b[143])^(a[407] & b[144])^(a[406] & b[145])^(a[405] & b[146])^(a[404] & b[147])^(a[403] & b[148])^(a[402] & b[149])^(a[401] & b[150])^(a[400] & b[151])^(a[399] & b[152])^(a[398] & b[153])^(a[397] & b[154])^(a[396] & b[155])^(a[395] & b[156])^(a[394] & b[157])^(a[393] & b[158])^(a[392] & b[159])^(a[391] & b[160])^(a[390] & b[161])^(a[389] & b[162])^(a[388] & b[163])^(a[387] & b[164])^(a[386] & b[165])^(a[385] & b[166])^(a[384] & b[167])^(a[383] & b[168])^(a[382] & b[169])^(a[381] & b[170])^(a[380] & b[171])^(a[379] & b[172])^(a[378] & b[173])^(a[377] & b[174])^(a[376] & b[175])^(a[375] & b[176])^(a[374] & b[177])^(a[373] & b[178])^(a[372] & b[179])^(a[371] & b[180])^(a[370] & b[181])^(a[369] & b[182])^(a[368] & b[183])^(a[367] & b[184])^(a[366] & b[185])^(a[365] & b[186])^(a[364] & b[187])^(a[363] & b[188])^(a[362] & b[189])^(a[361] & b[190])^(a[360] & b[191])^(a[359] & b[192])^(a[358] & b[193])^(a[357] & b[194])^(a[356] & b[195])^(a[355] & b[196])^(a[354] & b[197])^(a[353] & b[198])^(a[352] & b[199])^(a[351] & b[200])^(a[350] & b[201])^(a[349] & b[202])^(a[348] & b[203])^(a[347] & b[204])^(a[346] & b[205])^(a[345] & b[206])^(a[344] & b[207])^(a[343] & b[208])^(a[342] & b[209])^(a[341] & b[210])^(a[340] & b[211])^(a[339] & b[212])^(a[338] & b[213])^(a[337] & b[214])^(a[336] & b[215])^(a[335] & b[216])^(a[334] & b[217])^(a[333] & b[218])^(a[332] & b[219])^(a[331] & b[220])^(a[330] & b[221])^(a[329] & b[222])^(a[328] & b[223])^(a[327] & b[224])^(a[326] & b[225])^(a[325] & b[226])^(a[324] & b[227])^(a[323] & b[228])^(a[322] & b[229])^(a[321] & b[230])^(a[320] & b[231])^(a[319] & b[232])^(a[318] & b[233])^(a[317] & b[234])^(a[316] & b[235])^(a[315] & b[236])^(a[314] & b[237])^(a[313] & b[238])^(a[312] & b[239])^(a[311] & b[240])^(a[310] & b[241])^(a[309] & b[242])^(a[308] & b[243])^(a[307] & b[244])^(a[306] & b[245])^(a[305] & b[246])^(a[304] & b[247])^(a[303] & b[248])^(a[302] & b[249])^(a[301] & b[250])^(a[300] & b[251])^(a[299] & b[252])^(a[298] & b[253])^(a[297] & b[254])^(a[296] & b[255])^(a[295] & b[256])^(a[294] & b[257])^(a[293] & b[258])^(a[292] & b[259])^(a[291] & b[260])^(a[290] & b[261])^(a[289] & b[262])^(a[288] & b[263])^(a[287] & b[264])^(a[286] & b[265])^(a[285] & b[266])^(a[284] & b[267])^(a[283] & b[268])^(a[282] & b[269])^(a[281] & b[270])^(a[280] & b[271])^(a[279] & b[272])^(a[278] & b[273])^(a[277] & b[274])^(a[276] & b[275])^(a[275] & b[276])^(a[274] & b[277])^(a[273] & b[278])^(a[272] & b[279])^(a[271] & b[280])^(a[270] & b[281])^(a[269] & b[282])^(a[268] & b[283])^(a[267] & b[284])^(a[266] & b[285])^(a[265] & b[286])^(a[264] & b[287])^(a[263] & b[288])^(a[262] & b[289])^(a[261] & b[290])^(a[260] & b[291])^(a[259] & b[292])^(a[258] & b[293])^(a[257] & b[294])^(a[256] & b[295])^(a[255] & b[296])^(a[254] & b[297])^(a[253] & b[298])^(a[252] & b[299])^(a[251] & b[300])^(a[250] & b[301])^(a[249] & b[302])^(a[248] & b[303])^(a[247] & b[304])^(a[246] & b[305])^(a[245] & b[306])^(a[244] & b[307])^(a[243] & b[308])^(a[242] & b[309])^(a[241] & b[310])^(a[240] & b[311])^(a[239] & b[312])^(a[238] & b[313])^(a[237] & b[314])^(a[236] & b[315])^(a[235] & b[316])^(a[234] & b[317])^(a[233] & b[318])^(a[232] & b[319])^(a[231] & b[320])^(a[230] & b[321])^(a[229] & b[322])^(a[228] & b[323])^(a[227] & b[324])^(a[226] & b[325])^(a[225] & b[326])^(a[224] & b[327])^(a[223] & b[328])^(a[222] & b[329])^(a[221] & b[330])^(a[220] & b[331])^(a[219] & b[332])^(a[218] & b[333])^(a[217] & b[334])^(a[216] & b[335])^(a[215] & b[336])^(a[214] & b[337])^(a[213] & b[338])^(a[212] & b[339])^(a[211] & b[340])^(a[210] & b[341])^(a[209] & b[342])^(a[208] & b[343])^(a[207] & b[344])^(a[206] & b[345])^(a[205] & b[346])^(a[204] & b[347])^(a[203] & b[348])^(a[202] & b[349])^(a[201] & b[350])^(a[200] & b[351])^(a[199] & b[352])^(a[198] & b[353])^(a[197] & b[354])^(a[196] & b[355])^(a[195] & b[356])^(a[194] & b[357])^(a[193] & b[358])^(a[192] & b[359])^(a[191] & b[360])^(a[190] & b[361])^(a[189] & b[362])^(a[188] & b[363])^(a[187] & b[364])^(a[186] & b[365])^(a[185] & b[366])^(a[184] & b[367])^(a[183] & b[368])^(a[182] & b[369])^(a[181] & b[370])^(a[180] & b[371])^(a[179] & b[372])^(a[178] & b[373])^(a[177] & b[374])^(a[176] & b[375])^(a[175] & b[376])^(a[174] & b[377])^(a[173] & b[378])^(a[172] & b[379])^(a[171] & b[380])^(a[170] & b[381])^(a[169] & b[382])^(a[168] & b[383])^(a[167] & b[384])^(a[166] & b[385])^(a[165] & b[386])^(a[164] & b[387])^(a[163] & b[388])^(a[162] & b[389])^(a[161] & b[390])^(a[160] & b[391])^(a[159] & b[392])^(a[158] & b[393])^(a[157] & b[394])^(a[156] & b[395])^(a[155] & b[396])^(a[154] & b[397])^(a[153] & b[398])^(a[152] & b[399])^(a[151] & b[400])^(a[150] & b[401])^(a[149] & b[402])^(a[148] & b[403])^(a[147] & b[404])^(a[146] & b[405])^(a[145] & b[406])^(a[144] & b[407])^(a[143] & b[408]);
assign y[552] = (a[408] & b[144])^(a[407] & b[145])^(a[406] & b[146])^(a[405] & b[147])^(a[404] & b[148])^(a[403] & b[149])^(a[402] & b[150])^(a[401] & b[151])^(a[400] & b[152])^(a[399] & b[153])^(a[398] & b[154])^(a[397] & b[155])^(a[396] & b[156])^(a[395] & b[157])^(a[394] & b[158])^(a[393] & b[159])^(a[392] & b[160])^(a[391] & b[161])^(a[390] & b[162])^(a[389] & b[163])^(a[388] & b[164])^(a[387] & b[165])^(a[386] & b[166])^(a[385] & b[167])^(a[384] & b[168])^(a[383] & b[169])^(a[382] & b[170])^(a[381] & b[171])^(a[380] & b[172])^(a[379] & b[173])^(a[378] & b[174])^(a[377] & b[175])^(a[376] & b[176])^(a[375] & b[177])^(a[374] & b[178])^(a[373] & b[179])^(a[372] & b[180])^(a[371] & b[181])^(a[370] & b[182])^(a[369] & b[183])^(a[368] & b[184])^(a[367] & b[185])^(a[366] & b[186])^(a[365] & b[187])^(a[364] & b[188])^(a[363] & b[189])^(a[362] & b[190])^(a[361] & b[191])^(a[360] & b[192])^(a[359] & b[193])^(a[358] & b[194])^(a[357] & b[195])^(a[356] & b[196])^(a[355] & b[197])^(a[354] & b[198])^(a[353] & b[199])^(a[352] & b[200])^(a[351] & b[201])^(a[350] & b[202])^(a[349] & b[203])^(a[348] & b[204])^(a[347] & b[205])^(a[346] & b[206])^(a[345] & b[207])^(a[344] & b[208])^(a[343] & b[209])^(a[342] & b[210])^(a[341] & b[211])^(a[340] & b[212])^(a[339] & b[213])^(a[338] & b[214])^(a[337] & b[215])^(a[336] & b[216])^(a[335] & b[217])^(a[334] & b[218])^(a[333] & b[219])^(a[332] & b[220])^(a[331] & b[221])^(a[330] & b[222])^(a[329] & b[223])^(a[328] & b[224])^(a[327] & b[225])^(a[326] & b[226])^(a[325] & b[227])^(a[324] & b[228])^(a[323] & b[229])^(a[322] & b[230])^(a[321] & b[231])^(a[320] & b[232])^(a[319] & b[233])^(a[318] & b[234])^(a[317] & b[235])^(a[316] & b[236])^(a[315] & b[237])^(a[314] & b[238])^(a[313] & b[239])^(a[312] & b[240])^(a[311] & b[241])^(a[310] & b[242])^(a[309] & b[243])^(a[308] & b[244])^(a[307] & b[245])^(a[306] & b[246])^(a[305] & b[247])^(a[304] & b[248])^(a[303] & b[249])^(a[302] & b[250])^(a[301] & b[251])^(a[300] & b[252])^(a[299] & b[253])^(a[298] & b[254])^(a[297] & b[255])^(a[296] & b[256])^(a[295] & b[257])^(a[294] & b[258])^(a[293] & b[259])^(a[292] & b[260])^(a[291] & b[261])^(a[290] & b[262])^(a[289] & b[263])^(a[288] & b[264])^(a[287] & b[265])^(a[286] & b[266])^(a[285] & b[267])^(a[284] & b[268])^(a[283] & b[269])^(a[282] & b[270])^(a[281] & b[271])^(a[280] & b[272])^(a[279] & b[273])^(a[278] & b[274])^(a[277] & b[275])^(a[276] & b[276])^(a[275] & b[277])^(a[274] & b[278])^(a[273] & b[279])^(a[272] & b[280])^(a[271] & b[281])^(a[270] & b[282])^(a[269] & b[283])^(a[268] & b[284])^(a[267] & b[285])^(a[266] & b[286])^(a[265] & b[287])^(a[264] & b[288])^(a[263] & b[289])^(a[262] & b[290])^(a[261] & b[291])^(a[260] & b[292])^(a[259] & b[293])^(a[258] & b[294])^(a[257] & b[295])^(a[256] & b[296])^(a[255] & b[297])^(a[254] & b[298])^(a[253] & b[299])^(a[252] & b[300])^(a[251] & b[301])^(a[250] & b[302])^(a[249] & b[303])^(a[248] & b[304])^(a[247] & b[305])^(a[246] & b[306])^(a[245] & b[307])^(a[244] & b[308])^(a[243] & b[309])^(a[242] & b[310])^(a[241] & b[311])^(a[240] & b[312])^(a[239] & b[313])^(a[238] & b[314])^(a[237] & b[315])^(a[236] & b[316])^(a[235] & b[317])^(a[234] & b[318])^(a[233] & b[319])^(a[232] & b[320])^(a[231] & b[321])^(a[230] & b[322])^(a[229] & b[323])^(a[228] & b[324])^(a[227] & b[325])^(a[226] & b[326])^(a[225] & b[327])^(a[224] & b[328])^(a[223] & b[329])^(a[222] & b[330])^(a[221] & b[331])^(a[220] & b[332])^(a[219] & b[333])^(a[218] & b[334])^(a[217] & b[335])^(a[216] & b[336])^(a[215] & b[337])^(a[214] & b[338])^(a[213] & b[339])^(a[212] & b[340])^(a[211] & b[341])^(a[210] & b[342])^(a[209] & b[343])^(a[208] & b[344])^(a[207] & b[345])^(a[206] & b[346])^(a[205] & b[347])^(a[204] & b[348])^(a[203] & b[349])^(a[202] & b[350])^(a[201] & b[351])^(a[200] & b[352])^(a[199] & b[353])^(a[198] & b[354])^(a[197] & b[355])^(a[196] & b[356])^(a[195] & b[357])^(a[194] & b[358])^(a[193] & b[359])^(a[192] & b[360])^(a[191] & b[361])^(a[190] & b[362])^(a[189] & b[363])^(a[188] & b[364])^(a[187] & b[365])^(a[186] & b[366])^(a[185] & b[367])^(a[184] & b[368])^(a[183] & b[369])^(a[182] & b[370])^(a[181] & b[371])^(a[180] & b[372])^(a[179] & b[373])^(a[178] & b[374])^(a[177] & b[375])^(a[176] & b[376])^(a[175] & b[377])^(a[174] & b[378])^(a[173] & b[379])^(a[172] & b[380])^(a[171] & b[381])^(a[170] & b[382])^(a[169] & b[383])^(a[168] & b[384])^(a[167] & b[385])^(a[166] & b[386])^(a[165] & b[387])^(a[164] & b[388])^(a[163] & b[389])^(a[162] & b[390])^(a[161] & b[391])^(a[160] & b[392])^(a[159] & b[393])^(a[158] & b[394])^(a[157] & b[395])^(a[156] & b[396])^(a[155] & b[397])^(a[154] & b[398])^(a[153] & b[399])^(a[152] & b[400])^(a[151] & b[401])^(a[150] & b[402])^(a[149] & b[403])^(a[148] & b[404])^(a[147] & b[405])^(a[146] & b[406])^(a[145] & b[407])^(a[144] & b[408]);
assign y[553] = (a[408] & b[145])^(a[407] & b[146])^(a[406] & b[147])^(a[405] & b[148])^(a[404] & b[149])^(a[403] & b[150])^(a[402] & b[151])^(a[401] & b[152])^(a[400] & b[153])^(a[399] & b[154])^(a[398] & b[155])^(a[397] & b[156])^(a[396] & b[157])^(a[395] & b[158])^(a[394] & b[159])^(a[393] & b[160])^(a[392] & b[161])^(a[391] & b[162])^(a[390] & b[163])^(a[389] & b[164])^(a[388] & b[165])^(a[387] & b[166])^(a[386] & b[167])^(a[385] & b[168])^(a[384] & b[169])^(a[383] & b[170])^(a[382] & b[171])^(a[381] & b[172])^(a[380] & b[173])^(a[379] & b[174])^(a[378] & b[175])^(a[377] & b[176])^(a[376] & b[177])^(a[375] & b[178])^(a[374] & b[179])^(a[373] & b[180])^(a[372] & b[181])^(a[371] & b[182])^(a[370] & b[183])^(a[369] & b[184])^(a[368] & b[185])^(a[367] & b[186])^(a[366] & b[187])^(a[365] & b[188])^(a[364] & b[189])^(a[363] & b[190])^(a[362] & b[191])^(a[361] & b[192])^(a[360] & b[193])^(a[359] & b[194])^(a[358] & b[195])^(a[357] & b[196])^(a[356] & b[197])^(a[355] & b[198])^(a[354] & b[199])^(a[353] & b[200])^(a[352] & b[201])^(a[351] & b[202])^(a[350] & b[203])^(a[349] & b[204])^(a[348] & b[205])^(a[347] & b[206])^(a[346] & b[207])^(a[345] & b[208])^(a[344] & b[209])^(a[343] & b[210])^(a[342] & b[211])^(a[341] & b[212])^(a[340] & b[213])^(a[339] & b[214])^(a[338] & b[215])^(a[337] & b[216])^(a[336] & b[217])^(a[335] & b[218])^(a[334] & b[219])^(a[333] & b[220])^(a[332] & b[221])^(a[331] & b[222])^(a[330] & b[223])^(a[329] & b[224])^(a[328] & b[225])^(a[327] & b[226])^(a[326] & b[227])^(a[325] & b[228])^(a[324] & b[229])^(a[323] & b[230])^(a[322] & b[231])^(a[321] & b[232])^(a[320] & b[233])^(a[319] & b[234])^(a[318] & b[235])^(a[317] & b[236])^(a[316] & b[237])^(a[315] & b[238])^(a[314] & b[239])^(a[313] & b[240])^(a[312] & b[241])^(a[311] & b[242])^(a[310] & b[243])^(a[309] & b[244])^(a[308] & b[245])^(a[307] & b[246])^(a[306] & b[247])^(a[305] & b[248])^(a[304] & b[249])^(a[303] & b[250])^(a[302] & b[251])^(a[301] & b[252])^(a[300] & b[253])^(a[299] & b[254])^(a[298] & b[255])^(a[297] & b[256])^(a[296] & b[257])^(a[295] & b[258])^(a[294] & b[259])^(a[293] & b[260])^(a[292] & b[261])^(a[291] & b[262])^(a[290] & b[263])^(a[289] & b[264])^(a[288] & b[265])^(a[287] & b[266])^(a[286] & b[267])^(a[285] & b[268])^(a[284] & b[269])^(a[283] & b[270])^(a[282] & b[271])^(a[281] & b[272])^(a[280] & b[273])^(a[279] & b[274])^(a[278] & b[275])^(a[277] & b[276])^(a[276] & b[277])^(a[275] & b[278])^(a[274] & b[279])^(a[273] & b[280])^(a[272] & b[281])^(a[271] & b[282])^(a[270] & b[283])^(a[269] & b[284])^(a[268] & b[285])^(a[267] & b[286])^(a[266] & b[287])^(a[265] & b[288])^(a[264] & b[289])^(a[263] & b[290])^(a[262] & b[291])^(a[261] & b[292])^(a[260] & b[293])^(a[259] & b[294])^(a[258] & b[295])^(a[257] & b[296])^(a[256] & b[297])^(a[255] & b[298])^(a[254] & b[299])^(a[253] & b[300])^(a[252] & b[301])^(a[251] & b[302])^(a[250] & b[303])^(a[249] & b[304])^(a[248] & b[305])^(a[247] & b[306])^(a[246] & b[307])^(a[245] & b[308])^(a[244] & b[309])^(a[243] & b[310])^(a[242] & b[311])^(a[241] & b[312])^(a[240] & b[313])^(a[239] & b[314])^(a[238] & b[315])^(a[237] & b[316])^(a[236] & b[317])^(a[235] & b[318])^(a[234] & b[319])^(a[233] & b[320])^(a[232] & b[321])^(a[231] & b[322])^(a[230] & b[323])^(a[229] & b[324])^(a[228] & b[325])^(a[227] & b[326])^(a[226] & b[327])^(a[225] & b[328])^(a[224] & b[329])^(a[223] & b[330])^(a[222] & b[331])^(a[221] & b[332])^(a[220] & b[333])^(a[219] & b[334])^(a[218] & b[335])^(a[217] & b[336])^(a[216] & b[337])^(a[215] & b[338])^(a[214] & b[339])^(a[213] & b[340])^(a[212] & b[341])^(a[211] & b[342])^(a[210] & b[343])^(a[209] & b[344])^(a[208] & b[345])^(a[207] & b[346])^(a[206] & b[347])^(a[205] & b[348])^(a[204] & b[349])^(a[203] & b[350])^(a[202] & b[351])^(a[201] & b[352])^(a[200] & b[353])^(a[199] & b[354])^(a[198] & b[355])^(a[197] & b[356])^(a[196] & b[357])^(a[195] & b[358])^(a[194] & b[359])^(a[193] & b[360])^(a[192] & b[361])^(a[191] & b[362])^(a[190] & b[363])^(a[189] & b[364])^(a[188] & b[365])^(a[187] & b[366])^(a[186] & b[367])^(a[185] & b[368])^(a[184] & b[369])^(a[183] & b[370])^(a[182] & b[371])^(a[181] & b[372])^(a[180] & b[373])^(a[179] & b[374])^(a[178] & b[375])^(a[177] & b[376])^(a[176] & b[377])^(a[175] & b[378])^(a[174] & b[379])^(a[173] & b[380])^(a[172] & b[381])^(a[171] & b[382])^(a[170] & b[383])^(a[169] & b[384])^(a[168] & b[385])^(a[167] & b[386])^(a[166] & b[387])^(a[165] & b[388])^(a[164] & b[389])^(a[163] & b[390])^(a[162] & b[391])^(a[161] & b[392])^(a[160] & b[393])^(a[159] & b[394])^(a[158] & b[395])^(a[157] & b[396])^(a[156] & b[397])^(a[155] & b[398])^(a[154] & b[399])^(a[153] & b[400])^(a[152] & b[401])^(a[151] & b[402])^(a[150] & b[403])^(a[149] & b[404])^(a[148] & b[405])^(a[147] & b[406])^(a[146] & b[407])^(a[145] & b[408]);
assign y[554] = (a[408] & b[146])^(a[407] & b[147])^(a[406] & b[148])^(a[405] & b[149])^(a[404] & b[150])^(a[403] & b[151])^(a[402] & b[152])^(a[401] & b[153])^(a[400] & b[154])^(a[399] & b[155])^(a[398] & b[156])^(a[397] & b[157])^(a[396] & b[158])^(a[395] & b[159])^(a[394] & b[160])^(a[393] & b[161])^(a[392] & b[162])^(a[391] & b[163])^(a[390] & b[164])^(a[389] & b[165])^(a[388] & b[166])^(a[387] & b[167])^(a[386] & b[168])^(a[385] & b[169])^(a[384] & b[170])^(a[383] & b[171])^(a[382] & b[172])^(a[381] & b[173])^(a[380] & b[174])^(a[379] & b[175])^(a[378] & b[176])^(a[377] & b[177])^(a[376] & b[178])^(a[375] & b[179])^(a[374] & b[180])^(a[373] & b[181])^(a[372] & b[182])^(a[371] & b[183])^(a[370] & b[184])^(a[369] & b[185])^(a[368] & b[186])^(a[367] & b[187])^(a[366] & b[188])^(a[365] & b[189])^(a[364] & b[190])^(a[363] & b[191])^(a[362] & b[192])^(a[361] & b[193])^(a[360] & b[194])^(a[359] & b[195])^(a[358] & b[196])^(a[357] & b[197])^(a[356] & b[198])^(a[355] & b[199])^(a[354] & b[200])^(a[353] & b[201])^(a[352] & b[202])^(a[351] & b[203])^(a[350] & b[204])^(a[349] & b[205])^(a[348] & b[206])^(a[347] & b[207])^(a[346] & b[208])^(a[345] & b[209])^(a[344] & b[210])^(a[343] & b[211])^(a[342] & b[212])^(a[341] & b[213])^(a[340] & b[214])^(a[339] & b[215])^(a[338] & b[216])^(a[337] & b[217])^(a[336] & b[218])^(a[335] & b[219])^(a[334] & b[220])^(a[333] & b[221])^(a[332] & b[222])^(a[331] & b[223])^(a[330] & b[224])^(a[329] & b[225])^(a[328] & b[226])^(a[327] & b[227])^(a[326] & b[228])^(a[325] & b[229])^(a[324] & b[230])^(a[323] & b[231])^(a[322] & b[232])^(a[321] & b[233])^(a[320] & b[234])^(a[319] & b[235])^(a[318] & b[236])^(a[317] & b[237])^(a[316] & b[238])^(a[315] & b[239])^(a[314] & b[240])^(a[313] & b[241])^(a[312] & b[242])^(a[311] & b[243])^(a[310] & b[244])^(a[309] & b[245])^(a[308] & b[246])^(a[307] & b[247])^(a[306] & b[248])^(a[305] & b[249])^(a[304] & b[250])^(a[303] & b[251])^(a[302] & b[252])^(a[301] & b[253])^(a[300] & b[254])^(a[299] & b[255])^(a[298] & b[256])^(a[297] & b[257])^(a[296] & b[258])^(a[295] & b[259])^(a[294] & b[260])^(a[293] & b[261])^(a[292] & b[262])^(a[291] & b[263])^(a[290] & b[264])^(a[289] & b[265])^(a[288] & b[266])^(a[287] & b[267])^(a[286] & b[268])^(a[285] & b[269])^(a[284] & b[270])^(a[283] & b[271])^(a[282] & b[272])^(a[281] & b[273])^(a[280] & b[274])^(a[279] & b[275])^(a[278] & b[276])^(a[277] & b[277])^(a[276] & b[278])^(a[275] & b[279])^(a[274] & b[280])^(a[273] & b[281])^(a[272] & b[282])^(a[271] & b[283])^(a[270] & b[284])^(a[269] & b[285])^(a[268] & b[286])^(a[267] & b[287])^(a[266] & b[288])^(a[265] & b[289])^(a[264] & b[290])^(a[263] & b[291])^(a[262] & b[292])^(a[261] & b[293])^(a[260] & b[294])^(a[259] & b[295])^(a[258] & b[296])^(a[257] & b[297])^(a[256] & b[298])^(a[255] & b[299])^(a[254] & b[300])^(a[253] & b[301])^(a[252] & b[302])^(a[251] & b[303])^(a[250] & b[304])^(a[249] & b[305])^(a[248] & b[306])^(a[247] & b[307])^(a[246] & b[308])^(a[245] & b[309])^(a[244] & b[310])^(a[243] & b[311])^(a[242] & b[312])^(a[241] & b[313])^(a[240] & b[314])^(a[239] & b[315])^(a[238] & b[316])^(a[237] & b[317])^(a[236] & b[318])^(a[235] & b[319])^(a[234] & b[320])^(a[233] & b[321])^(a[232] & b[322])^(a[231] & b[323])^(a[230] & b[324])^(a[229] & b[325])^(a[228] & b[326])^(a[227] & b[327])^(a[226] & b[328])^(a[225] & b[329])^(a[224] & b[330])^(a[223] & b[331])^(a[222] & b[332])^(a[221] & b[333])^(a[220] & b[334])^(a[219] & b[335])^(a[218] & b[336])^(a[217] & b[337])^(a[216] & b[338])^(a[215] & b[339])^(a[214] & b[340])^(a[213] & b[341])^(a[212] & b[342])^(a[211] & b[343])^(a[210] & b[344])^(a[209] & b[345])^(a[208] & b[346])^(a[207] & b[347])^(a[206] & b[348])^(a[205] & b[349])^(a[204] & b[350])^(a[203] & b[351])^(a[202] & b[352])^(a[201] & b[353])^(a[200] & b[354])^(a[199] & b[355])^(a[198] & b[356])^(a[197] & b[357])^(a[196] & b[358])^(a[195] & b[359])^(a[194] & b[360])^(a[193] & b[361])^(a[192] & b[362])^(a[191] & b[363])^(a[190] & b[364])^(a[189] & b[365])^(a[188] & b[366])^(a[187] & b[367])^(a[186] & b[368])^(a[185] & b[369])^(a[184] & b[370])^(a[183] & b[371])^(a[182] & b[372])^(a[181] & b[373])^(a[180] & b[374])^(a[179] & b[375])^(a[178] & b[376])^(a[177] & b[377])^(a[176] & b[378])^(a[175] & b[379])^(a[174] & b[380])^(a[173] & b[381])^(a[172] & b[382])^(a[171] & b[383])^(a[170] & b[384])^(a[169] & b[385])^(a[168] & b[386])^(a[167] & b[387])^(a[166] & b[388])^(a[165] & b[389])^(a[164] & b[390])^(a[163] & b[391])^(a[162] & b[392])^(a[161] & b[393])^(a[160] & b[394])^(a[159] & b[395])^(a[158] & b[396])^(a[157] & b[397])^(a[156] & b[398])^(a[155] & b[399])^(a[154] & b[400])^(a[153] & b[401])^(a[152] & b[402])^(a[151] & b[403])^(a[150] & b[404])^(a[149] & b[405])^(a[148] & b[406])^(a[147] & b[407])^(a[146] & b[408]);
assign y[555] = (a[408] & b[147])^(a[407] & b[148])^(a[406] & b[149])^(a[405] & b[150])^(a[404] & b[151])^(a[403] & b[152])^(a[402] & b[153])^(a[401] & b[154])^(a[400] & b[155])^(a[399] & b[156])^(a[398] & b[157])^(a[397] & b[158])^(a[396] & b[159])^(a[395] & b[160])^(a[394] & b[161])^(a[393] & b[162])^(a[392] & b[163])^(a[391] & b[164])^(a[390] & b[165])^(a[389] & b[166])^(a[388] & b[167])^(a[387] & b[168])^(a[386] & b[169])^(a[385] & b[170])^(a[384] & b[171])^(a[383] & b[172])^(a[382] & b[173])^(a[381] & b[174])^(a[380] & b[175])^(a[379] & b[176])^(a[378] & b[177])^(a[377] & b[178])^(a[376] & b[179])^(a[375] & b[180])^(a[374] & b[181])^(a[373] & b[182])^(a[372] & b[183])^(a[371] & b[184])^(a[370] & b[185])^(a[369] & b[186])^(a[368] & b[187])^(a[367] & b[188])^(a[366] & b[189])^(a[365] & b[190])^(a[364] & b[191])^(a[363] & b[192])^(a[362] & b[193])^(a[361] & b[194])^(a[360] & b[195])^(a[359] & b[196])^(a[358] & b[197])^(a[357] & b[198])^(a[356] & b[199])^(a[355] & b[200])^(a[354] & b[201])^(a[353] & b[202])^(a[352] & b[203])^(a[351] & b[204])^(a[350] & b[205])^(a[349] & b[206])^(a[348] & b[207])^(a[347] & b[208])^(a[346] & b[209])^(a[345] & b[210])^(a[344] & b[211])^(a[343] & b[212])^(a[342] & b[213])^(a[341] & b[214])^(a[340] & b[215])^(a[339] & b[216])^(a[338] & b[217])^(a[337] & b[218])^(a[336] & b[219])^(a[335] & b[220])^(a[334] & b[221])^(a[333] & b[222])^(a[332] & b[223])^(a[331] & b[224])^(a[330] & b[225])^(a[329] & b[226])^(a[328] & b[227])^(a[327] & b[228])^(a[326] & b[229])^(a[325] & b[230])^(a[324] & b[231])^(a[323] & b[232])^(a[322] & b[233])^(a[321] & b[234])^(a[320] & b[235])^(a[319] & b[236])^(a[318] & b[237])^(a[317] & b[238])^(a[316] & b[239])^(a[315] & b[240])^(a[314] & b[241])^(a[313] & b[242])^(a[312] & b[243])^(a[311] & b[244])^(a[310] & b[245])^(a[309] & b[246])^(a[308] & b[247])^(a[307] & b[248])^(a[306] & b[249])^(a[305] & b[250])^(a[304] & b[251])^(a[303] & b[252])^(a[302] & b[253])^(a[301] & b[254])^(a[300] & b[255])^(a[299] & b[256])^(a[298] & b[257])^(a[297] & b[258])^(a[296] & b[259])^(a[295] & b[260])^(a[294] & b[261])^(a[293] & b[262])^(a[292] & b[263])^(a[291] & b[264])^(a[290] & b[265])^(a[289] & b[266])^(a[288] & b[267])^(a[287] & b[268])^(a[286] & b[269])^(a[285] & b[270])^(a[284] & b[271])^(a[283] & b[272])^(a[282] & b[273])^(a[281] & b[274])^(a[280] & b[275])^(a[279] & b[276])^(a[278] & b[277])^(a[277] & b[278])^(a[276] & b[279])^(a[275] & b[280])^(a[274] & b[281])^(a[273] & b[282])^(a[272] & b[283])^(a[271] & b[284])^(a[270] & b[285])^(a[269] & b[286])^(a[268] & b[287])^(a[267] & b[288])^(a[266] & b[289])^(a[265] & b[290])^(a[264] & b[291])^(a[263] & b[292])^(a[262] & b[293])^(a[261] & b[294])^(a[260] & b[295])^(a[259] & b[296])^(a[258] & b[297])^(a[257] & b[298])^(a[256] & b[299])^(a[255] & b[300])^(a[254] & b[301])^(a[253] & b[302])^(a[252] & b[303])^(a[251] & b[304])^(a[250] & b[305])^(a[249] & b[306])^(a[248] & b[307])^(a[247] & b[308])^(a[246] & b[309])^(a[245] & b[310])^(a[244] & b[311])^(a[243] & b[312])^(a[242] & b[313])^(a[241] & b[314])^(a[240] & b[315])^(a[239] & b[316])^(a[238] & b[317])^(a[237] & b[318])^(a[236] & b[319])^(a[235] & b[320])^(a[234] & b[321])^(a[233] & b[322])^(a[232] & b[323])^(a[231] & b[324])^(a[230] & b[325])^(a[229] & b[326])^(a[228] & b[327])^(a[227] & b[328])^(a[226] & b[329])^(a[225] & b[330])^(a[224] & b[331])^(a[223] & b[332])^(a[222] & b[333])^(a[221] & b[334])^(a[220] & b[335])^(a[219] & b[336])^(a[218] & b[337])^(a[217] & b[338])^(a[216] & b[339])^(a[215] & b[340])^(a[214] & b[341])^(a[213] & b[342])^(a[212] & b[343])^(a[211] & b[344])^(a[210] & b[345])^(a[209] & b[346])^(a[208] & b[347])^(a[207] & b[348])^(a[206] & b[349])^(a[205] & b[350])^(a[204] & b[351])^(a[203] & b[352])^(a[202] & b[353])^(a[201] & b[354])^(a[200] & b[355])^(a[199] & b[356])^(a[198] & b[357])^(a[197] & b[358])^(a[196] & b[359])^(a[195] & b[360])^(a[194] & b[361])^(a[193] & b[362])^(a[192] & b[363])^(a[191] & b[364])^(a[190] & b[365])^(a[189] & b[366])^(a[188] & b[367])^(a[187] & b[368])^(a[186] & b[369])^(a[185] & b[370])^(a[184] & b[371])^(a[183] & b[372])^(a[182] & b[373])^(a[181] & b[374])^(a[180] & b[375])^(a[179] & b[376])^(a[178] & b[377])^(a[177] & b[378])^(a[176] & b[379])^(a[175] & b[380])^(a[174] & b[381])^(a[173] & b[382])^(a[172] & b[383])^(a[171] & b[384])^(a[170] & b[385])^(a[169] & b[386])^(a[168] & b[387])^(a[167] & b[388])^(a[166] & b[389])^(a[165] & b[390])^(a[164] & b[391])^(a[163] & b[392])^(a[162] & b[393])^(a[161] & b[394])^(a[160] & b[395])^(a[159] & b[396])^(a[158] & b[397])^(a[157] & b[398])^(a[156] & b[399])^(a[155] & b[400])^(a[154] & b[401])^(a[153] & b[402])^(a[152] & b[403])^(a[151] & b[404])^(a[150] & b[405])^(a[149] & b[406])^(a[148] & b[407])^(a[147] & b[408]);
assign y[556] = (a[408] & b[148])^(a[407] & b[149])^(a[406] & b[150])^(a[405] & b[151])^(a[404] & b[152])^(a[403] & b[153])^(a[402] & b[154])^(a[401] & b[155])^(a[400] & b[156])^(a[399] & b[157])^(a[398] & b[158])^(a[397] & b[159])^(a[396] & b[160])^(a[395] & b[161])^(a[394] & b[162])^(a[393] & b[163])^(a[392] & b[164])^(a[391] & b[165])^(a[390] & b[166])^(a[389] & b[167])^(a[388] & b[168])^(a[387] & b[169])^(a[386] & b[170])^(a[385] & b[171])^(a[384] & b[172])^(a[383] & b[173])^(a[382] & b[174])^(a[381] & b[175])^(a[380] & b[176])^(a[379] & b[177])^(a[378] & b[178])^(a[377] & b[179])^(a[376] & b[180])^(a[375] & b[181])^(a[374] & b[182])^(a[373] & b[183])^(a[372] & b[184])^(a[371] & b[185])^(a[370] & b[186])^(a[369] & b[187])^(a[368] & b[188])^(a[367] & b[189])^(a[366] & b[190])^(a[365] & b[191])^(a[364] & b[192])^(a[363] & b[193])^(a[362] & b[194])^(a[361] & b[195])^(a[360] & b[196])^(a[359] & b[197])^(a[358] & b[198])^(a[357] & b[199])^(a[356] & b[200])^(a[355] & b[201])^(a[354] & b[202])^(a[353] & b[203])^(a[352] & b[204])^(a[351] & b[205])^(a[350] & b[206])^(a[349] & b[207])^(a[348] & b[208])^(a[347] & b[209])^(a[346] & b[210])^(a[345] & b[211])^(a[344] & b[212])^(a[343] & b[213])^(a[342] & b[214])^(a[341] & b[215])^(a[340] & b[216])^(a[339] & b[217])^(a[338] & b[218])^(a[337] & b[219])^(a[336] & b[220])^(a[335] & b[221])^(a[334] & b[222])^(a[333] & b[223])^(a[332] & b[224])^(a[331] & b[225])^(a[330] & b[226])^(a[329] & b[227])^(a[328] & b[228])^(a[327] & b[229])^(a[326] & b[230])^(a[325] & b[231])^(a[324] & b[232])^(a[323] & b[233])^(a[322] & b[234])^(a[321] & b[235])^(a[320] & b[236])^(a[319] & b[237])^(a[318] & b[238])^(a[317] & b[239])^(a[316] & b[240])^(a[315] & b[241])^(a[314] & b[242])^(a[313] & b[243])^(a[312] & b[244])^(a[311] & b[245])^(a[310] & b[246])^(a[309] & b[247])^(a[308] & b[248])^(a[307] & b[249])^(a[306] & b[250])^(a[305] & b[251])^(a[304] & b[252])^(a[303] & b[253])^(a[302] & b[254])^(a[301] & b[255])^(a[300] & b[256])^(a[299] & b[257])^(a[298] & b[258])^(a[297] & b[259])^(a[296] & b[260])^(a[295] & b[261])^(a[294] & b[262])^(a[293] & b[263])^(a[292] & b[264])^(a[291] & b[265])^(a[290] & b[266])^(a[289] & b[267])^(a[288] & b[268])^(a[287] & b[269])^(a[286] & b[270])^(a[285] & b[271])^(a[284] & b[272])^(a[283] & b[273])^(a[282] & b[274])^(a[281] & b[275])^(a[280] & b[276])^(a[279] & b[277])^(a[278] & b[278])^(a[277] & b[279])^(a[276] & b[280])^(a[275] & b[281])^(a[274] & b[282])^(a[273] & b[283])^(a[272] & b[284])^(a[271] & b[285])^(a[270] & b[286])^(a[269] & b[287])^(a[268] & b[288])^(a[267] & b[289])^(a[266] & b[290])^(a[265] & b[291])^(a[264] & b[292])^(a[263] & b[293])^(a[262] & b[294])^(a[261] & b[295])^(a[260] & b[296])^(a[259] & b[297])^(a[258] & b[298])^(a[257] & b[299])^(a[256] & b[300])^(a[255] & b[301])^(a[254] & b[302])^(a[253] & b[303])^(a[252] & b[304])^(a[251] & b[305])^(a[250] & b[306])^(a[249] & b[307])^(a[248] & b[308])^(a[247] & b[309])^(a[246] & b[310])^(a[245] & b[311])^(a[244] & b[312])^(a[243] & b[313])^(a[242] & b[314])^(a[241] & b[315])^(a[240] & b[316])^(a[239] & b[317])^(a[238] & b[318])^(a[237] & b[319])^(a[236] & b[320])^(a[235] & b[321])^(a[234] & b[322])^(a[233] & b[323])^(a[232] & b[324])^(a[231] & b[325])^(a[230] & b[326])^(a[229] & b[327])^(a[228] & b[328])^(a[227] & b[329])^(a[226] & b[330])^(a[225] & b[331])^(a[224] & b[332])^(a[223] & b[333])^(a[222] & b[334])^(a[221] & b[335])^(a[220] & b[336])^(a[219] & b[337])^(a[218] & b[338])^(a[217] & b[339])^(a[216] & b[340])^(a[215] & b[341])^(a[214] & b[342])^(a[213] & b[343])^(a[212] & b[344])^(a[211] & b[345])^(a[210] & b[346])^(a[209] & b[347])^(a[208] & b[348])^(a[207] & b[349])^(a[206] & b[350])^(a[205] & b[351])^(a[204] & b[352])^(a[203] & b[353])^(a[202] & b[354])^(a[201] & b[355])^(a[200] & b[356])^(a[199] & b[357])^(a[198] & b[358])^(a[197] & b[359])^(a[196] & b[360])^(a[195] & b[361])^(a[194] & b[362])^(a[193] & b[363])^(a[192] & b[364])^(a[191] & b[365])^(a[190] & b[366])^(a[189] & b[367])^(a[188] & b[368])^(a[187] & b[369])^(a[186] & b[370])^(a[185] & b[371])^(a[184] & b[372])^(a[183] & b[373])^(a[182] & b[374])^(a[181] & b[375])^(a[180] & b[376])^(a[179] & b[377])^(a[178] & b[378])^(a[177] & b[379])^(a[176] & b[380])^(a[175] & b[381])^(a[174] & b[382])^(a[173] & b[383])^(a[172] & b[384])^(a[171] & b[385])^(a[170] & b[386])^(a[169] & b[387])^(a[168] & b[388])^(a[167] & b[389])^(a[166] & b[390])^(a[165] & b[391])^(a[164] & b[392])^(a[163] & b[393])^(a[162] & b[394])^(a[161] & b[395])^(a[160] & b[396])^(a[159] & b[397])^(a[158] & b[398])^(a[157] & b[399])^(a[156] & b[400])^(a[155] & b[401])^(a[154] & b[402])^(a[153] & b[403])^(a[152] & b[404])^(a[151] & b[405])^(a[150] & b[406])^(a[149] & b[407])^(a[148] & b[408]);
assign y[557] = (a[408] & b[149])^(a[407] & b[150])^(a[406] & b[151])^(a[405] & b[152])^(a[404] & b[153])^(a[403] & b[154])^(a[402] & b[155])^(a[401] & b[156])^(a[400] & b[157])^(a[399] & b[158])^(a[398] & b[159])^(a[397] & b[160])^(a[396] & b[161])^(a[395] & b[162])^(a[394] & b[163])^(a[393] & b[164])^(a[392] & b[165])^(a[391] & b[166])^(a[390] & b[167])^(a[389] & b[168])^(a[388] & b[169])^(a[387] & b[170])^(a[386] & b[171])^(a[385] & b[172])^(a[384] & b[173])^(a[383] & b[174])^(a[382] & b[175])^(a[381] & b[176])^(a[380] & b[177])^(a[379] & b[178])^(a[378] & b[179])^(a[377] & b[180])^(a[376] & b[181])^(a[375] & b[182])^(a[374] & b[183])^(a[373] & b[184])^(a[372] & b[185])^(a[371] & b[186])^(a[370] & b[187])^(a[369] & b[188])^(a[368] & b[189])^(a[367] & b[190])^(a[366] & b[191])^(a[365] & b[192])^(a[364] & b[193])^(a[363] & b[194])^(a[362] & b[195])^(a[361] & b[196])^(a[360] & b[197])^(a[359] & b[198])^(a[358] & b[199])^(a[357] & b[200])^(a[356] & b[201])^(a[355] & b[202])^(a[354] & b[203])^(a[353] & b[204])^(a[352] & b[205])^(a[351] & b[206])^(a[350] & b[207])^(a[349] & b[208])^(a[348] & b[209])^(a[347] & b[210])^(a[346] & b[211])^(a[345] & b[212])^(a[344] & b[213])^(a[343] & b[214])^(a[342] & b[215])^(a[341] & b[216])^(a[340] & b[217])^(a[339] & b[218])^(a[338] & b[219])^(a[337] & b[220])^(a[336] & b[221])^(a[335] & b[222])^(a[334] & b[223])^(a[333] & b[224])^(a[332] & b[225])^(a[331] & b[226])^(a[330] & b[227])^(a[329] & b[228])^(a[328] & b[229])^(a[327] & b[230])^(a[326] & b[231])^(a[325] & b[232])^(a[324] & b[233])^(a[323] & b[234])^(a[322] & b[235])^(a[321] & b[236])^(a[320] & b[237])^(a[319] & b[238])^(a[318] & b[239])^(a[317] & b[240])^(a[316] & b[241])^(a[315] & b[242])^(a[314] & b[243])^(a[313] & b[244])^(a[312] & b[245])^(a[311] & b[246])^(a[310] & b[247])^(a[309] & b[248])^(a[308] & b[249])^(a[307] & b[250])^(a[306] & b[251])^(a[305] & b[252])^(a[304] & b[253])^(a[303] & b[254])^(a[302] & b[255])^(a[301] & b[256])^(a[300] & b[257])^(a[299] & b[258])^(a[298] & b[259])^(a[297] & b[260])^(a[296] & b[261])^(a[295] & b[262])^(a[294] & b[263])^(a[293] & b[264])^(a[292] & b[265])^(a[291] & b[266])^(a[290] & b[267])^(a[289] & b[268])^(a[288] & b[269])^(a[287] & b[270])^(a[286] & b[271])^(a[285] & b[272])^(a[284] & b[273])^(a[283] & b[274])^(a[282] & b[275])^(a[281] & b[276])^(a[280] & b[277])^(a[279] & b[278])^(a[278] & b[279])^(a[277] & b[280])^(a[276] & b[281])^(a[275] & b[282])^(a[274] & b[283])^(a[273] & b[284])^(a[272] & b[285])^(a[271] & b[286])^(a[270] & b[287])^(a[269] & b[288])^(a[268] & b[289])^(a[267] & b[290])^(a[266] & b[291])^(a[265] & b[292])^(a[264] & b[293])^(a[263] & b[294])^(a[262] & b[295])^(a[261] & b[296])^(a[260] & b[297])^(a[259] & b[298])^(a[258] & b[299])^(a[257] & b[300])^(a[256] & b[301])^(a[255] & b[302])^(a[254] & b[303])^(a[253] & b[304])^(a[252] & b[305])^(a[251] & b[306])^(a[250] & b[307])^(a[249] & b[308])^(a[248] & b[309])^(a[247] & b[310])^(a[246] & b[311])^(a[245] & b[312])^(a[244] & b[313])^(a[243] & b[314])^(a[242] & b[315])^(a[241] & b[316])^(a[240] & b[317])^(a[239] & b[318])^(a[238] & b[319])^(a[237] & b[320])^(a[236] & b[321])^(a[235] & b[322])^(a[234] & b[323])^(a[233] & b[324])^(a[232] & b[325])^(a[231] & b[326])^(a[230] & b[327])^(a[229] & b[328])^(a[228] & b[329])^(a[227] & b[330])^(a[226] & b[331])^(a[225] & b[332])^(a[224] & b[333])^(a[223] & b[334])^(a[222] & b[335])^(a[221] & b[336])^(a[220] & b[337])^(a[219] & b[338])^(a[218] & b[339])^(a[217] & b[340])^(a[216] & b[341])^(a[215] & b[342])^(a[214] & b[343])^(a[213] & b[344])^(a[212] & b[345])^(a[211] & b[346])^(a[210] & b[347])^(a[209] & b[348])^(a[208] & b[349])^(a[207] & b[350])^(a[206] & b[351])^(a[205] & b[352])^(a[204] & b[353])^(a[203] & b[354])^(a[202] & b[355])^(a[201] & b[356])^(a[200] & b[357])^(a[199] & b[358])^(a[198] & b[359])^(a[197] & b[360])^(a[196] & b[361])^(a[195] & b[362])^(a[194] & b[363])^(a[193] & b[364])^(a[192] & b[365])^(a[191] & b[366])^(a[190] & b[367])^(a[189] & b[368])^(a[188] & b[369])^(a[187] & b[370])^(a[186] & b[371])^(a[185] & b[372])^(a[184] & b[373])^(a[183] & b[374])^(a[182] & b[375])^(a[181] & b[376])^(a[180] & b[377])^(a[179] & b[378])^(a[178] & b[379])^(a[177] & b[380])^(a[176] & b[381])^(a[175] & b[382])^(a[174] & b[383])^(a[173] & b[384])^(a[172] & b[385])^(a[171] & b[386])^(a[170] & b[387])^(a[169] & b[388])^(a[168] & b[389])^(a[167] & b[390])^(a[166] & b[391])^(a[165] & b[392])^(a[164] & b[393])^(a[163] & b[394])^(a[162] & b[395])^(a[161] & b[396])^(a[160] & b[397])^(a[159] & b[398])^(a[158] & b[399])^(a[157] & b[400])^(a[156] & b[401])^(a[155] & b[402])^(a[154] & b[403])^(a[153] & b[404])^(a[152] & b[405])^(a[151] & b[406])^(a[150] & b[407])^(a[149] & b[408]);
assign y[558] = (a[408] & b[150])^(a[407] & b[151])^(a[406] & b[152])^(a[405] & b[153])^(a[404] & b[154])^(a[403] & b[155])^(a[402] & b[156])^(a[401] & b[157])^(a[400] & b[158])^(a[399] & b[159])^(a[398] & b[160])^(a[397] & b[161])^(a[396] & b[162])^(a[395] & b[163])^(a[394] & b[164])^(a[393] & b[165])^(a[392] & b[166])^(a[391] & b[167])^(a[390] & b[168])^(a[389] & b[169])^(a[388] & b[170])^(a[387] & b[171])^(a[386] & b[172])^(a[385] & b[173])^(a[384] & b[174])^(a[383] & b[175])^(a[382] & b[176])^(a[381] & b[177])^(a[380] & b[178])^(a[379] & b[179])^(a[378] & b[180])^(a[377] & b[181])^(a[376] & b[182])^(a[375] & b[183])^(a[374] & b[184])^(a[373] & b[185])^(a[372] & b[186])^(a[371] & b[187])^(a[370] & b[188])^(a[369] & b[189])^(a[368] & b[190])^(a[367] & b[191])^(a[366] & b[192])^(a[365] & b[193])^(a[364] & b[194])^(a[363] & b[195])^(a[362] & b[196])^(a[361] & b[197])^(a[360] & b[198])^(a[359] & b[199])^(a[358] & b[200])^(a[357] & b[201])^(a[356] & b[202])^(a[355] & b[203])^(a[354] & b[204])^(a[353] & b[205])^(a[352] & b[206])^(a[351] & b[207])^(a[350] & b[208])^(a[349] & b[209])^(a[348] & b[210])^(a[347] & b[211])^(a[346] & b[212])^(a[345] & b[213])^(a[344] & b[214])^(a[343] & b[215])^(a[342] & b[216])^(a[341] & b[217])^(a[340] & b[218])^(a[339] & b[219])^(a[338] & b[220])^(a[337] & b[221])^(a[336] & b[222])^(a[335] & b[223])^(a[334] & b[224])^(a[333] & b[225])^(a[332] & b[226])^(a[331] & b[227])^(a[330] & b[228])^(a[329] & b[229])^(a[328] & b[230])^(a[327] & b[231])^(a[326] & b[232])^(a[325] & b[233])^(a[324] & b[234])^(a[323] & b[235])^(a[322] & b[236])^(a[321] & b[237])^(a[320] & b[238])^(a[319] & b[239])^(a[318] & b[240])^(a[317] & b[241])^(a[316] & b[242])^(a[315] & b[243])^(a[314] & b[244])^(a[313] & b[245])^(a[312] & b[246])^(a[311] & b[247])^(a[310] & b[248])^(a[309] & b[249])^(a[308] & b[250])^(a[307] & b[251])^(a[306] & b[252])^(a[305] & b[253])^(a[304] & b[254])^(a[303] & b[255])^(a[302] & b[256])^(a[301] & b[257])^(a[300] & b[258])^(a[299] & b[259])^(a[298] & b[260])^(a[297] & b[261])^(a[296] & b[262])^(a[295] & b[263])^(a[294] & b[264])^(a[293] & b[265])^(a[292] & b[266])^(a[291] & b[267])^(a[290] & b[268])^(a[289] & b[269])^(a[288] & b[270])^(a[287] & b[271])^(a[286] & b[272])^(a[285] & b[273])^(a[284] & b[274])^(a[283] & b[275])^(a[282] & b[276])^(a[281] & b[277])^(a[280] & b[278])^(a[279] & b[279])^(a[278] & b[280])^(a[277] & b[281])^(a[276] & b[282])^(a[275] & b[283])^(a[274] & b[284])^(a[273] & b[285])^(a[272] & b[286])^(a[271] & b[287])^(a[270] & b[288])^(a[269] & b[289])^(a[268] & b[290])^(a[267] & b[291])^(a[266] & b[292])^(a[265] & b[293])^(a[264] & b[294])^(a[263] & b[295])^(a[262] & b[296])^(a[261] & b[297])^(a[260] & b[298])^(a[259] & b[299])^(a[258] & b[300])^(a[257] & b[301])^(a[256] & b[302])^(a[255] & b[303])^(a[254] & b[304])^(a[253] & b[305])^(a[252] & b[306])^(a[251] & b[307])^(a[250] & b[308])^(a[249] & b[309])^(a[248] & b[310])^(a[247] & b[311])^(a[246] & b[312])^(a[245] & b[313])^(a[244] & b[314])^(a[243] & b[315])^(a[242] & b[316])^(a[241] & b[317])^(a[240] & b[318])^(a[239] & b[319])^(a[238] & b[320])^(a[237] & b[321])^(a[236] & b[322])^(a[235] & b[323])^(a[234] & b[324])^(a[233] & b[325])^(a[232] & b[326])^(a[231] & b[327])^(a[230] & b[328])^(a[229] & b[329])^(a[228] & b[330])^(a[227] & b[331])^(a[226] & b[332])^(a[225] & b[333])^(a[224] & b[334])^(a[223] & b[335])^(a[222] & b[336])^(a[221] & b[337])^(a[220] & b[338])^(a[219] & b[339])^(a[218] & b[340])^(a[217] & b[341])^(a[216] & b[342])^(a[215] & b[343])^(a[214] & b[344])^(a[213] & b[345])^(a[212] & b[346])^(a[211] & b[347])^(a[210] & b[348])^(a[209] & b[349])^(a[208] & b[350])^(a[207] & b[351])^(a[206] & b[352])^(a[205] & b[353])^(a[204] & b[354])^(a[203] & b[355])^(a[202] & b[356])^(a[201] & b[357])^(a[200] & b[358])^(a[199] & b[359])^(a[198] & b[360])^(a[197] & b[361])^(a[196] & b[362])^(a[195] & b[363])^(a[194] & b[364])^(a[193] & b[365])^(a[192] & b[366])^(a[191] & b[367])^(a[190] & b[368])^(a[189] & b[369])^(a[188] & b[370])^(a[187] & b[371])^(a[186] & b[372])^(a[185] & b[373])^(a[184] & b[374])^(a[183] & b[375])^(a[182] & b[376])^(a[181] & b[377])^(a[180] & b[378])^(a[179] & b[379])^(a[178] & b[380])^(a[177] & b[381])^(a[176] & b[382])^(a[175] & b[383])^(a[174] & b[384])^(a[173] & b[385])^(a[172] & b[386])^(a[171] & b[387])^(a[170] & b[388])^(a[169] & b[389])^(a[168] & b[390])^(a[167] & b[391])^(a[166] & b[392])^(a[165] & b[393])^(a[164] & b[394])^(a[163] & b[395])^(a[162] & b[396])^(a[161] & b[397])^(a[160] & b[398])^(a[159] & b[399])^(a[158] & b[400])^(a[157] & b[401])^(a[156] & b[402])^(a[155] & b[403])^(a[154] & b[404])^(a[153] & b[405])^(a[152] & b[406])^(a[151] & b[407])^(a[150] & b[408]);
assign y[559] = (a[408] & b[151])^(a[407] & b[152])^(a[406] & b[153])^(a[405] & b[154])^(a[404] & b[155])^(a[403] & b[156])^(a[402] & b[157])^(a[401] & b[158])^(a[400] & b[159])^(a[399] & b[160])^(a[398] & b[161])^(a[397] & b[162])^(a[396] & b[163])^(a[395] & b[164])^(a[394] & b[165])^(a[393] & b[166])^(a[392] & b[167])^(a[391] & b[168])^(a[390] & b[169])^(a[389] & b[170])^(a[388] & b[171])^(a[387] & b[172])^(a[386] & b[173])^(a[385] & b[174])^(a[384] & b[175])^(a[383] & b[176])^(a[382] & b[177])^(a[381] & b[178])^(a[380] & b[179])^(a[379] & b[180])^(a[378] & b[181])^(a[377] & b[182])^(a[376] & b[183])^(a[375] & b[184])^(a[374] & b[185])^(a[373] & b[186])^(a[372] & b[187])^(a[371] & b[188])^(a[370] & b[189])^(a[369] & b[190])^(a[368] & b[191])^(a[367] & b[192])^(a[366] & b[193])^(a[365] & b[194])^(a[364] & b[195])^(a[363] & b[196])^(a[362] & b[197])^(a[361] & b[198])^(a[360] & b[199])^(a[359] & b[200])^(a[358] & b[201])^(a[357] & b[202])^(a[356] & b[203])^(a[355] & b[204])^(a[354] & b[205])^(a[353] & b[206])^(a[352] & b[207])^(a[351] & b[208])^(a[350] & b[209])^(a[349] & b[210])^(a[348] & b[211])^(a[347] & b[212])^(a[346] & b[213])^(a[345] & b[214])^(a[344] & b[215])^(a[343] & b[216])^(a[342] & b[217])^(a[341] & b[218])^(a[340] & b[219])^(a[339] & b[220])^(a[338] & b[221])^(a[337] & b[222])^(a[336] & b[223])^(a[335] & b[224])^(a[334] & b[225])^(a[333] & b[226])^(a[332] & b[227])^(a[331] & b[228])^(a[330] & b[229])^(a[329] & b[230])^(a[328] & b[231])^(a[327] & b[232])^(a[326] & b[233])^(a[325] & b[234])^(a[324] & b[235])^(a[323] & b[236])^(a[322] & b[237])^(a[321] & b[238])^(a[320] & b[239])^(a[319] & b[240])^(a[318] & b[241])^(a[317] & b[242])^(a[316] & b[243])^(a[315] & b[244])^(a[314] & b[245])^(a[313] & b[246])^(a[312] & b[247])^(a[311] & b[248])^(a[310] & b[249])^(a[309] & b[250])^(a[308] & b[251])^(a[307] & b[252])^(a[306] & b[253])^(a[305] & b[254])^(a[304] & b[255])^(a[303] & b[256])^(a[302] & b[257])^(a[301] & b[258])^(a[300] & b[259])^(a[299] & b[260])^(a[298] & b[261])^(a[297] & b[262])^(a[296] & b[263])^(a[295] & b[264])^(a[294] & b[265])^(a[293] & b[266])^(a[292] & b[267])^(a[291] & b[268])^(a[290] & b[269])^(a[289] & b[270])^(a[288] & b[271])^(a[287] & b[272])^(a[286] & b[273])^(a[285] & b[274])^(a[284] & b[275])^(a[283] & b[276])^(a[282] & b[277])^(a[281] & b[278])^(a[280] & b[279])^(a[279] & b[280])^(a[278] & b[281])^(a[277] & b[282])^(a[276] & b[283])^(a[275] & b[284])^(a[274] & b[285])^(a[273] & b[286])^(a[272] & b[287])^(a[271] & b[288])^(a[270] & b[289])^(a[269] & b[290])^(a[268] & b[291])^(a[267] & b[292])^(a[266] & b[293])^(a[265] & b[294])^(a[264] & b[295])^(a[263] & b[296])^(a[262] & b[297])^(a[261] & b[298])^(a[260] & b[299])^(a[259] & b[300])^(a[258] & b[301])^(a[257] & b[302])^(a[256] & b[303])^(a[255] & b[304])^(a[254] & b[305])^(a[253] & b[306])^(a[252] & b[307])^(a[251] & b[308])^(a[250] & b[309])^(a[249] & b[310])^(a[248] & b[311])^(a[247] & b[312])^(a[246] & b[313])^(a[245] & b[314])^(a[244] & b[315])^(a[243] & b[316])^(a[242] & b[317])^(a[241] & b[318])^(a[240] & b[319])^(a[239] & b[320])^(a[238] & b[321])^(a[237] & b[322])^(a[236] & b[323])^(a[235] & b[324])^(a[234] & b[325])^(a[233] & b[326])^(a[232] & b[327])^(a[231] & b[328])^(a[230] & b[329])^(a[229] & b[330])^(a[228] & b[331])^(a[227] & b[332])^(a[226] & b[333])^(a[225] & b[334])^(a[224] & b[335])^(a[223] & b[336])^(a[222] & b[337])^(a[221] & b[338])^(a[220] & b[339])^(a[219] & b[340])^(a[218] & b[341])^(a[217] & b[342])^(a[216] & b[343])^(a[215] & b[344])^(a[214] & b[345])^(a[213] & b[346])^(a[212] & b[347])^(a[211] & b[348])^(a[210] & b[349])^(a[209] & b[350])^(a[208] & b[351])^(a[207] & b[352])^(a[206] & b[353])^(a[205] & b[354])^(a[204] & b[355])^(a[203] & b[356])^(a[202] & b[357])^(a[201] & b[358])^(a[200] & b[359])^(a[199] & b[360])^(a[198] & b[361])^(a[197] & b[362])^(a[196] & b[363])^(a[195] & b[364])^(a[194] & b[365])^(a[193] & b[366])^(a[192] & b[367])^(a[191] & b[368])^(a[190] & b[369])^(a[189] & b[370])^(a[188] & b[371])^(a[187] & b[372])^(a[186] & b[373])^(a[185] & b[374])^(a[184] & b[375])^(a[183] & b[376])^(a[182] & b[377])^(a[181] & b[378])^(a[180] & b[379])^(a[179] & b[380])^(a[178] & b[381])^(a[177] & b[382])^(a[176] & b[383])^(a[175] & b[384])^(a[174] & b[385])^(a[173] & b[386])^(a[172] & b[387])^(a[171] & b[388])^(a[170] & b[389])^(a[169] & b[390])^(a[168] & b[391])^(a[167] & b[392])^(a[166] & b[393])^(a[165] & b[394])^(a[164] & b[395])^(a[163] & b[396])^(a[162] & b[397])^(a[161] & b[398])^(a[160] & b[399])^(a[159] & b[400])^(a[158] & b[401])^(a[157] & b[402])^(a[156] & b[403])^(a[155] & b[404])^(a[154] & b[405])^(a[153] & b[406])^(a[152] & b[407])^(a[151] & b[408]);
assign y[560] = (a[408] & b[152])^(a[407] & b[153])^(a[406] & b[154])^(a[405] & b[155])^(a[404] & b[156])^(a[403] & b[157])^(a[402] & b[158])^(a[401] & b[159])^(a[400] & b[160])^(a[399] & b[161])^(a[398] & b[162])^(a[397] & b[163])^(a[396] & b[164])^(a[395] & b[165])^(a[394] & b[166])^(a[393] & b[167])^(a[392] & b[168])^(a[391] & b[169])^(a[390] & b[170])^(a[389] & b[171])^(a[388] & b[172])^(a[387] & b[173])^(a[386] & b[174])^(a[385] & b[175])^(a[384] & b[176])^(a[383] & b[177])^(a[382] & b[178])^(a[381] & b[179])^(a[380] & b[180])^(a[379] & b[181])^(a[378] & b[182])^(a[377] & b[183])^(a[376] & b[184])^(a[375] & b[185])^(a[374] & b[186])^(a[373] & b[187])^(a[372] & b[188])^(a[371] & b[189])^(a[370] & b[190])^(a[369] & b[191])^(a[368] & b[192])^(a[367] & b[193])^(a[366] & b[194])^(a[365] & b[195])^(a[364] & b[196])^(a[363] & b[197])^(a[362] & b[198])^(a[361] & b[199])^(a[360] & b[200])^(a[359] & b[201])^(a[358] & b[202])^(a[357] & b[203])^(a[356] & b[204])^(a[355] & b[205])^(a[354] & b[206])^(a[353] & b[207])^(a[352] & b[208])^(a[351] & b[209])^(a[350] & b[210])^(a[349] & b[211])^(a[348] & b[212])^(a[347] & b[213])^(a[346] & b[214])^(a[345] & b[215])^(a[344] & b[216])^(a[343] & b[217])^(a[342] & b[218])^(a[341] & b[219])^(a[340] & b[220])^(a[339] & b[221])^(a[338] & b[222])^(a[337] & b[223])^(a[336] & b[224])^(a[335] & b[225])^(a[334] & b[226])^(a[333] & b[227])^(a[332] & b[228])^(a[331] & b[229])^(a[330] & b[230])^(a[329] & b[231])^(a[328] & b[232])^(a[327] & b[233])^(a[326] & b[234])^(a[325] & b[235])^(a[324] & b[236])^(a[323] & b[237])^(a[322] & b[238])^(a[321] & b[239])^(a[320] & b[240])^(a[319] & b[241])^(a[318] & b[242])^(a[317] & b[243])^(a[316] & b[244])^(a[315] & b[245])^(a[314] & b[246])^(a[313] & b[247])^(a[312] & b[248])^(a[311] & b[249])^(a[310] & b[250])^(a[309] & b[251])^(a[308] & b[252])^(a[307] & b[253])^(a[306] & b[254])^(a[305] & b[255])^(a[304] & b[256])^(a[303] & b[257])^(a[302] & b[258])^(a[301] & b[259])^(a[300] & b[260])^(a[299] & b[261])^(a[298] & b[262])^(a[297] & b[263])^(a[296] & b[264])^(a[295] & b[265])^(a[294] & b[266])^(a[293] & b[267])^(a[292] & b[268])^(a[291] & b[269])^(a[290] & b[270])^(a[289] & b[271])^(a[288] & b[272])^(a[287] & b[273])^(a[286] & b[274])^(a[285] & b[275])^(a[284] & b[276])^(a[283] & b[277])^(a[282] & b[278])^(a[281] & b[279])^(a[280] & b[280])^(a[279] & b[281])^(a[278] & b[282])^(a[277] & b[283])^(a[276] & b[284])^(a[275] & b[285])^(a[274] & b[286])^(a[273] & b[287])^(a[272] & b[288])^(a[271] & b[289])^(a[270] & b[290])^(a[269] & b[291])^(a[268] & b[292])^(a[267] & b[293])^(a[266] & b[294])^(a[265] & b[295])^(a[264] & b[296])^(a[263] & b[297])^(a[262] & b[298])^(a[261] & b[299])^(a[260] & b[300])^(a[259] & b[301])^(a[258] & b[302])^(a[257] & b[303])^(a[256] & b[304])^(a[255] & b[305])^(a[254] & b[306])^(a[253] & b[307])^(a[252] & b[308])^(a[251] & b[309])^(a[250] & b[310])^(a[249] & b[311])^(a[248] & b[312])^(a[247] & b[313])^(a[246] & b[314])^(a[245] & b[315])^(a[244] & b[316])^(a[243] & b[317])^(a[242] & b[318])^(a[241] & b[319])^(a[240] & b[320])^(a[239] & b[321])^(a[238] & b[322])^(a[237] & b[323])^(a[236] & b[324])^(a[235] & b[325])^(a[234] & b[326])^(a[233] & b[327])^(a[232] & b[328])^(a[231] & b[329])^(a[230] & b[330])^(a[229] & b[331])^(a[228] & b[332])^(a[227] & b[333])^(a[226] & b[334])^(a[225] & b[335])^(a[224] & b[336])^(a[223] & b[337])^(a[222] & b[338])^(a[221] & b[339])^(a[220] & b[340])^(a[219] & b[341])^(a[218] & b[342])^(a[217] & b[343])^(a[216] & b[344])^(a[215] & b[345])^(a[214] & b[346])^(a[213] & b[347])^(a[212] & b[348])^(a[211] & b[349])^(a[210] & b[350])^(a[209] & b[351])^(a[208] & b[352])^(a[207] & b[353])^(a[206] & b[354])^(a[205] & b[355])^(a[204] & b[356])^(a[203] & b[357])^(a[202] & b[358])^(a[201] & b[359])^(a[200] & b[360])^(a[199] & b[361])^(a[198] & b[362])^(a[197] & b[363])^(a[196] & b[364])^(a[195] & b[365])^(a[194] & b[366])^(a[193] & b[367])^(a[192] & b[368])^(a[191] & b[369])^(a[190] & b[370])^(a[189] & b[371])^(a[188] & b[372])^(a[187] & b[373])^(a[186] & b[374])^(a[185] & b[375])^(a[184] & b[376])^(a[183] & b[377])^(a[182] & b[378])^(a[181] & b[379])^(a[180] & b[380])^(a[179] & b[381])^(a[178] & b[382])^(a[177] & b[383])^(a[176] & b[384])^(a[175] & b[385])^(a[174] & b[386])^(a[173] & b[387])^(a[172] & b[388])^(a[171] & b[389])^(a[170] & b[390])^(a[169] & b[391])^(a[168] & b[392])^(a[167] & b[393])^(a[166] & b[394])^(a[165] & b[395])^(a[164] & b[396])^(a[163] & b[397])^(a[162] & b[398])^(a[161] & b[399])^(a[160] & b[400])^(a[159] & b[401])^(a[158] & b[402])^(a[157] & b[403])^(a[156] & b[404])^(a[155] & b[405])^(a[154] & b[406])^(a[153] & b[407])^(a[152] & b[408]);
assign y[561] = (a[408] & b[153])^(a[407] & b[154])^(a[406] & b[155])^(a[405] & b[156])^(a[404] & b[157])^(a[403] & b[158])^(a[402] & b[159])^(a[401] & b[160])^(a[400] & b[161])^(a[399] & b[162])^(a[398] & b[163])^(a[397] & b[164])^(a[396] & b[165])^(a[395] & b[166])^(a[394] & b[167])^(a[393] & b[168])^(a[392] & b[169])^(a[391] & b[170])^(a[390] & b[171])^(a[389] & b[172])^(a[388] & b[173])^(a[387] & b[174])^(a[386] & b[175])^(a[385] & b[176])^(a[384] & b[177])^(a[383] & b[178])^(a[382] & b[179])^(a[381] & b[180])^(a[380] & b[181])^(a[379] & b[182])^(a[378] & b[183])^(a[377] & b[184])^(a[376] & b[185])^(a[375] & b[186])^(a[374] & b[187])^(a[373] & b[188])^(a[372] & b[189])^(a[371] & b[190])^(a[370] & b[191])^(a[369] & b[192])^(a[368] & b[193])^(a[367] & b[194])^(a[366] & b[195])^(a[365] & b[196])^(a[364] & b[197])^(a[363] & b[198])^(a[362] & b[199])^(a[361] & b[200])^(a[360] & b[201])^(a[359] & b[202])^(a[358] & b[203])^(a[357] & b[204])^(a[356] & b[205])^(a[355] & b[206])^(a[354] & b[207])^(a[353] & b[208])^(a[352] & b[209])^(a[351] & b[210])^(a[350] & b[211])^(a[349] & b[212])^(a[348] & b[213])^(a[347] & b[214])^(a[346] & b[215])^(a[345] & b[216])^(a[344] & b[217])^(a[343] & b[218])^(a[342] & b[219])^(a[341] & b[220])^(a[340] & b[221])^(a[339] & b[222])^(a[338] & b[223])^(a[337] & b[224])^(a[336] & b[225])^(a[335] & b[226])^(a[334] & b[227])^(a[333] & b[228])^(a[332] & b[229])^(a[331] & b[230])^(a[330] & b[231])^(a[329] & b[232])^(a[328] & b[233])^(a[327] & b[234])^(a[326] & b[235])^(a[325] & b[236])^(a[324] & b[237])^(a[323] & b[238])^(a[322] & b[239])^(a[321] & b[240])^(a[320] & b[241])^(a[319] & b[242])^(a[318] & b[243])^(a[317] & b[244])^(a[316] & b[245])^(a[315] & b[246])^(a[314] & b[247])^(a[313] & b[248])^(a[312] & b[249])^(a[311] & b[250])^(a[310] & b[251])^(a[309] & b[252])^(a[308] & b[253])^(a[307] & b[254])^(a[306] & b[255])^(a[305] & b[256])^(a[304] & b[257])^(a[303] & b[258])^(a[302] & b[259])^(a[301] & b[260])^(a[300] & b[261])^(a[299] & b[262])^(a[298] & b[263])^(a[297] & b[264])^(a[296] & b[265])^(a[295] & b[266])^(a[294] & b[267])^(a[293] & b[268])^(a[292] & b[269])^(a[291] & b[270])^(a[290] & b[271])^(a[289] & b[272])^(a[288] & b[273])^(a[287] & b[274])^(a[286] & b[275])^(a[285] & b[276])^(a[284] & b[277])^(a[283] & b[278])^(a[282] & b[279])^(a[281] & b[280])^(a[280] & b[281])^(a[279] & b[282])^(a[278] & b[283])^(a[277] & b[284])^(a[276] & b[285])^(a[275] & b[286])^(a[274] & b[287])^(a[273] & b[288])^(a[272] & b[289])^(a[271] & b[290])^(a[270] & b[291])^(a[269] & b[292])^(a[268] & b[293])^(a[267] & b[294])^(a[266] & b[295])^(a[265] & b[296])^(a[264] & b[297])^(a[263] & b[298])^(a[262] & b[299])^(a[261] & b[300])^(a[260] & b[301])^(a[259] & b[302])^(a[258] & b[303])^(a[257] & b[304])^(a[256] & b[305])^(a[255] & b[306])^(a[254] & b[307])^(a[253] & b[308])^(a[252] & b[309])^(a[251] & b[310])^(a[250] & b[311])^(a[249] & b[312])^(a[248] & b[313])^(a[247] & b[314])^(a[246] & b[315])^(a[245] & b[316])^(a[244] & b[317])^(a[243] & b[318])^(a[242] & b[319])^(a[241] & b[320])^(a[240] & b[321])^(a[239] & b[322])^(a[238] & b[323])^(a[237] & b[324])^(a[236] & b[325])^(a[235] & b[326])^(a[234] & b[327])^(a[233] & b[328])^(a[232] & b[329])^(a[231] & b[330])^(a[230] & b[331])^(a[229] & b[332])^(a[228] & b[333])^(a[227] & b[334])^(a[226] & b[335])^(a[225] & b[336])^(a[224] & b[337])^(a[223] & b[338])^(a[222] & b[339])^(a[221] & b[340])^(a[220] & b[341])^(a[219] & b[342])^(a[218] & b[343])^(a[217] & b[344])^(a[216] & b[345])^(a[215] & b[346])^(a[214] & b[347])^(a[213] & b[348])^(a[212] & b[349])^(a[211] & b[350])^(a[210] & b[351])^(a[209] & b[352])^(a[208] & b[353])^(a[207] & b[354])^(a[206] & b[355])^(a[205] & b[356])^(a[204] & b[357])^(a[203] & b[358])^(a[202] & b[359])^(a[201] & b[360])^(a[200] & b[361])^(a[199] & b[362])^(a[198] & b[363])^(a[197] & b[364])^(a[196] & b[365])^(a[195] & b[366])^(a[194] & b[367])^(a[193] & b[368])^(a[192] & b[369])^(a[191] & b[370])^(a[190] & b[371])^(a[189] & b[372])^(a[188] & b[373])^(a[187] & b[374])^(a[186] & b[375])^(a[185] & b[376])^(a[184] & b[377])^(a[183] & b[378])^(a[182] & b[379])^(a[181] & b[380])^(a[180] & b[381])^(a[179] & b[382])^(a[178] & b[383])^(a[177] & b[384])^(a[176] & b[385])^(a[175] & b[386])^(a[174] & b[387])^(a[173] & b[388])^(a[172] & b[389])^(a[171] & b[390])^(a[170] & b[391])^(a[169] & b[392])^(a[168] & b[393])^(a[167] & b[394])^(a[166] & b[395])^(a[165] & b[396])^(a[164] & b[397])^(a[163] & b[398])^(a[162] & b[399])^(a[161] & b[400])^(a[160] & b[401])^(a[159] & b[402])^(a[158] & b[403])^(a[157] & b[404])^(a[156] & b[405])^(a[155] & b[406])^(a[154] & b[407])^(a[153] & b[408]);
assign y[562] = (a[408] & b[154])^(a[407] & b[155])^(a[406] & b[156])^(a[405] & b[157])^(a[404] & b[158])^(a[403] & b[159])^(a[402] & b[160])^(a[401] & b[161])^(a[400] & b[162])^(a[399] & b[163])^(a[398] & b[164])^(a[397] & b[165])^(a[396] & b[166])^(a[395] & b[167])^(a[394] & b[168])^(a[393] & b[169])^(a[392] & b[170])^(a[391] & b[171])^(a[390] & b[172])^(a[389] & b[173])^(a[388] & b[174])^(a[387] & b[175])^(a[386] & b[176])^(a[385] & b[177])^(a[384] & b[178])^(a[383] & b[179])^(a[382] & b[180])^(a[381] & b[181])^(a[380] & b[182])^(a[379] & b[183])^(a[378] & b[184])^(a[377] & b[185])^(a[376] & b[186])^(a[375] & b[187])^(a[374] & b[188])^(a[373] & b[189])^(a[372] & b[190])^(a[371] & b[191])^(a[370] & b[192])^(a[369] & b[193])^(a[368] & b[194])^(a[367] & b[195])^(a[366] & b[196])^(a[365] & b[197])^(a[364] & b[198])^(a[363] & b[199])^(a[362] & b[200])^(a[361] & b[201])^(a[360] & b[202])^(a[359] & b[203])^(a[358] & b[204])^(a[357] & b[205])^(a[356] & b[206])^(a[355] & b[207])^(a[354] & b[208])^(a[353] & b[209])^(a[352] & b[210])^(a[351] & b[211])^(a[350] & b[212])^(a[349] & b[213])^(a[348] & b[214])^(a[347] & b[215])^(a[346] & b[216])^(a[345] & b[217])^(a[344] & b[218])^(a[343] & b[219])^(a[342] & b[220])^(a[341] & b[221])^(a[340] & b[222])^(a[339] & b[223])^(a[338] & b[224])^(a[337] & b[225])^(a[336] & b[226])^(a[335] & b[227])^(a[334] & b[228])^(a[333] & b[229])^(a[332] & b[230])^(a[331] & b[231])^(a[330] & b[232])^(a[329] & b[233])^(a[328] & b[234])^(a[327] & b[235])^(a[326] & b[236])^(a[325] & b[237])^(a[324] & b[238])^(a[323] & b[239])^(a[322] & b[240])^(a[321] & b[241])^(a[320] & b[242])^(a[319] & b[243])^(a[318] & b[244])^(a[317] & b[245])^(a[316] & b[246])^(a[315] & b[247])^(a[314] & b[248])^(a[313] & b[249])^(a[312] & b[250])^(a[311] & b[251])^(a[310] & b[252])^(a[309] & b[253])^(a[308] & b[254])^(a[307] & b[255])^(a[306] & b[256])^(a[305] & b[257])^(a[304] & b[258])^(a[303] & b[259])^(a[302] & b[260])^(a[301] & b[261])^(a[300] & b[262])^(a[299] & b[263])^(a[298] & b[264])^(a[297] & b[265])^(a[296] & b[266])^(a[295] & b[267])^(a[294] & b[268])^(a[293] & b[269])^(a[292] & b[270])^(a[291] & b[271])^(a[290] & b[272])^(a[289] & b[273])^(a[288] & b[274])^(a[287] & b[275])^(a[286] & b[276])^(a[285] & b[277])^(a[284] & b[278])^(a[283] & b[279])^(a[282] & b[280])^(a[281] & b[281])^(a[280] & b[282])^(a[279] & b[283])^(a[278] & b[284])^(a[277] & b[285])^(a[276] & b[286])^(a[275] & b[287])^(a[274] & b[288])^(a[273] & b[289])^(a[272] & b[290])^(a[271] & b[291])^(a[270] & b[292])^(a[269] & b[293])^(a[268] & b[294])^(a[267] & b[295])^(a[266] & b[296])^(a[265] & b[297])^(a[264] & b[298])^(a[263] & b[299])^(a[262] & b[300])^(a[261] & b[301])^(a[260] & b[302])^(a[259] & b[303])^(a[258] & b[304])^(a[257] & b[305])^(a[256] & b[306])^(a[255] & b[307])^(a[254] & b[308])^(a[253] & b[309])^(a[252] & b[310])^(a[251] & b[311])^(a[250] & b[312])^(a[249] & b[313])^(a[248] & b[314])^(a[247] & b[315])^(a[246] & b[316])^(a[245] & b[317])^(a[244] & b[318])^(a[243] & b[319])^(a[242] & b[320])^(a[241] & b[321])^(a[240] & b[322])^(a[239] & b[323])^(a[238] & b[324])^(a[237] & b[325])^(a[236] & b[326])^(a[235] & b[327])^(a[234] & b[328])^(a[233] & b[329])^(a[232] & b[330])^(a[231] & b[331])^(a[230] & b[332])^(a[229] & b[333])^(a[228] & b[334])^(a[227] & b[335])^(a[226] & b[336])^(a[225] & b[337])^(a[224] & b[338])^(a[223] & b[339])^(a[222] & b[340])^(a[221] & b[341])^(a[220] & b[342])^(a[219] & b[343])^(a[218] & b[344])^(a[217] & b[345])^(a[216] & b[346])^(a[215] & b[347])^(a[214] & b[348])^(a[213] & b[349])^(a[212] & b[350])^(a[211] & b[351])^(a[210] & b[352])^(a[209] & b[353])^(a[208] & b[354])^(a[207] & b[355])^(a[206] & b[356])^(a[205] & b[357])^(a[204] & b[358])^(a[203] & b[359])^(a[202] & b[360])^(a[201] & b[361])^(a[200] & b[362])^(a[199] & b[363])^(a[198] & b[364])^(a[197] & b[365])^(a[196] & b[366])^(a[195] & b[367])^(a[194] & b[368])^(a[193] & b[369])^(a[192] & b[370])^(a[191] & b[371])^(a[190] & b[372])^(a[189] & b[373])^(a[188] & b[374])^(a[187] & b[375])^(a[186] & b[376])^(a[185] & b[377])^(a[184] & b[378])^(a[183] & b[379])^(a[182] & b[380])^(a[181] & b[381])^(a[180] & b[382])^(a[179] & b[383])^(a[178] & b[384])^(a[177] & b[385])^(a[176] & b[386])^(a[175] & b[387])^(a[174] & b[388])^(a[173] & b[389])^(a[172] & b[390])^(a[171] & b[391])^(a[170] & b[392])^(a[169] & b[393])^(a[168] & b[394])^(a[167] & b[395])^(a[166] & b[396])^(a[165] & b[397])^(a[164] & b[398])^(a[163] & b[399])^(a[162] & b[400])^(a[161] & b[401])^(a[160] & b[402])^(a[159] & b[403])^(a[158] & b[404])^(a[157] & b[405])^(a[156] & b[406])^(a[155] & b[407])^(a[154] & b[408]);
assign y[563] = (a[408] & b[155])^(a[407] & b[156])^(a[406] & b[157])^(a[405] & b[158])^(a[404] & b[159])^(a[403] & b[160])^(a[402] & b[161])^(a[401] & b[162])^(a[400] & b[163])^(a[399] & b[164])^(a[398] & b[165])^(a[397] & b[166])^(a[396] & b[167])^(a[395] & b[168])^(a[394] & b[169])^(a[393] & b[170])^(a[392] & b[171])^(a[391] & b[172])^(a[390] & b[173])^(a[389] & b[174])^(a[388] & b[175])^(a[387] & b[176])^(a[386] & b[177])^(a[385] & b[178])^(a[384] & b[179])^(a[383] & b[180])^(a[382] & b[181])^(a[381] & b[182])^(a[380] & b[183])^(a[379] & b[184])^(a[378] & b[185])^(a[377] & b[186])^(a[376] & b[187])^(a[375] & b[188])^(a[374] & b[189])^(a[373] & b[190])^(a[372] & b[191])^(a[371] & b[192])^(a[370] & b[193])^(a[369] & b[194])^(a[368] & b[195])^(a[367] & b[196])^(a[366] & b[197])^(a[365] & b[198])^(a[364] & b[199])^(a[363] & b[200])^(a[362] & b[201])^(a[361] & b[202])^(a[360] & b[203])^(a[359] & b[204])^(a[358] & b[205])^(a[357] & b[206])^(a[356] & b[207])^(a[355] & b[208])^(a[354] & b[209])^(a[353] & b[210])^(a[352] & b[211])^(a[351] & b[212])^(a[350] & b[213])^(a[349] & b[214])^(a[348] & b[215])^(a[347] & b[216])^(a[346] & b[217])^(a[345] & b[218])^(a[344] & b[219])^(a[343] & b[220])^(a[342] & b[221])^(a[341] & b[222])^(a[340] & b[223])^(a[339] & b[224])^(a[338] & b[225])^(a[337] & b[226])^(a[336] & b[227])^(a[335] & b[228])^(a[334] & b[229])^(a[333] & b[230])^(a[332] & b[231])^(a[331] & b[232])^(a[330] & b[233])^(a[329] & b[234])^(a[328] & b[235])^(a[327] & b[236])^(a[326] & b[237])^(a[325] & b[238])^(a[324] & b[239])^(a[323] & b[240])^(a[322] & b[241])^(a[321] & b[242])^(a[320] & b[243])^(a[319] & b[244])^(a[318] & b[245])^(a[317] & b[246])^(a[316] & b[247])^(a[315] & b[248])^(a[314] & b[249])^(a[313] & b[250])^(a[312] & b[251])^(a[311] & b[252])^(a[310] & b[253])^(a[309] & b[254])^(a[308] & b[255])^(a[307] & b[256])^(a[306] & b[257])^(a[305] & b[258])^(a[304] & b[259])^(a[303] & b[260])^(a[302] & b[261])^(a[301] & b[262])^(a[300] & b[263])^(a[299] & b[264])^(a[298] & b[265])^(a[297] & b[266])^(a[296] & b[267])^(a[295] & b[268])^(a[294] & b[269])^(a[293] & b[270])^(a[292] & b[271])^(a[291] & b[272])^(a[290] & b[273])^(a[289] & b[274])^(a[288] & b[275])^(a[287] & b[276])^(a[286] & b[277])^(a[285] & b[278])^(a[284] & b[279])^(a[283] & b[280])^(a[282] & b[281])^(a[281] & b[282])^(a[280] & b[283])^(a[279] & b[284])^(a[278] & b[285])^(a[277] & b[286])^(a[276] & b[287])^(a[275] & b[288])^(a[274] & b[289])^(a[273] & b[290])^(a[272] & b[291])^(a[271] & b[292])^(a[270] & b[293])^(a[269] & b[294])^(a[268] & b[295])^(a[267] & b[296])^(a[266] & b[297])^(a[265] & b[298])^(a[264] & b[299])^(a[263] & b[300])^(a[262] & b[301])^(a[261] & b[302])^(a[260] & b[303])^(a[259] & b[304])^(a[258] & b[305])^(a[257] & b[306])^(a[256] & b[307])^(a[255] & b[308])^(a[254] & b[309])^(a[253] & b[310])^(a[252] & b[311])^(a[251] & b[312])^(a[250] & b[313])^(a[249] & b[314])^(a[248] & b[315])^(a[247] & b[316])^(a[246] & b[317])^(a[245] & b[318])^(a[244] & b[319])^(a[243] & b[320])^(a[242] & b[321])^(a[241] & b[322])^(a[240] & b[323])^(a[239] & b[324])^(a[238] & b[325])^(a[237] & b[326])^(a[236] & b[327])^(a[235] & b[328])^(a[234] & b[329])^(a[233] & b[330])^(a[232] & b[331])^(a[231] & b[332])^(a[230] & b[333])^(a[229] & b[334])^(a[228] & b[335])^(a[227] & b[336])^(a[226] & b[337])^(a[225] & b[338])^(a[224] & b[339])^(a[223] & b[340])^(a[222] & b[341])^(a[221] & b[342])^(a[220] & b[343])^(a[219] & b[344])^(a[218] & b[345])^(a[217] & b[346])^(a[216] & b[347])^(a[215] & b[348])^(a[214] & b[349])^(a[213] & b[350])^(a[212] & b[351])^(a[211] & b[352])^(a[210] & b[353])^(a[209] & b[354])^(a[208] & b[355])^(a[207] & b[356])^(a[206] & b[357])^(a[205] & b[358])^(a[204] & b[359])^(a[203] & b[360])^(a[202] & b[361])^(a[201] & b[362])^(a[200] & b[363])^(a[199] & b[364])^(a[198] & b[365])^(a[197] & b[366])^(a[196] & b[367])^(a[195] & b[368])^(a[194] & b[369])^(a[193] & b[370])^(a[192] & b[371])^(a[191] & b[372])^(a[190] & b[373])^(a[189] & b[374])^(a[188] & b[375])^(a[187] & b[376])^(a[186] & b[377])^(a[185] & b[378])^(a[184] & b[379])^(a[183] & b[380])^(a[182] & b[381])^(a[181] & b[382])^(a[180] & b[383])^(a[179] & b[384])^(a[178] & b[385])^(a[177] & b[386])^(a[176] & b[387])^(a[175] & b[388])^(a[174] & b[389])^(a[173] & b[390])^(a[172] & b[391])^(a[171] & b[392])^(a[170] & b[393])^(a[169] & b[394])^(a[168] & b[395])^(a[167] & b[396])^(a[166] & b[397])^(a[165] & b[398])^(a[164] & b[399])^(a[163] & b[400])^(a[162] & b[401])^(a[161] & b[402])^(a[160] & b[403])^(a[159] & b[404])^(a[158] & b[405])^(a[157] & b[406])^(a[156] & b[407])^(a[155] & b[408]);
assign y[564] = (a[408] & b[156])^(a[407] & b[157])^(a[406] & b[158])^(a[405] & b[159])^(a[404] & b[160])^(a[403] & b[161])^(a[402] & b[162])^(a[401] & b[163])^(a[400] & b[164])^(a[399] & b[165])^(a[398] & b[166])^(a[397] & b[167])^(a[396] & b[168])^(a[395] & b[169])^(a[394] & b[170])^(a[393] & b[171])^(a[392] & b[172])^(a[391] & b[173])^(a[390] & b[174])^(a[389] & b[175])^(a[388] & b[176])^(a[387] & b[177])^(a[386] & b[178])^(a[385] & b[179])^(a[384] & b[180])^(a[383] & b[181])^(a[382] & b[182])^(a[381] & b[183])^(a[380] & b[184])^(a[379] & b[185])^(a[378] & b[186])^(a[377] & b[187])^(a[376] & b[188])^(a[375] & b[189])^(a[374] & b[190])^(a[373] & b[191])^(a[372] & b[192])^(a[371] & b[193])^(a[370] & b[194])^(a[369] & b[195])^(a[368] & b[196])^(a[367] & b[197])^(a[366] & b[198])^(a[365] & b[199])^(a[364] & b[200])^(a[363] & b[201])^(a[362] & b[202])^(a[361] & b[203])^(a[360] & b[204])^(a[359] & b[205])^(a[358] & b[206])^(a[357] & b[207])^(a[356] & b[208])^(a[355] & b[209])^(a[354] & b[210])^(a[353] & b[211])^(a[352] & b[212])^(a[351] & b[213])^(a[350] & b[214])^(a[349] & b[215])^(a[348] & b[216])^(a[347] & b[217])^(a[346] & b[218])^(a[345] & b[219])^(a[344] & b[220])^(a[343] & b[221])^(a[342] & b[222])^(a[341] & b[223])^(a[340] & b[224])^(a[339] & b[225])^(a[338] & b[226])^(a[337] & b[227])^(a[336] & b[228])^(a[335] & b[229])^(a[334] & b[230])^(a[333] & b[231])^(a[332] & b[232])^(a[331] & b[233])^(a[330] & b[234])^(a[329] & b[235])^(a[328] & b[236])^(a[327] & b[237])^(a[326] & b[238])^(a[325] & b[239])^(a[324] & b[240])^(a[323] & b[241])^(a[322] & b[242])^(a[321] & b[243])^(a[320] & b[244])^(a[319] & b[245])^(a[318] & b[246])^(a[317] & b[247])^(a[316] & b[248])^(a[315] & b[249])^(a[314] & b[250])^(a[313] & b[251])^(a[312] & b[252])^(a[311] & b[253])^(a[310] & b[254])^(a[309] & b[255])^(a[308] & b[256])^(a[307] & b[257])^(a[306] & b[258])^(a[305] & b[259])^(a[304] & b[260])^(a[303] & b[261])^(a[302] & b[262])^(a[301] & b[263])^(a[300] & b[264])^(a[299] & b[265])^(a[298] & b[266])^(a[297] & b[267])^(a[296] & b[268])^(a[295] & b[269])^(a[294] & b[270])^(a[293] & b[271])^(a[292] & b[272])^(a[291] & b[273])^(a[290] & b[274])^(a[289] & b[275])^(a[288] & b[276])^(a[287] & b[277])^(a[286] & b[278])^(a[285] & b[279])^(a[284] & b[280])^(a[283] & b[281])^(a[282] & b[282])^(a[281] & b[283])^(a[280] & b[284])^(a[279] & b[285])^(a[278] & b[286])^(a[277] & b[287])^(a[276] & b[288])^(a[275] & b[289])^(a[274] & b[290])^(a[273] & b[291])^(a[272] & b[292])^(a[271] & b[293])^(a[270] & b[294])^(a[269] & b[295])^(a[268] & b[296])^(a[267] & b[297])^(a[266] & b[298])^(a[265] & b[299])^(a[264] & b[300])^(a[263] & b[301])^(a[262] & b[302])^(a[261] & b[303])^(a[260] & b[304])^(a[259] & b[305])^(a[258] & b[306])^(a[257] & b[307])^(a[256] & b[308])^(a[255] & b[309])^(a[254] & b[310])^(a[253] & b[311])^(a[252] & b[312])^(a[251] & b[313])^(a[250] & b[314])^(a[249] & b[315])^(a[248] & b[316])^(a[247] & b[317])^(a[246] & b[318])^(a[245] & b[319])^(a[244] & b[320])^(a[243] & b[321])^(a[242] & b[322])^(a[241] & b[323])^(a[240] & b[324])^(a[239] & b[325])^(a[238] & b[326])^(a[237] & b[327])^(a[236] & b[328])^(a[235] & b[329])^(a[234] & b[330])^(a[233] & b[331])^(a[232] & b[332])^(a[231] & b[333])^(a[230] & b[334])^(a[229] & b[335])^(a[228] & b[336])^(a[227] & b[337])^(a[226] & b[338])^(a[225] & b[339])^(a[224] & b[340])^(a[223] & b[341])^(a[222] & b[342])^(a[221] & b[343])^(a[220] & b[344])^(a[219] & b[345])^(a[218] & b[346])^(a[217] & b[347])^(a[216] & b[348])^(a[215] & b[349])^(a[214] & b[350])^(a[213] & b[351])^(a[212] & b[352])^(a[211] & b[353])^(a[210] & b[354])^(a[209] & b[355])^(a[208] & b[356])^(a[207] & b[357])^(a[206] & b[358])^(a[205] & b[359])^(a[204] & b[360])^(a[203] & b[361])^(a[202] & b[362])^(a[201] & b[363])^(a[200] & b[364])^(a[199] & b[365])^(a[198] & b[366])^(a[197] & b[367])^(a[196] & b[368])^(a[195] & b[369])^(a[194] & b[370])^(a[193] & b[371])^(a[192] & b[372])^(a[191] & b[373])^(a[190] & b[374])^(a[189] & b[375])^(a[188] & b[376])^(a[187] & b[377])^(a[186] & b[378])^(a[185] & b[379])^(a[184] & b[380])^(a[183] & b[381])^(a[182] & b[382])^(a[181] & b[383])^(a[180] & b[384])^(a[179] & b[385])^(a[178] & b[386])^(a[177] & b[387])^(a[176] & b[388])^(a[175] & b[389])^(a[174] & b[390])^(a[173] & b[391])^(a[172] & b[392])^(a[171] & b[393])^(a[170] & b[394])^(a[169] & b[395])^(a[168] & b[396])^(a[167] & b[397])^(a[166] & b[398])^(a[165] & b[399])^(a[164] & b[400])^(a[163] & b[401])^(a[162] & b[402])^(a[161] & b[403])^(a[160] & b[404])^(a[159] & b[405])^(a[158] & b[406])^(a[157] & b[407])^(a[156] & b[408]);
assign y[565] = (a[408] & b[157])^(a[407] & b[158])^(a[406] & b[159])^(a[405] & b[160])^(a[404] & b[161])^(a[403] & b[162])^(a[402] & b[163])^(a[401] & b[164])^(a[400] & b[165])^(a[399] & b[166])^(a[398] & b[167])^(a[397] & b[168])^(a[396] & b[169])^(a[395] & b[170])^(a[394] & b[171])^(a[393] & b[172])^(a[392] & b[173])^(a[391] & b[174])^(a[390] & b[175])^(a[389] & b[176])^(a[388] & b[177])^(a[387] & b[178])^(a[386] & b[179])^(a[385] & b[180])^(a[384] & b[181])^(a[383] & b[182])^(a[382] & b[183])^(a[381] & b[184])^(a[380] & b[185])^(a[379] & b[186])^(a[378] & b[187])^(a[377] & b[188])^(a[376] & b[189])^(a[375] & b[190])^(a[374] & b[191])^(a[373] & b[192])^(a[372] & b[193])^(a[371] & b[194])^(a[370] & b[195])^(a[369] & b[196])^(a[368] & b[197])^(a[367] & b[198])^(a[366] & b[199])^(a[365] & b[200])^(a[364] & b[201])^(a[363] & b[202])^(a[362] & b[203])^(a[361] & b[204])^(a[360] & b[205])^(a[359] & b[206])^(a[358] & b[207])^(a[357] & b[208])^(a[356] & b[209])^(a[355] & b[210])^(a[354] & b[211])^(a[353] & b[212])^(a[352] & b[213])^(a[351] & b[214])^(a[350] & b[215])^(a[349] & b[216])^(a[348] & b[217])^(a[347] & b[218])^(a[346] & b[219])^(a[345] & b[220])^(a[344] & b[221])^(a[343] & b[222])^(a[342] & b[223])^(a[341] & b[224])^(a[340] & b[225])^(a[339] & b[226])^(a[338] & b[227])^(a[337] & b[228])^(a[336] & b[229])^(a[335] & b[230])^(a[334] & b[231])^(a[333] & b[232])^(a[332] & b[233])^(a[331] & b[234])^(a[330] & b[235])^(a[329] & b[236])^(a[328] & b[237])^(a[327] & b[238])^(a[326] & b[239])^(a[325] & b[240])^(a[324] & b[241])^(a[323] & b[242])^(a[322] & b[243])^(a[321] & b[244])^(a[320] & b[245])^(a[319] & b[246])^(a[318] & b[247])^(a[317] & b[248])^(a[316] & b[249])^(a[315] & b[250])^(a[314] & b[251])^(a[313] & b[252])^(a[312] & b[253])^(a[311] & b[254])^(a[310] & b[255])^(a[309] & b[256])^(a[308] & b[257])^(a[307] & b[258])^(a[306] & b[259])^(a[305] & b[260])^(a[304] & b[261])^(a[303] & b[262])^(a[302] & b[263])^(a[301] & b[264])^(a[300] & b[265])^(a[299] & b[266])^(a[298] & b[267])^(a[297] & b[268])^(a[296] & b[269])^(a[295] & b[270])^(a[294] & b[271])^(a[293] & b[272])^(a[292] & b[273])^(a[291] & b[274])^(a[290] & b[275])^(a[289] & b[276])^(a[288] & b[277])^(a[287] & b[278])^(a[286] & b[279])^(a[285] & b[280])^(a[284] & b[281])^(a[283] & b[282])^(a[282] & b[283])^(a[281] & b[284])^(a[280] & b[285])^(a[279] & b[286])^(a[278] & b[287])^(a[277] & b[288])^(a[276] & b[289])^(a[275] & b[290])^(a[274] & b[291])^(a[273] & b[292])^(a[272] & b[293])^(a[271] & b[294])^(a[270] & b[295])^(a[269] & b[296])^(a[268] & b[297])^(a[267] & b[298])^(a[266] & b[299])^(a[265] & b[300])^(a[264] & b[301])^(a[263] & b[302])^(a[262] & b[303])^(a[261] & b[304])^(a[260] & b[305])^(a[259] & b[306])^(a[258] & b[307])^(a[257] & b[308])^(a[256] & b[309])^(a[255] & b[310])^(a[254] & b[311])^(a[253] & b[312])^(a[252] & b[313])^(a[251] & b[314])^(a[250] & b[315])^(a[249] & b[316])^(a[248] & b[317])^(a[247] & b[318])^(a[246] & b[319])^(a[245] & b[320])^(a[244] & b[321])^(a[243] & b[322])^(a[242] & b[323])^(a[241] & b[324])^(a[240] & b[325])^(a[239] & b[326])^(a[238] & b[327])^(a[237] & b[328])^(a[236] & b[329])^(a[235] & b[330])^(a[234] & b[331])^(a[233] & b[332])^(a[232] & b[333])^(a[231] & b[334])^(a[230] & b[335])^(a[229] & b[336])^(a[228] & b[337])^(a[227] & b[338])^(a[226] & b[339])^(a[225] & b[340])^(a[224] & b[341])^(a[223] & b[342])^(a[222] & b[343])^(a[221] & b[344])^(a[220] & b[345])^(a[219] & b[346])^(a[218] & b[347])^(a[217] & b[348])^(a[216] & b[349])^(a[215] & b[350])^(a[214] & b[351])^(a[213] & b[352])^(a[212] & b[353])^(a[211] & b[354])^(a[210] & b[355])^(a[209] & b[356])^(a[208] & b[357])^(a[207] & b[358])^(a[206] & b[359])^(a[205] & b[360])^(a[204] & b[361])^(a[203] & b[362])^(a[202] & b[363])^(a[201] & b[364])^(a[200] & b[365])^(a[199] & b[366])^(a[198] & b[367])^(a[197] & b[368])^(a[196] & b[369])^(a[195] & b[370])^(a[194] & b[371])^(a[193] & b[372])^(a[192] & b[373])^(a[191] & b[374])^(a[190] & b[375])^(a[189] & b[376])^(a[188] & b[377])^(a[187] & b[378])^(a[186] & b[379])^(a[185] & b[380])^(a[184] & b[381])^(a[183] & b[382])^(a[182] & b[383])^(a[181] & b[384])^(a[180] & b[385])^(a[179] & b[386])^(a[178] & b[387])^(a[177] & b[388])^(a[176] & b[389])^(a[175] & b[390])^(a[174] & b[391])^(a[173] & b[392])^(a[172] & b[393])^(a[171] & b[394])^(a[170] & b[395])^(a[169] & b[396])^(a[168] & b[397])^(a[167] & b[398])^(a[166] & b[399])^(a[165] & b[400])^(a[164] & b[401])^(a[163] & b[402])^(a[162] & b[403])^(a[161] & b[404])^(a[160] & b[405])^(a[159] & b[406])^(a[158] & b[407])^(a[157] & b[408]);
assign y[566] = (a[408] & b[158])^(a[407] & b[159])^(a[406] & b[160])^(a[405] & b[161])^(a[404] & b[162])^(a[403] & b[163])^(a[402] & b[164])^(a[401] & b[165])^(a[400] & b[166])^(a[399] & b[167])^(a[398] & b[168])^(a[397] & b[169])^(a[396] & b[170])^(a[395] & b[171])^(a[394] & b[172])^(a[393] & b[173])^(a[392] & b[174])^(a[391] & b[175])^(a[390] & b[176])^(a[389] & b[177])^(a[388] & b[178])^(a[387] & b[179])^(a[386] & b[180])^(a[385] & b[181])^(a[384] & b[182])^(a[383] & b[183])^(a[382] & b[184])^(a[381] & b[185])^(a[380] & b[186])^(a[379] & b[187])^(a[378] & b[188])^(a[377] & b[189])^(a[376] & b[190])^(a[375] & b[191])^(a[374] & b[192])^(a[373] & b[193])^(a[372] & b[194])^(a[371] & b[195])^(a[370] & b[196])^(a[369] & b[197])^(a[368] & b[198])^(a[367] & b[199])^(a[366] & b[200])^(a[365] & b[201])^(a[364] & b[202])^(a[363] & b[203])^(a[362] & b[204])^(a[361] & b[205])^(a[360] & b[206])^(a[359] & b[207])^(a[358] & b[208])^(a[357] & b[209])^(a[356] & b[210])^(a[355] & b[211])^(a[354] & b[212])^(a[353] & b[213])^(a[352] & b[214])^(a[351] & b[215])^(a[350] & b[216])^(a[349] & b[217])^(a[348] & b[218])^(a[347] & b[219])^(a[346] & b[220])^(a[345] & b[221])^(a[344] & b[222])^(a[343] & b[223])^(a[342] & b[224])^(a[341] & b[225])^(a[340] & b[226])^(a[339] & b[227])^(a[338] & b[228])^(a[337] & b[229])^(a[336] & b[230])^(a[335] & b[231])^(a[334] & b[232])^(a[333] & b[233])^(a[332] & b[234])^(a[331] & b[235])^(a[330] & b[236])^(a[329] & b[237])^(a[328] & b[238])^(a[327] & b[239])^(a[326] & b[240])^(a[325] & b[241])^(a[324] & b[242])^(a[323] & b[243])^(a[322] & b[244])^(a[321] & b[245])^(a[320] & b[246])^(a[319] & b[247])^(a[318] & b[248])^(a[317] & b[249])^(a[316] & b[250])^(a[315] & b[251])^(a[314] & b[252])^(a[313] & b[253])^(a[312] & b[254])^(a[311] & b[255])^(a[310] & b[256])^(a[309] & b[257])^(a[308] & b[258])^(a[307] & b[259])^(a[306] & b[260])^(a[305] & b[261])^(a[304] & b[262])^(a[303] & b[263])^(a[302] & b[264])^(a[301] & b[265])^(a[300] & b[266])^(a[299] & b[267])^(a[298] & b[268])^(a[297] & b[269])^(a[296] & b[270])^(a[295] & b[271])^(a[294] & b[272])^(a[293] & b[273])^(a[292] & b[274])^(a[291] & b[275])^(a[290] & b[276])^(a[289] & b[277])^(a[288] & b[278])^(a[287] & b[279])^(a[286] & b[280])^(a[285] & b[281])^(a[284] & b[282])^(a[283] & b[283])^(a[282] & b[284])^(a[281] & b[285])^(a[280] & b[286])^(a[279] & b[287])^(a[278] & b[288])^(a[277] & b[289])^(a[276] & b[290])^(a[275] & b[291])^(a[274] & b[292])^(a[273] & b[293])^(a[272] & b[294])^(a[271] & b[295])^(a[270] & b[296])^(a[269] & b[297])^(a[268] & b[298])^(a[267] & b[299])^(a[266] & b[300])^(a[265] & b[301])^(a[264] & b[302])^(a[263] & b[303])^(a[262] & b[304])^(a[261] & b[305])^(a[260] & b[306])^(a[259] & b[307])^(a[258] & b[308])^(a[257] & b[309])^(a[256] & b[310])^(a[255] & b[311])^(a[254] & b[312])^(a[253] & b[313])^(a[252] & b[314])^(a[251] & b[315])^(a[250] & b[316])^(a[249] & b[317])^(a[248] & b[318])^(a[247] & b[319])^(a[246] & b[320])^(a[245] & b[321])^(a[244] & b[322])^(a[243] & b[323])^(a[242] & b[324])^(a[241] & b[325])^(a[240] & b[326])^(a[239] & b[327])^(a[238] & b[328])^(a[237] & b[329])^(a[236] & b[330])^(a[235] & b[331])^(a[234] & b[332])^(a[233] & b[333])^(a[232] & b[334])^(a[231] & b[335])^(a[230] & b[336])^(a[229] & b[337])^(a[228] & b[338])^(a[227] & b[339])^(a[226] & b[340])^(a[225] & b[341])^(a[224] & b[342])^(a[223] & b[343])^(a[222] & b[344])^(a[221] & b[345])^(a[220] & b[346])^(a[219] & b[347])^(a[218] & b[348])^(a[217] & b[349])^(a[216] & b[350])^(a[215] & b[351])^(a[214] & b[352])^(a[213] & b[353])^(a[212] & b[354])^(a[211] & b[355])^(a[210] & b[356])^(a[209] & b[357])^(a[208] & b[358])^(a[207] & b[359])^(a[206] & b[360])^(a[205] & b[361])^(a[204] & b[362])^(a[203] & b[363])^(a[202] & b[364])^(a[201] & b[365])^(a[200] & b[366])^(a[199] & b[367])^(a[198] & b[368])^(a[197] & b[369])^(a[196] & b[370])^(a[195] & b[371])^(a[194] & b[372])^(a[193] & b[373])^(a[192] & b[374])^(a[191] & b[375])^(a[190] & b[376])^(a[189] & b[377])^(a[188] & b[378])^(a[187] & b[379])^(a[186] & b[380])^(a[185] & b[381])^(a[184] & b[382])^(a[183] & b[383])^(a[182] & b[384])^(a[181] & b[385])^(a[180] & b[386])^(a[179] & b[387])^(a[178] & b[388])^(a[177] & b[389])^(a[176] & b[390])^(a[175] & b[391])^(a[174] & b[392])^(a[173] & b[393])^(a[172] & b[394])^(a[171] & b[395])^(a[170] & b[396])^(a[169] & b[397])^(a[168] & b[398])^(a[167] & b[399])^(a[166] & b[400])^(a[165] & b[401])^(a[164] & b[402])^(a[163] & b[403])^(a[162] & b[404])^(a[161] & b[405])^(a[160] & b[406])^(a[159] & b[407])^(a[158] & b[408]);
assign y[567] = (a[408] & b[159])^(a[407] & b[160])^(a[406] & b[161])^(a[405] & b[162])^(a[404] & b[163])^(a[403] & b[164])^(a[402] & b[165])^(a[401] & b[166])^(a[400] & b[167])^(a[399] & b[168])^(a[398] & b[169])^(a[397] & b[170])^(a[396] & b[171])^(a[395] & b[172])^(a[394] & b[173])^(a[393] & b[174])^(a[392] & b[175])^(a[391] & b[176])^(a[390] & b[177])^(a[389] & b[178])^(a[388] & b[179])^(a[387] & b[180])^(a[386] & b[181])^(a[385] & b[182])^(a[384] & b[183])^(a[383] & b[184])^(a[382] & b[185])^(a[381] & b[186])^(a[380] & b[187])^(a[379] & b[188])^(a[378] & b[189])^(a[377] & b[190])^(a[376] & b[191])^(a[375] & b[192])^(a[374] & b[193])^(a[373] & b[194])^(a[372] & b[195])^(a[371] & b[196])^(a[370] & b[197])^(a[369] & b[198])^(a[368] & b[199])^(a[367] & b[200])^(a[366] & b[201])^(a[365] & b[202])^(a[364] & b[203])^(a[363] & b[204])^(a[362] & b[205])^(a[361] & b[206])^(a[360] & b[207])^(a[359] & b[208])^(a[358] & b[209])^(a[357] & b[210])^(a[356] & b[211])^(a[355] & b[212])^(a[354] & b[213])^(a[353] & b[214])^(a[352] & b[215])^(a[351] & b[216])^(a[350] & b[217])^(a[349] & b[218])^(a[348] & b[219])^(a[347] & b[220])^(a[346] & b[221])^(a[345] & b[222])^(a[344] & b[223])^(a[343] & b[224])^(a[342] & b[225])^(a[341] & b[226])^(a[340] & b[227])^(a[339] & b[228])^(a[338] & b[229])^(a[337] & b[230])^(a[336] & b[231])^(a[335] & b[232])^(a[334] & b[233])^(a[333] & b[234])^(a[332] & b[235])^(a[331] & b[236])^(a[330] & b[237])^(a[329] & b[238])^(a[328] & b[239])^(a[327] & b[240])^(a[326] & b[241])^(a[325] & b[242])^(a[324] & b[243])^(a[323] & b[244])^(a[322] & b[245])^(a[321] & b[246])^(a[320] & b[247])^(a[319] & b[248])^(a[318] & b[249])^(a[317] & b[250])^(a[316] & b[251])^(a[315] & b[252])^(a[314] & b[253])^(a[313] & b[254])^(a[312] & b[255])^(a[311] & b[256])^(a[310] & b[257])^(a[309] & b[258])^(a[308] & b[259])^(a[307] & b[260])^(a[306] & b[261])^(a[305] & b[262])^(a[304] & b[263])^(a[303] & b[264])^(a[302] & b[265])^(a[301] & b[266])^(a[300] & b[267])^(a[299] & b[268])^(a[298] & b[269])^(a[297] & b[270])^(a[296] & b[271])^(a[295] & b[272])^(a[294] & b[273])^(a[293] & b[274])^(a[292] & b[275])^(a[291] & b[276])^(a[290] & b[277])^(a[289] & b[278])^(a[288] & b[279])^(a[287] & b[280])^(a[286] & b[281])^(a[285] & b[282])^(a[284] & b[283])^(a[283] & b[284])^(a[282] & b[285])^(a[281] & b[286])^(a[280] & b[287])^(a[279] & b[288])^(a[278] & b[289])^(a[277] & b[290])^(a[276] & b[291])^(a[275] & b[292])^(a[274] & b[293])^(a[273] & b[294])^(a[272] & b[295])^(a[271] & b[296])^(a[270] & b[297])^(a[269] & b[298])^(a[268] & b[299])^(a[267] & b[300])^(a[266] & b[301])^(a[265] & b[302])^(a[264] & b[303])^(a[263] & b[304])^(a[262] & b[305])^(a[261] & b[306])^(a[260] & b[307])^(a[259] & b[308])^(a[258] & b[309])^(a[257] & b[310])^(a[256] & b[311])^(a[255] & b[312])^(a[254] & b[313])^(a[253] & b[314])^(a[252] & b[315])^(a[251] & b[316])^(a[250] & b[317])^(a[249] & b[318])^(a[248] & b[319])^(a[247] & b[320])^(a[246] & b[321])^(a[245] & b[322])^(a[244] & b[323])^(a[243] & b[324])^(a[242] & b[325])^(a[241] & b[326])^(a[240] & b[327])^(a[239] & b[328])^(a[238] & b[329])^(a[237] & b[330])^(a[236] & b[331])^(a[235] & b[332])^(a[234] & b[333])^(a[233] & b[334])^(a[232] & b[335])^(a[231] & b[336])^(a[230] & b[337])^(a[229] & b[338])^(a[228] & b[339])^(a[227] & b[340])^(a[226] & b[341])^(a[225] & b[342])^(a[224] & b[343])^(a[223] & b[344])^(a[222] & b[345])^(a[221] & b[346])^(a[220] & b[347])^(a[219] & b[348])^(a[218] & b[349])^(a[217] & b[350])^(a[216] & b[351])^(a[215] & b[352])^(a[214] & b[353])^(a[213] & b[354])^(a[212] & b[355])^(a[211] & b[356])^(a[210] & b[357])^(a[209] & b[358])^(a[208] & b[359])^(a[207] & b[360])^(a[206] & b[361])^(a[205] & b[362])^(a[204] & b[363])^(a[203] & b[364])^(a[202] & b[365])^(a[201] & b[366])^(a[200] & b[367])^(a[199] & b[368])^(a[198] & b[369])^(a[197] & b[370])^(a[196] & b[371])^(a[195] & b[372])^(a[194] & b[373])^(a[193] & b[374])^(a[192] & b[375])^(a[191] & b[376])^(a[190] & b[377])^(a[189] & b[378])^(a[188] & b[379])^(a[187] & b[380])^(a[186] & b[381])^(a[185] & b[382])^(a[184] & b[383])^(a[183] & b[384])^(a[182] & b[385])^(a[181] & b[386])^(a[180] & b[387])^(a[179] & b[388])^(a[178] & b[389])^(a[177] & b[390])^(a[176] & b[391])^(a[175] & b[392])^(a[174] & b[393])^(a[173] & b[394])^(a[172] & b[395])^(a[171] & b[396])^(a[170] & b[397])^(a[169] & b[398])^(a[168] & b[399])^(a[167] & b[400])^(a[166] & b[401])^(a[165] & b[402])^(a[164] & b[403])^(a[163] & b[404])^(a[162] & b[405])^(a[161] & b[406])^(a[160] & b[407])^(a[159] & b[408]);
assign y[568] = (a[408] & b[160])^(a[407] & b[161])^(a[406] & b[162])^(a[405] & b[163])^(a[404] & b[164])^(a[403] & b[165])^(a[402] & b[166])^(a[401] & b[167])^(a[400] & b[168])^(a[399] & b[169])^(a[398] & b[170])^(a[397] & b[171])^(a[396] & b[172])^(a[395] & b[173])^(a[394] & b[174])^(a[393] & b[175])^(a[392] & b[176])^(a[391] & b[177])^(a[390] & b[178])^(a[389] & b[179])^(a[388] & b[180])^(a[387] & b[181])^(a[386] & b[182])^(a[385] & b[183])^(a[384] & b[184])^(a[383] & b[185])^(a[382] & b[186])^(a[381] & b[187])^(a[380] & b[188])^(a[379] & b[189])^(a[378] & b[190])^(a[377] & b[191])^(a[376] & b[192])^(a[375] & b[193])^(a[374] & b[194])^(a[373] & b[195])^(a[372] & b[196])^(a[371] & b[197])^(a[370] & b[198])^(a[369] & b[199])^(a[368] & b[200])^(a[367] & b[201])^(a[366] & b[202])^(a[365] & b[203])^(a[364] & b[204])^(a[363] & b[205])^(a[362] & b[206])^(a[361] & b[207])^(a[360] & b[208])^(a[359] & b[209])^(a[358] & b[210])^(a[357] & b[211])^(a[356] & b[212])^(a[355] & b[213])^(a[354] & b[214])^(a[353] & b[215])^(a[352] & b[216])^(a[351] & b[217])^(a[350] & b[218])^(a[349] & b[219])^(a[348] & b[220])^(a[347] & b[221])^(a[346] & b[222])^(a[345] & b[223])^(a[344] & b[224])^(a[343] & b[225])^(a[342] & b[226])^(a[341] & b[227])^(a[340] & b[228])^(a[339] & b[229])^(a[338] & b[230])^(a[337] & b[231])^(a[336] & b[232])^(a[335] & b[233])^(a[334] & b[234])^(a[333] & b[235])^(a[332] & b[236])^(a[331] & b[237])^(a[330] & b[238])^(a[329] & b[239])^(a[328] & b[240])^(a[327] & b[241])^(a[326] & b[242])^(a[325] & b[243])^(a[324] & b[244])^(a[323] & b[245])^(a[322] & b[246])^(a[321] & b[247])^(a[320] & b[248])^(a[319] & b[249])^(a[318] & b[250])^(a[317] & b[251])^(a[316] & b[252])^(a[315] & b[253])^(a[314] & b[254])^(a[313] & b[255])^(a[312] & b[256])^(a[311] & b[257])^(a[310] & b[258])^(a[309] & b[259])^(a[308] & b[260])^(a[307] & b[261])^(a[306] & b[262])^(a[305] & b[263])^(a[304] & b[264])^(a[303] & b[265])^(a[302] & b[266])^(a[301] & b[267])^(a[300] & b[268])^(a[299] & b[269])^(a[298] & b[270])^(a[297] & b[271])^(a[296] & b[272])^(a[295] & b[273])^(a[294] & b[274])^(a[293] & b[275])^(a[292] & b[276])^(a[291] & b[277])^(a[290] & b[278])^(a[289] & b[279])^(a[288] & b[280])^(a[287] & b[281])^(a[286] & b[282])^(a[285] & b[283])^(a[284] & b[284])^(a[283] & b[285])^(a[282] & b[286])^(a[281] & b[287])^(a[280] & b[288])^(a[279] & b[289])^(a[278] & b[290])^(a[277] & b[291])^(a[276] & b[292])^(a[275] & b[293])^(a[274] & b[294])^(a[273] & b[295])^(a[272] & b[296])^(a[271] & b[297])^(a[270] & b[298])^(a[269] & b[299])^(a[268] & b[300])^(a[267] & b[301])^(a[266] & b[302])^(a[265] & b[303])^(a[264] & b[304])^(a[263] & b[305])^(a[262] & b[306])^(a[261] & b[307])^(a[260] & b[308])^(a[259] & b[309])^(a[258] & b[310])^(a[257] & b[311])^(a[256] & b[312])^(a[255] & b[313])^(a[254] & b[314])^(a[253] & b[315])^(a[252] & b[316])^(a[251] & b[317])^(a[250] & b[318])^(a[249] & b[319])^(a[248] & b[320])^(a[247] & b[321])^(a[246] & b[322])^(a[245] & b[323])^(a[244] & b[324])^(a[243] & b[325])^(a[242] & b[326])^(a[241] & b[327])^(a[240] & b[328])^(a[239] & b[329])^(a[238] & b[330])^(a[237] & b[331])^(a[236] & b[332])^(a[235] & b[333])^(a[234] & b[334])^(a[233] & b[335])^(a[232] & b[336])^(a[231] & b[337])^(a[230] & b[338])^(a[229] & b[339])^(a[228] & b[340])^(a[227] & b[341])^(a[226] & b[342])^(a[225] & b[343])^(a[224] & b[344])^(a[223] & b[345])^(a[222] & b[346])^(a[221] & b[347])^(a[220] & b[348])^(a[219] & b[349])^(a[218] & b[350])^(a[217] & b[351])^(a[216] & b[352])^(a[215] & b[353])^(a[214] & b[354])^(a[213] & b[355])^(a[212] & b[356])^(a[211] & b[357])^(a[210] & b[358])^(a[209] & b[359])^(a[208] & b[360])^(a[207] & b[361])^(a[206] & b[362])^(a[205] & b[363])^(a[204] & b[364])^(a[203] & b[365])^(a[202] & b[366])^(a[201] & b[367])^(a[200] & b[368])^(a[199] & b[369])^(a[198] & b[370])^(a[197] & b[371])^(a[196] & b[372])^(a[195] & b[373])^(a[194] & b[374])^(a[193] & b[375])^(a[192] & b[376])^(a[191] & b[377])^(a[190] & b[378])^(a[189] & b[379])^(a[188] & b[380])^(a[187] & b[381])^(a[186] & b[382])^(a[185] & b[383])^(a[184] & b[384])^(a[183] & b[385])^(a[182] & b[386])^(a[181] & b[387])^(a[180] & b[388])^(a[179] & b[389])^(a[178] & b[390])^(a[177] & b[391])^(a[176] & b[392])^(a[175] & b[393])^(a[174] & b[394])^(a[173] & b[395])^(a[172] & b[396])^(a[171] & b[397])^(a[170] & b[398])^(a[169] & b[399])^(a[168] & b[400])^(a[167] & b[401])^(a[166] & b[402])^(a[165] & b[403])^(a[164] & b[404])^(a[163] & b[405])^(a[162] & b[406])^(a[161] & b[407])^(a[160] & b[408]);
assign y[569] = (a[408] & b[161])^(a[407] & b[162])^(a[406] & b[163])^(a[405] & b[164])^(a[404] & b[165])^(a[403] & b[166])^(a[402] & b[167])^(a[401] & b[168])^(a[400] & b[169])^(a[399] & b[170])^(a[398] & b[171])^(a[397] & b[172])^(a[396] & b[173])^(a[395] & b[174])^(a[394] & b[175])^(a[393] & b[176])^(a[392] & b[177])^(a[391] & b[178])^(a[390] & b[179])^(a[389] & b[180])^(a[388] & b[181])^(a[387] & b[182])^(a[386] & b[183])^(a[385] & b[184])^(a[384] & b[185])^(a[383] & b[186])^(a[382] & b[187])^(a[381] & b[188])^(a[380] & b[189])^(a[379] & b[190])^(a[378] & b[191])^(a[377] & b[192])^(a[376] & b[193])^(a[375] & b[194])^(a[374] & b[195])^(a[373] & b[196])^(a[372] & b[197])^(a[371] & b[198])^(a[370] & b[199])^(a[369] & b[200])^(a[368] & b[201])^(a[367] & b[202])^(a[366] & b[203])^(a[365] & b[204])^(a[364] & b[205])^(a[363] & b[206])^(a[362] & b[207])^(a[361] & b[208])^(a[360] & b[209])^(a[359] & b[210])^(a[358] & b[211])^(a[357] & b[212])^(a[356] & b[213])^(a[355] & b[214])^(a[354] & b[215])^(a[353] & b[216])^(a[352] & b[217])^(a[351] & b[218])^(a[350] & b[219])^(a[349] & b[220])^(a[348] & b[221])^(a[347] & b[222])^(a[346] & b[223])^(a[345] & b[224])^(a[344] & b[225])^(a[343] & b[226])^(a[342] & b[227])^(a[341] & b[228])^(a[340] & b[229])^(a[339] & b[230])^(a[338] & b[231])^(a[337] & b[232])^(a[336] & b[233])^(a[335] & b[234])^(a[334] & b[235])^(a[333] & b[236])^(a[332] & b[237])^(a[331] & b[238])^(a[330] & b[239])^(a[329] & b[240])^(a[328] & b[241])^(a[327] & b[242])^(a[326] & b[243])^(a[325] & b[244])^(a[324] & b[245])^(a[323] & b[246])^(a[322] & b[247])^(a[321] & b[248])^(a[320] & b[249])^(a[319] & b[250])^(a[318] & b[251])^(a[317] & b[252])^(a[316] & b[253])^(a[315] & b[254])^(a[314] & b[255])^(a[313] & b[256])^(a[312] & b[257])^(a[311] & b[258])^(a[310] & b[259])^(a[309] & b[260])^(a[308] & b[261])^(a[307] & b[262])^(a[306] & b[263])^(a[305] & b[264])^(a[304] & b[265])^(a[303] & b[266])^(a[302] & b[267])^(a[301] & b[268])^(a[300] & b[269])^(a[299] & b[270])^(a[298] & b[271])^(a[297] & b[272])^(a[296] & b[273])^(a[295] & b[274])^(a[294] & b[275])^(a[293] & b[276])^(a[292] & b[277])^(a[291] & b[278])^(a[290] & b[279])^(a[289] & b[280])^(a[288] & b[281])^(a[287] & b[282])^(a[286] & b[283])^(a[285] & b[284])^(a[284] & b[285])^(a[283] & b[286])^(a[282] & b[287])^(a[281] & b[288])^(a[280] & b[289])^(a[279] & b[290])^(a[278] & b[291])^(a[277] & b[292])^(a[276] & b[293])^(a[275] & b[294])^(a[274] & b[295])^(a[273] & b[296])^(a[272] & b[297])^(a[271] & b[298])^(a[270] & b[299])^(a[269] & b[300])^(a[268] & b[301])^(a[267] & b[302])^(a[266] & b[303])^(a[265] & b[304])^(a[264] & b[305])^(a[263] & b[306])^(a[262] & b[307])^(a[261] & b[308])^(a[260] & b[309])^(a[259] & b[310])^(a[258] & b[311])^(a[257] & b[312])^(a[256] & b[313])^(a[255] & b[314])^(a[254] & b[315])^(a[253] & b[316])^(a[252] & b[317])^(a[251] & b[318])^(a[250] & b[319])^(a[249] & b[320])^(a[248] & b[321])^(a[247] & b[322])^(a[246] & b[323])^(a[245] & b[324])^(a[244] & b[325])^(a[243] & b[326])^(a[242] & b[327])^(a[241] & b[328])^(a[240] & b[329])^(a[239] & b[330])^(a[238] & b[331])^(a[237] & b[332])^(a[236] & b[333])^(a[235] & b[334])^(a[234] & b[335])^(a[233] & b[336])^(a[232] & b[337])^(a[231] & b[338])^(a[230] & b[339])^(a[229] & b[340])^(a[228] & b[341])^(a[227] & b[342])^(a[226] & b[343])^(a[225] & b[344])^(a[224] & b[345])^(a[223] & b[346])^(a[222] & b[347])^(a[221] & b[348])^(a[220] & b[349])^(a[219] & b[350])^(a[218] & b[351])^(a[217] & b[352])^(a[216] & b[353])^(a[215] & b[354])^(a[214] & b[355])^(a[213] & b[356])^(a[212] & b[357])^(a[211] & b[358])^(a[210] & b[359])^(a[209] & b[360])^(a[208] & b[361])^(a[207] & b[362])^(a[206] & b[363])^(a[205] & b[364])^(a[204] & b[365])^(a[203] & b[366])^(a[202] & b[367])^(a[201] & b[368])^(a[200] & b[369])^(a[199] & b[370])^(a[198] & b[371])^(a[197] & b[372])^(a[196] & b[373])^(a[195] & b[374])^(a[194] & b[375])^(a[193] & b[376])^(a[192] & b[377])^(a[191] & b[378])^(a[190] & b[379])^(a[189] & b[380])^(a[188] & b[381])^(a[187] & b[382])^(a[186] & b[383])^(a[185] & b[384])^(a[184] & b[385])^(a[183] & b[386])^(a[182] & b[387])^(a[181] & b[388])^(a[180] & b[389])^(a[179] & b[390])^(a[178] & b[391])^(a[177] & b[392])^(a[176] & b[393])^(a[175] & b[394])^(a[174] & b[395])^(a[173] & b[396])^(a[172] & b[397])^(a[171] & b[398])^(a[170] & b[399])^(a[169] & b[400])^(a[168] & b[401])^(a[167] & b[402])^(a[166] & b[403])^(a[165] & b[404])^(a[164] & b[405])^(a[163] & b[406])^(a[162] & b[407])^(a[161] & b[408]);
assign y[570] = (a[408] & b[162])^(a[407] & b[163])^(a[406] & b[164])^(a[405] & b[165])^(a[404] & b[166])^(a[403] & b[167])^(a[402] & b[168])^(a[401] & b[169])^(a[400] & b[170])^(a[399] & b[171])^(a[398] & b[172])^(a[397] & b[173])^(a[396] & b[174])^(a[395] & b[175])^(a[394] & b[176])^(a[393] & b[177])^(a[392] & b[178])^(a[391] & b[179])^(a[390] & b[180])^(a[389] & b[181])^(a[388] & b[182])^(a[387] & b[183])^(a[386] & b[184])^(a[385] & b[185])^(a[384] & b[186])^(a[383] & b[187])^(a[382] & b[188])^(a[381] & b[189])^(a[380] & b[190])^(a[379] & b[191])^(a[378] & b[192])^(a[377] & b[193])^(a[376] & b[194])^(a[375] & b[195])^(a[374] & b[196])^(a[373] & b[197])^(a[372] & b[198])^(a[371] & b[199])^(a[370] & b[200])^(a[369] & b[201])^(a[368] & b[202])^(a[367] & b[203])^(a[366] & b[204])^(a[365] & b[205])^(a[364] & b[206])^(a[363] & b[207])^(a[362] & b[208])^(a[361] & b[209])^(a[360] & b[210])^(a[359] & b[211])^(a[358] & b[212])^(a[357] & b[213])^(a[356] & b[214])^(a[355] & b[215])^(a[354] & b[216])^(a[353] & b[217])^(a[352] & b[218])^(a[351] & b[219])^(a[350] & b[220])^(a[349] & b[221])^(a[348] & b[222])^(a[347] & b[223])^(a[346] & b[224])^(a[345] & b[225])^(a[344] & b[226])^(a[343] & b[227])^(a[342] & b[228])^(a[341] & b[229])^(a[340] & b[230])^(a[339] & b[231])^(a[338] & b[232])^(a[337] & b[233])^(a[336] & b[234])^(a[335] & b[235])^(a[334] & b[236])^(a[333] & b[237])^(a[332] & b[238])^(a[331] & b[239])^(a[330] & b[240])^(a[329] & b[241])^(a[328] & b[242])^(a[327] & b[243])^(a[326] & b[244])^(a[325] & b[245])^(a[324] & b[246])^(a[323] & b[247])^(a[322] & b[248])^(a[321] & b[249])^(a[320] & b[250])^(a[319] & b[251])^(a[318] & b[252])^(a[317] & b[253])^(a[316] & b[254])^(a[315] & b[255])^(a[314] & b[256])^(a[313] & b[257])^(a[312] & b[258])^(a[311] & b[259])^(a[310] & b[260])^(a[309] & b[261])^(a[308] & b[262])^(a[307] & b[263])^(a[306] & b[264])^(a[305] & b[265])^(a[304] & b[266])^(a[303] & b[267])^(a[302] & b[268])^(a[301] & b[269])^(a[300] & b[270])^(a[299] & b[271])^(a[298] & b[272])^(a[297] & b[273])^(a[296] & b[274])^(a[295] & b[275])^(a[294] & b[276])^(a[293] & b[277])^(a[292] & b[278])^(a[291] & b[279])^(a[290] & b[280])^(a[289] & b[281])^(a[288] & b[282])^(a[287] & b[283])^(a[286] & b[284])^(a[285] & b[285])^(a[284] & b[286])^(a[283] & b[287])^(a[282] & b[288])^(a[281] & b[289])^(a[280] & b[290])^(a[279] & b[291])^(a[278] & b[292])^(a[277] & b[293])^(a[276] & b[294])^(a[275] & b[295])^(a[274] & b[296])^(a[273] & b[297])^(a[272] & b[298])^(a[271] & b[299])^(a[270] & b[300])^(a[269] & b[301])^(a[268] & b[302])^(a[267] & b[303])^(a[266] & b[304])^(a[265] & b[305])^(a[264] & b[306])^(a[263] & b[307])^(a[262] & b[308])^(a[261] & b[309])^(a[260] & b[310])^(a[259] & b[311])^(a[258] & b[312])^(a[257] & b[313])^(a[256] & b[314])^(a[255] & b[315])^(a[254] & b[316])^(a[253] & b[317])^(a[252] & b[318])^(a[251] & b[319])^(a[250] & b[320])^(a[249] & b[321])^(a[248] & b[322])^(a[247] & b[323])^(a[246] & b[324])^(a[245] & b[325])^(a[244] & b[326])^(a[243] & b[327])^(a[242] & b[328])^(a[241] & b[329])^(a[240] & b[330])^(a[239] & b[331])^(a[238] & b[332])^(a[237] & b[333])^(a[236] & b[334])^(a[235] & b[335])^(a[234] & b[336])^(a[233] & b[337])^(a[232] & b[338])^(a[231] & b[339])^(a[230] & b[340])^(a[229] & b[341])^(a[228] & b[342])^(a[227] & b[343])^(a[226] & b[344])^(a[225] & b[345])^(a[224] & b[346])^(a[223] & b[347])^(a[222] & b[348])^(a[221] & b[349])^(a[220] & b[350])^(a[219] & b[351])^(a[218] & b[352])^(a[217] & b[353])^(a[216] & b[354])^(a[215] & b[355])^(a[214] & b[356])^(a[213] & b[357])^(a[212] & b[358])^(a[211] & b[359])^(a[210] & b[360])^(a[209] & b[361])^(a[208] & b[362])^(a[207] & b[363])^(a[206] & b[364])^(a[205] & b[365])^(a[204] & b[366])^(a[203] & b[367])^(a[202] & b[368])^(a[201] & b[369])^(a[200] & b[370])^(a[199] & b[371])^(a[198] & b[372])^(a[197] & b[373])^(a[196] & b[374])^(a[195] & b[375])^(a[194] & b[376])^(a[193] & b[377])^(a[192] & b[378])^(a[191] & b[379])^(a[190] & b[380])^(a[189] & b[381])^(a[188] & b[382])^(a[187] & b[383])^(a[186] & b[384])^(a[185] & b[385])^(a[184] & b[386])^(a[183] & b[387])^(a[182] & b[388])^(a[181] & b[389])^(a[180] & b[390])^(a[179] & b[391])^(a[178] & b[392])^(a[177] & b[393])^(a[176] & b[394])^(a[175] & b[395])^(a[174] & b[396])^(a[173] & b[397])^(a[172] & b[398])^(a[171] & b[399])^(a[170] & b[400])^(a[169] & b[401])^(a[168] & b[402])^(a[167] & b[403])^(a[166] & b[404])^(a[165] & b[405])^(a[164] & b[406])^(a[163] & b[407])^(a[162] & b[408]);
assign y[571] = (a[408] & b[163])^(a[407] & b[164])^(a[406] & b[165])^(a[405] & b[166])^(a[404] & b[167])^(a[403] & b[168])^(a[402] & b[169])^(a[401] & b[170])^(a[400] & b[171])^(a[399] & b[172])^(a[398] & b[173])^(a[397] & b[174])^(a[396] & b[175])^(a[395] & b[176])^(a[394] & b[177])^(a[393] & b[178])^(a[392] & b[179])^(a[391] & b[180])^(a[390] & b[181])^(a[389] & b[182])^(a[388] & b[183])^(a[387] & b[184])^(a[386] & b[185])^(a[385] & b[186])^(a[384] & b[187])^(a[383] & b[188])^(a[382] & b[189])^(a[381] & b[190])^(a[380] & b[191])^(a[379] & b[192])^(a[378] & b[193])^(a[377] & b[194])^(a[376] & b[195])^(a[375] & b[196])^(a[374] & b[197])^(a[373] & b[198])^(a[372] & b[199])^(a[371] & b[200])^(a[370] & b[201])^(a[369] & b[202])^(a[368] & b[203])^(a[367] & b[204])^(a[366] & b[205])^(a[365] & b[206])^(a[364] & b[207])^(a[363] & b[208])^(a[362] & b[209])^(a[361] & b[210])^(a[360] & b[211])^(a[359] & b[212])^(a[358] & b[213])^(a[357] & b[214])^(a[356] & b[215])^(a[355] & b[216])^(a[354] & b[217])^(a[353] & b[218])^(a[352] & b[219])^(a[351] & b[220])^(a[350] & b[221])^(a[349] & b[222])^(a[348] & b[223])^(a[347] & b[224])^(a[346] & b[225])^(a[345] & b[226])^(a[344] & b[227])^(a[343] & b[228])^(a[342] & b[229])^(a[341] & b[230])^(a[340] & b[231])^(a[339] & b[232])^(a[338] & b[233])^(a[337] & b[234])^(a[336] & b[235])^(a[335] & b[236])^(a[334] & b[237])^(a[333] & b[238])^(a[332] & b[239])^(a[331] & b[240])^(a[330] & b[241])^(a[329] & b[242])^(a[328] & b[243])^(a[327] & b[244])^(a[326] & b[245])^(a[325] & b[246])^(a[324] & b[247])^(a[323] & b[248])^(a[322] & b[249])^(a[321] & b[250])^(a[320] & b[251])^(a[319] & b[252])^(a[318] & b[253])^(a[317] & b[254])^(a[316] & b[255])^(a[315] & b[256])^(a[314] & b[257])^(a[313] & b[258])^(a[312] & b[259])^(a[311] & b[260])^(a[310] & b[261])^(a[309] & b[262])^(a[308] & b[263])^(a[307] & b[264])^(a[306] & b[265])^(a[305] & b[266])^(a[304] & b[267])^(a[303] & b[268])^(a[302] & b[269])^(a[301] & b[270])^(a[300] & b[271])^(a[299] & b[272])^(a[298] & b[273])^(a[297] & b[274])^(a[296] & b[275])^(a[295] & b[276])^(a[294] & b[277])^(a[293] & b[278])^(a[292] & b[279])^(a[291] & b[280])^(a[290] & b[281])^(a[289] & b[282])^(a[288] & b[283])^(a[287] & b[284])^(a[286] & b[285])^(a[285] & b[286])^(a[284] & b[287])^(a[283] & b[288])^(a[282] & b[289])^(a[281] & b[290])^(a[280] & b[291])^(a[279] & b[292])^(a[278] & b[293])^(a[277] & b[294])^(a[276] & b[295])^(a[275] & b[296])^(a[274] & b[297])^(a[273] & b[298])^(a[272] & b[299])^(a[271] & b[300])^(a[270] & b[301])^(a[269] & b[302])^(a[268] & b[303])^(a[267] & b[304])^(a[266] & b[305])^(a[265] & b[306])^(a[264] & b[307])^(a[263] & b[308])^(a[262] & b[309])^(a[261] & b[310])^(a[260] & b[311])^(a[259] & b[312])^(a[258] & b[313])^(a[257] & b[314])^(a[256] & b[315])^(a[255] & b[316])^(a[254] & b[317])^(a[253] & b[318])^(a[252] & b[319])^(a[251] & b[320])^(a[250] & b[321])^(a[249] & b[322])^(a[248] & b[323])^(a[247] & b[324])^(a[246] & b[325])^(a[245] & b[326])^(a[244] & b[327])^(a[243] & b[328])^(a[242] & b[329])^(a[241] & b[330])^(a[240] & b[331])^(a[239] & b[332])^(a[238] & b[333])^(a[237] & b[334])^(a[236] & b[335])^(a[235] & b[336])^(a[234] & b[337])^(a[233] & b[338])^(a[232] & b[339])^(a[231] & b[340])^(a[230] & b[341])^(a[229] & b[342])^(a[228] & b[343])^(a[227] & b[344])^(a[226] & b[345])^(a[225] & b[346])^(a[224] & b[347])^(a[223] & b[348])^(a[222] & b[349])^(a[221] & b[350])^(a[220] & b[351])^(a[219] & b[352])^(a[218] & b[353])^(a[217] & b[354])^(a[216] & b[355])^(a[215] & b[356])^(a[214] & b[357])^(a[213] & b[358])^(a[212] & b[359])^(a[211] & b[360])^(a[210] & b[361])^(a[209] & b[362])^(a[208] & b[363])^(a[207] & b[364])^(a[206] & b[365])^(a[205] & b[366])^(a[204] & b[367])^(a[203] & b[368])^(a[202] & b[369])^(a[201] & b[370])^(a[200] & b[371])^(a[199] & b[372])^(a[198] & b[373])^(a[197] & b[374])^(a[196] & b[375])^(a[195] & b[376])^(a[194] & b[377])^(a[193] & b[378])^(a[192] & b[379])^(a[191] & b[380])^(a[190] & b[381])^(a[189] & b[382])^(a[188] & b[383])^(a[187] & b[384])^(a[186] & b[385])^(a[185] & b[386])^(a[184] & b[387])^(a[183] & b[388])^(a[182] & b[389])^(a[181] & b[390])^(a[180] & b[391])^(a[179] & b[392])^(a[178] & b[393])^(a[177] & b[394])^(a[176] & b[395])^(a[175] & b[396])^(a[174] & b[397])^(a[173] & b[398])^(a[172] & b[399])^(a[171] & b[400])^(a[170] & b[401])^(a[169] & b[402])^(a[168] & b[403])^(a[167] & b[404])^(a[166] & b[405])^(a[165] & b[406])^(a[164] & b[407])^(a[163] & b[408]);
assign y[572] = (a[408] & b[164])^(a[407] & b[165])^(a[406] & b[166])^(a[405] & b[167])^(a[404] & b[168])^(a[403] & b[169])^(a[402] & b[170])^(a[401] & b[171])^(a[400] & b[172])^(a[399] & b[173])^(a[398] & b[174])^(a[397] & b[175])^(a[396] & b[176])^(a[395] & b[177])^(a[394] & b[178])^(a[393] & b[179])^(a[392] & b[180])^(a[391] & b[181])^(a[390] & b[182])^(a[389] & b[183])^(a[388] & b[184])^(a[387] & b[185])^(a[386] & b[186])^(a[385] & b[187])^(a[384] & b[188])^(a[383] & b[189])^(a[382] & b[190])^(a[381] & b[191])^(a[380] & b[192])^(a[379] & b[193])^(a[378] & b[194])^(a[377] & b[195])^(a[376] & b[196])^(a[375] & b[197])^(a[374] & b[198])^(a[373] & b[199])^(a[372] & b[200])^(a[371] & b[201])^(a[370] & b[202])^(a[369] & b[203])^(a[368] & b[204])^(a[367] & b[205])^(a[366] & b[206])^(a[365] & b[207])^(a[364] & b[208])^(a[363] & b[209])^(a[362] & b[210])^(a[361] & b[211])^(a[360] & b[212])^(a[359] & b[213])^(a[358] & b[214])^(a[357] & b[215])^(a[356] & b[216])^(a[355] & b[217])^(a[354] & b[218])^(a[353] & b[219])^(a[352] & b[220])^(a[351] & b[221])^(a[350] & b[222])^(a[349] & b[223])^(a[348] & b[224])^(a[347] & b[225])^(a[346] & b[226])^(a[345] & b[227])^(a[344] & b[228])^(a[343] & b[229])^(a[342] & b[230])^(a[341] & b[231])^(a[340] & b[232])^(a[339] & b[233])^(a[338] & b[234])^(a[337] & b[235])^(a[336] & b[236])^(a[335] & b[237])^(a[334] & b[238])^(a[333] & b[239])^(a[332] & b[240])^(a[331] & b[241])^(a[330] & b[242])^(a[329] & b[243])^(a[328] & b[244])^(a[327] & b[245])^(a[326] & b[246])^(a[325] & b[247])^(a[324] & b[248])^(a[323] & b[249])^(a[322] & b[250])^(a[321] & b[251])^(a[320] & b[252])^(a[319] & b[253])^(a[318] & b[254])^(a[317] & b[255])^(a[316] & b[256])^(a[315] & b[257])^(a[314] & b[258])^(a[313] & b[259])^(a[312] & b[260])^(a[311] & b[261])^(a[310] & b[262])^(a[309] & b[263])^(a[308] & b[264])^(a[307] & b[265])^(a[306] & b[266])^(a[305] & b[267])^(a[304] & b[268])^(a[303] & b[269])^(a[302] & b[270])^(a[301] & b[271])^(a[300] & b[272])^(a[299] & b[273])^(a[298] & b[274])^(a[297] & b[275])^(a[296] & b[276])^(a[295] & b[277])^(a[294] & b[278])^(a[293] & b[279])^(a[292] & b[280])^(a[291] & b[281])^(a[290] & b[282])^(a[289] & b[283])^(a[288] & b[284])^(a[287] & b[285])^(a[286] & b[286])^(a[285] & b[287])^(a[284] & b[288])^(a[283] & b[289])^(a[282] & b[290])^(a[281] & b[291])^(a[280] & b[292])^(a[279] & b[293])^(a[278] & b[294])^(a[277] & b[295])^(a[276] & b[296])^(a[275] & b[297])^(a[274] & b[298])^(a[273] & b[299])^(a[272] & b[300])^(a[271] & b[301])^(a[270] & b[302])^(a[269] & b[303])^(a[268] & b[304])^(a[267] & b[305])^(a[266] & b[306])^(a[265] & b[307])^(a[264] & b[308])^(a[263] & b[309])^(a[262] & b[310])^(a[261] & b[311])^(a[260] & b[312])^(a[259] & b[313])^(a[258] & b[314])^(a[257] & b[315])^(a[256] & b[316])^(a[255] & b[317])^(a[254] & b[318])^(a[253] & b[319])^(a[252] & b[320])^(a[251] & b[321])^(a[250] & b[322])^(a[249] & b[323])^(a[248] & b[324])^(a[247] & b[325])^(a[246] & b[326])^(a[245] & b[327])^(a[244] & b[328])^(a[243] & b[329])^(a[242] & b[330])^(a[241] & b[331])^(a[240] & b[332])^(a[239] & b[333])^(a[238] & b[334])^(a[237] & b[335])^(a[236] & b[336])^(a[235] & b[337])^(a[234] & b[338])^(a[233] & b[339])^(a[232] & b[340])^(a[231] & b[341])^(a[230] & b[342])^(a[229] & b[343])^(a[228] & b[344])^(a[227] & b[345])^(a[226] & b[346])^(a[225] & b[347])^(a[224] & b[348])^(a[223] & b[349])^(a[222] & b[350])^(a[221] & b[351])^(a[220] & b[352])^(a[219] & b[353])^(a[218] & b[354])^(a[217] & b[355])^(a[216] & b[356])^(a[215] & b[357])^(a[214] & b[358])^(a[213] & b[359])^(a[212] & b[360])^(a[211] & b[361])^(a[210] & b[362])^(a[209] & b[363])^(a[208] & b[364])^(a[207] & b[365])^(a[206] & b[366])^(a[205] & b[367])^(a[204] & b[368])^(a[203] & b[369])^(a[202] & b[370])^(a[201] & b[371])^(a[200] & b[372])^(a[199] & b[373])^(a[198] & b[374])^(a[197] & b[375])^(a[196] & b[376])^(a[195] & b[377])^(a[194] & b[378])^(a[193] & b[379])^(a[192] & b[380])^(a[191] & b[381])^(a[190] & b[382])^(a[189] & b[383])^(a[188] & b[384])^(a[187] & b[385])^(a[186] & b[386])^(a[185] & b[387])^(a[184] & b[388])^(a[183] & b[389])^(a[182] & b[390])^(a[181] & b[391])^(a[180] & b[392])^(a[179] & b[393])^(a[178] & b[394])^(a[177] & b[395])^(a[176] & b[396])^(a[175] & b[397])^(a[174] & b[398])^(a[173] & b[399])^(a[172] & b[400])^(a[171] & b[401])^(a[170] & b[402])^(a[169] & b[403])^(a[168] & b[404])^(a[167] & b[405])^(a[166] & b[406])^(a[165] & b[407])^(a[164] & b[408]);
assign y[573] = (a[408] & b[165])^(a[407] & b[166])^(a[406] & b[167])^(a[405] & b[168])^(a[404] & b[169])^(a[403] & b[170])^(a[402] & b[171])^(a[401] & b[172])^(a[400] & b[173])^(a[399] & b[174])^(a[398] & b[175])^(a[397] & b[176])^(a[396] & b[177])^(a[395] & b[178])^(a[394] & b[179])^(a[393] & b[180])^(a[392] & b[181])^(a[391] & b[182])^(a[390] & b[183])^(a[389] & b[184])^(a[388] & b[185])^(a[387] & b[186])^(a[386] & b[187])^(a[385] & b[188])^(a[384] & b[189])^(a[383] & b[190])^(a[382] & b[191])^(a[381] & b[192])^(a[380] & b[193])^(a[379] & b[194])^(a[378] & b[195])^(a[377] & b[196])^(a[376] & b[197])^(a[375] & b[198])^(a[374] & b[199])^(a[373] & b[200])^(a[372] & b[201])^(a[371] & b[202])^(a[370] & b[203])^(a[369] & b[204])^(a[368] & b[205])^(a[367] & b[206])^(a[366] & b[207])^(a[365] & b[208])^(a[364] & b[209])^(a[363] & b[210])^(a[362] & b[211])^(a[361] & b[212])^(a[360] & b[213])^(a[359] & b[214])^(a[358] & b[215])^(a[357] & b[216])^(a[356] & b[217])^(a[355] & b[218])^(a[354] & b[219])^(a[353] & b[220])^(a[352] & b[221])^(a[351] & b[222])^(a[350] & b[223])^(a[349] & b[224])^(a[348] & b[225])^(a[347] & b[226])^(a[346] & b[227])^(a[345] & b[228])^(a[344] & b[229])^(a[343] & b[230])^(a[342] & b[231])^(a[341] & b[232])^(a[340] & b[233])^(a[339] & b[234])^(a[338] & b[235])^(a[337] & b[236])^(a[336] & b[237])^(a[335] & b[238])^(a[334] & b[239])^(a[333] & b[240])^(a[332] & b[241])^(a[331] & b[242])^(a[330] & b[243])^(a[329] & b[244])^(a[328] & b[245])^(a[327] & b[246])^(a[326] & b[247])^(a[325] & b[248])^(a[324] & b[249])^(a[323] & b[250])^(a[322] & b[251])^(a[321] & b[252])^(a[320] & b[253])^(a[319] & b[254])^(a[318] & b[255])^(a[317] & b[256])^(a[316] & b[257])^(a[315] & b[258])^(a[314] & b[259])^(a[313] & b[260])^(a[312] & b[261])^(a[311] & b[262])^(a[310] & b[263])^(a[309] & b[264])^(a[308] & b[265])^(a[307] & b[266])^(a[306] & b[267])^(a[305] & b[268])^(a[304] & b[269])^(a[303] & b[270])^(a[302] & b[271])^(a[301] & b[272])^(a[300] & b[273])^(a[299] & b[274])^(a[298] & b[275])^(a[297] & b[276])^(a[296] & b[277])^(a[295] & b[278])^(a[294] & b[279])^(a[293] & b[280])^(a[292] & b[281])^(a[291] & b[282])^(a[290] & b[283])^(a[289] & b[284])^(a[288] & b[285])^(a[287] & b[286])^(a[286] & b[287])^(a[285] & b[288])^(a[284] & b[289])^(a[283] & b[290])^(a[282] & b[291])^(a[281] & b[292])^(a[280] & b[293])^(a[279] & b[294])^(a[278] & b[295])^(a[277] & b[296])^(a[276] & b[297])^(a[275] & b[298])^(a[274] & b[299])^(a[273] & b[300])^(a[272] & b[301])^(a[271] & b[302])^(a[270] & b[303])^(a[269] & b[304])^(a[268] & b[305])^(a[267] & b[306])^(a[266] & b[307])^(a[265] & b[308])^(a[264] & b[309])^(a[263] & b[310])^(a[262] & b[311])^(a[261] & b[312])^(a[260] & b[313])^(a[259] & b[314])^(a[258] & b[315])^(a[257] & b[316])^(a[256] & b[317])^(a[255] & b[318])^(a[254] & b[319])^(a[253] & b[320])^(a[252] & b[321])^(a[251] & b[322])^(a[250] & b[323])^(a[249] & b[324])^(a[248] & b[325])^(a[247] & b[326])^(a[246] & b[327])^(a[245] & b[328])^(a[244] & b[329])^(a[243] & b[330])^(a[242] & b[331])^(a[241] & b[332])^(a[240] & b[333])^(a[239] & b[334])^(a[238] & b[335])^(a[237] & b[336])^(a[236] & b[337])^(a[235] & b[338])^(a[234] & b[339])^(a[233] & b[340])^(a[232] & b[341])^(a[231] & b[342])^(a[230] & b[343])^(a[229] & b[344])^(a[228] & b[345])^(a[227] & b[346])^(a[226] & b[347])^(a[225] & b[348])^(a[224] & b[349])^(a[223] & b[350])^(a[222] & b[351])^(a[221] & b[352])^(a[220] & b[353])^(a[219] & b[354])^(a[218] & b[355])^(a[217] & b[356])^(a[216] & b[357])^(a[215] & b[358])^(a[214] & b[359])^(a[213] & b[360])^(a[212] & b[361])^(a[211] & b[362])^(a[210] & b[363])^(a[209] & b[364])^(a[208] & b[365])^(a[207] & b[366])^(a[206] & b[367])^(a[205] & b[368])^(a[204] & b[369])^(a[203] & b[370])^(a[202] & b[371])^(a[201] & b[372])^(a[200] & b[373])^(a[199] & b[374])^(a[198] & b[375])^(a[197] & b[376])^(a[196] & b[377])^(a[195] & b[378])^(a[194] & b[379])^(a[193] & b[380])^(a[192] & b[381])^(a[191] & b[382])^(a[190] & b[383])^(a[189] & b[384])^(a[188] & b[385])^(a[187] & b[386])^(a[186] & b[387])^(a[185] & b[388])^(a[184] & b[389])^(a[183] & b[390])^(a[182] & b[391])^(a[181] & b[392])^(a[180] & b[393])^(a[179] & b[394])^(a[178] & b[395])^(a[177] & b[396])^(a[176] & b[397])^(a[175] & b[398])^(a[174] & b[399])^(a[173] & b[400])^(a[172] & b[401])^(a[171] & b[402])^(a[170] & b[403])^(a[169] & b[404])^(a[168] & b[405])^(a[167] & b[406])^(a[166] & b[407])^(a[165] & b[408]);
assign y[574] = (a[408] & b[166])^(a[407] & b[167])^(a[406] & b[168])^(a[405] & b[169])^(a[404] & b[170])^(a[403] & b[171])^(a[402] & b[172])^(a[401] & b[173])^(a[400] & b[174])^(a[399] & b[175])^(a[398] & b[176])^(a[397] & b[177])^(a[396] & b[178])^(a[395] & b[179])^(a[394] & b[180])^(a[393] & b[181])^(a[392] & b[182])^(a[391] & b[183])^(a[390] & b[184])^(a[389] & b[185])^(a[388] & b[186])^(a[387] & b[187])^(a[386] & b[188])^(a[385] & b[189])^(a[384] & b[190])^(a[383] & b[191])^(a[382] & b[192])^(a[381] & b[193])^(a[380] & b[194])^(a[379] & b[195])^(a[378] & b[196])^(a[377] & b[197])^(a[376] & b[198])^(a[375] & b[199])^(a[374] & b[200])^(a[373] & b[201])^(a[372] & b[202])^(a[371] & b[203])^(a[370] & b[204])^(a[369] & b[205])^(a[368] & b[206])^(a[367] & b[207])^(a[366] & b[208])^(a[365] & b[209])^(a[364] & b[210])^(a[363] & b[211])^(a[362] & b[212])^(a[361] & b[213])^(a[360] & b[214])^(a[359] & b[215])^(a[358] & b[216])^(a[357] & b[217])^(a[356] & b[218])^(a[355] & b[219])^(a[354] & b[220])^(a[353] & b[221])^(a[352] & b[222])^(a[351] & b[223])^(a[350] & b[224])^(a[349] & b[225])^(a[348] & b[226])^(a[347] & b[227])^(a[346] & b[228])^(a[345] & b[229])^(a[344] & b[230])^(a[343] & b[231])^(a[342] & b[232])^(a[341] & b[233])^(a[340] & b[234])^(a[339] & b[235])^(a[338] & b[236])^(a[337] & b[237])^(a[336] & b[238])^(a[335] & b[239])^(a[334] & b[240])^(a[333] & b[241])^(a[332] & b[242])^(a[331] & b[243])^(a[330] & b[244])^(a[329] & b[245])^(a[328] & b[246])^(a[327] & b[247])^(a[326] & b[248])^(a[325] & b[249])^(a[324] & b[250])^(a[323] & b[251])^(a[322] & b[252])^(a[321] & b[253])^(a[320] & b[254])^(a[319] & b[255])^(a[318] & b[256])^(a[317] & b[257])^(a[316] & b[258])^(a[315] & b[259])^(a[314] & b[260])^(a[313] & b[261])^(a[312] & b[262])^(a[311] & b[263])^(a[310] & b[264])^(a[309] & b[265])^(a[308] & b[266])^(a[307] & b[267])^(a[306] & b[268])^(a[305] & b[269])^(a[304] & b[270])^(a[303] & b[271])^(a[302] & b[272])^(a[301] & b[273])^(a[300] & b[274])^(a[299] & b[275])^(a[298] & b[276])^(a[297] & b[277])^(a[296] & b[278])^(a[295] & b[279])^(a[294] & b[280])^(a[293] & b[281])^(a[292] & b[282])^(a[291] & b[283])^(a[290] & b[284])^(a[289] & b[285])^(a[288] & b[286])^(a[287] & b[287])^(a[286] & b[288])^(a[285] & b[289])^(a[284] & b[290])^(a[283] & b[291])^(a[282] & b[292])^(a[281] & b[293])^(a[280] & b[294])^(a[279] & b[295])^(a[278] & b[296])^(a[277] & b[297])^(a[276] & b[298])^(a[275] & b[299])^(a[274] & b[300])^(a[273] & b[301])^(a[272] & b[302])^(a[271] & b[303])^(a[270] & b[304])^(a[269] & b[305])^(a[268] & b[306])^(a[267] & b[307])^(a[266] & b[308])^(a[265] & b[309])^(a[264] & b[310])^(a[263] & b[311])^(a[262] & b[312])^(a[261] & b[313])^(a[260] & b[314])^(a[259] & b[315])^(a[258] & b[316])^(a[257] & b[317])^(a[256] & b[318])^(a[255] & b[319])^(a[254] & b[320])^(a[253] & b[321])^(a[252] & b[322])^(a[251] & b[323])^(a[250] & b[324])^(a[249] & b[325])^(a[248] & b[326])^(a[247] & b[327])^(a[246] & b[328])^(a[245] & b[329])^(a[244] & b[330])^(a[243] & b[331])^(a[242] & b[332])^(a[241] & b[333])^(a[240] & b[334])^(a[239] & b[335])^(a[238] & b[336])^(a[237] & b[337])^(a[236] & b[338])^(a[235] & b[339])^(a[234] & b[340])^(a[233] & b[341])^(a[232] & b[342])^(a[231] & b[343])^(a[230] & b[344])^(a[229] & b[345])^(a[228] & b[346])^(a[227] & b[347])^(a[226] & b[348])^(a[225] & b[349])^(a[224] & b[350])^(a[223] & b[351])^(a[222] & b[352])^(a[221] & b[353])^(a[220] & b[354])^(a[219] & b[355])^(a[218] & b[356])^(a[217] & b[357])^(a[216] & b[358])^(a[215] & b[359])^(a[214] & b[360])^(a[213] & b[361])^(a[212] & b[362])^(a[211] & b[363])^(a[210] & b[364])^(a[209] & b[365])^(a[208] & b[366])^(a[207] & b[367])^(a[206] & b[368])^(a[205] & b[369])^(a[204] & b[370])^(a[203] & b[371])^(a[202] & b[372])^(a[201] & b[373])^(a[200] & b[374])^(a[199] & b[375])^(a[198] & b[376])^(a[197] & b[377])^(a[196] & b[378])^(a[195] & b[379])^(a[194] & b[380])^(a[193] & b[381])^(a[192] & b[382])^(a[191] & b[383])^(a[190] & b[384])^(a[189] & b[385])^(a[188] & b[386])^(a[187] & b[387])^(a[186] & b[388])^(a[185] & b[389])^(a[184] & b[390])^(a[183] & b[391])^(a[182] & b[392])^(a[181] & b[393])^(a[180] & b[394])^(a[179] & b[395])^(a[178] & b[396])^(a[177] & b[397])^(a[176] & b[398])^(a[175] & b[399])^(a[174] & b[400])^(a[173] & b[401])^(a[172] & b[402])^(a[171] & b[403])^(a[170] & b[404])^(a[169] & b[405])^(a[168] & b[406])^(a[167] & b[407])^(a[166] & b[408]);
assign y[575] = (a[408] & b[167])^(a[407] & b[168])^(a[406] & b[169])^(a[405] & b[170])^(a[404] & b[171])^(a[403] & b[172])^(a[402] & b[173])^(a[401] & b[174])^(a[400] & b[175])^(a[399] & b[176])^(a[398] & b[177])^(a[397] & b[178])^(a[396] & b[179])^(a[395] & b[180])^(a[394] & b[181])^(a[393] & b[182])^(a[392] & b[183])^(a[391] & b[184])^(a[390] & b[185])^(a[389] & b[186])^(a[388] & b[187])^(a[387] & b[188])^(a[386] & b[189])^(a[385] & b[190])^(a[384] & b[191])^(a[383] & b[192])^(a[382] & b[193])^(a[381] & b[194])^(a[380] & b[195])^(a[379] & b[196])^(a[378] & b[197])^(a[377] & b[198])^(a[376] & b[199])^(a[375] & b[200])^(a[374] & b[201])^(a[373] & b[202])^(a[372] & b[203])^(a[371] & b[204])^(a[370] & b[205])^(a[369] & b[206])^(a[368] & b[207])^(a[367] & b[208])^(a[366] & b[209])^(a[365] & b[210])^(a[364] & b[211])^(a[363] & b[212])^(a[362] & b[213])^(a[361] & b[214])^(a[360] & b[215])^(a[359] & b[216])^(a[358] & b[217])^(a[357] & b[218])^(a[356] & b[219])^(a[355] & b[220])^(a[354] & b[221])^(a[353] & b[222])^(a[352] & b[223])^(a[351] & b[224])^(a[350] & b[225])^(a[349] & b[226])^(a[348] & b[227])^(a[347] & b[228])^(a[346] & b[229])^(a[345] & b[230])^(a[344] & b[231])^(a[343] & b[232])^(a[342] & b[233])^(a[341] & b[234])^(a[340] & b[235])^(a[339] & b[236])^(a[338] & b[237])^(a[337] & b[238])^(a[336] & b[239])^(a[335] & b[240])^(a[334] & b[241])^(a[333] & b[242])^(a[332] & b[243])^(a[331] & b[244])^(a[330] & b[245])^(a[329] & b[246])^(a[328] & b[247])^(a[327] & b[248])^(a[326] & b[249])^(a[325] & b[250])^(a[324] & b[251])^(a[323] & b[252])^(a[322] & b[253])^(a[321] & b[254])^(a[320] & b[255])^(a[319] & b[256])^(a[318] & b[257])^(a[317] & b[258])^(a[316] & b[259])^(a[315] & b[260])^(a[314] & b[261])^(a[313] & b[262])^(a[312] & b[263])^(a[311] & b[264])^(a[310] & b[265])^(a[309] & b[266])^(a[308] & b[267])^(a[307] & b[268])^(a[306] & b[269])^(a[305] & b[270])^(a[304] & b[271])^(a[303] & b[272])^(a[302] & b[273])^(a[301] & b[274])^(a[300] & b[275])^(a[299] & b[276])^(a[298] & b[277])^(a[297] & b[278])^(a[296] & b[279])^(a[295] & b[280])^(a[294] & b[281])^(a[293] & b[282])^(a[292] & b[283])^(a[291] & b[284])^(a[290] & b[285])^(a[289] & b[286])^(a[288] & b[287])^(a[287] & b[288])^(a[286] & b[289])^(a[285] & b[290])^(a[284] & b[291])^(a[283] & b[292])^(a[282] & b[293])^(a[281] & b[294])^(a[280] & b[295])^(a[279] & b[296])^(a[278] & b[297])^(a[277] & b[298])^(a[276] & b[299])^(a[275] & b[300])^(a[274] & b[301])^(a[273] & b[302])^(a[272] & b[303])^(a[271] & b[304])^(a[270] & b[305])^(a[269] & b[306])^(a[268] & b[307])^(a[267] & b[308])^(a[266] & b[309])^(a[265] & b[310])^(a[264] & b[311])^(a[263] & b[312])^(a[262] & b[313])^(a[261] & b[314])^(a[260] & b[315])^(a[259] & b[316])^(a[258] & b[317])^(a[257] & b[318])^(a[256] & b[319])^(a[255] & b[320])^(a[254] & b[321])^(a[253] & b[322])^(a[252] & b[323])^(a[251] & b[324])^(a[250] & b[325])^(a[249] & b[326])^(a[248] & b[327])^(a[247] & b[328])^(a[246] & b[329])^(a[245] & b[330])^(a[244] & b[331])^(a[243] & b[332])^(a[242] & b[333])^(a[241] & b[334])^(a[240] & b[335])^(a[239] & b[336])^(a[238] & b[337])^(a[237] & b[338])^(a[236] & b[339])^(a[235] & b[340])^(a[234] & b[341])^(a[233] & b[342])^(a[232] & b[343])^(a[231] & b[344])^(a[230] & b[345])^(a[229] & b[346])^(a[228] & b[347])^(a[227] & b[348])^(a[226] & b[349])^(a[225] & b[350])^(a[224] & b[351])^(a[223] & b[352])^(a[222] & b[353])^(a[221] & b[354])^(a[220] & b[355])^(a[219] & b[356])^(a[218] & b[357])^(a[217] & b[358])^(a[216] & b[359])^(a[215] & b[360])^(a[214] & b[361])^(a[213] & b[362])^(a[212] & b[363])^(a[211] & b[364])^(a[210] & b[365])^(a[209] & b[366])^(a[208] & b[367])^(a[207] & b[368])^(a[206] & b[369])^(a[205] & b[370])^(a[204] & b[371])^(a[203] & b[372])^(a[202] & b[373])^(a[201] & b[374])^(a[200] & b[375])^(a[199] & b[376])^(a[198] & b[377])^(a[197] & b[378])^(a[196] & b[379])^(a[195] & b[380])^(a[194] & b[381])^(a[193] & b[382])^(a[192] & b[383])^(a[191] & b[384])^(a[190] & b[385])^(a[189] & b[386])^(a[188] & b[387])^(a[187] & b[388])^(a[186] & b[389])^(a[185] & b[390])^(a[184] & b[391])^(a[183] & b[392])^(a[182] & b[393])^(a[181] & b[394])^(a[180] & b[395])^(a[179] & b[396])^(a[178] & b[397])^(a[177] & b[398])^(a[176] & b[399])^(a[175] & b[400])^(a[174] & b[401])^(a[173] & b[402])^(a[172] & b[403])^(a[171] & b[404])^(a[170] & b[405])^(a[169] & b[406])^(a[168] & b[407])^(a[167] & b[408]);
assign y[576] = (a[408] & b[168])^(a[407] & b[169])^(a[406] & b[170])^(a[405] & b[171])^(a[404] & b[172])^(a[403] & b[173])^(a[402] & b[174])^(a[401] & b[175])^(a[400] & b[176])^(a[399] & b[177])^(a[398] & b[178])^(a[397] & b[179])^(a[396] & b[180])^(a[395] & b[181])^(a[394] & b[182])^(a[393] & b[183])^(a[392] & b[184])^(a[391] & b[185])^(a[390] & b[186])^(a[389] & b[187])^(a[388] & b[188])^(a[387] & b[189])^(a[386] & b[190])^(a[385] & b[191])^(a[384] & b[192])^(a[383] & b[193])^(a[382] & b[194])^(a[381] & b[195])^(a[380] & b[196])^(a[379] & b[197])^(a[378] & b[198])^(a[377] & b[199])^(a[376] & b[200])^(a[375] & b[201])^(a[374] & b[202])^(a[373] & b[203])^(a[372] & b[204])^(a[371] & b[205])^(a[370] & b[206])^(a[369] & b[207])^(a[368] & b[208])^(a[367] & b[209])^(a[366] & b[210])^(a[365] & b[211])^(a[364] & b[212])^(a[363] & b[213])^(a[362] & b[214])^(a[361] & b[215])^(a[360] & b[216])^(a[359] & b[217])^(a[358] & b[218])^(a[357] & b[219])^(a[356] & b[220])^(a[355] & b[221])^(a[354] & b[222])^(a[353] & b[223])^(a[352] & b[224])^(a[351] & b[225])^(a[350] & b[226])^(a[349] & b[227])^(a[348] & b[228])^(a[347] & b[229])^(a[346] & b[230])^(a[345] & b[231])^(a[344] & b[232])^(a[343] & b[233])^(a[342] & b[234])^(a[341] & b[235])^(a[340] & b[236])^(a[339] & b[237])^(a[338] & b[238])^(a[337] & b[239])^(a[336] & b[240])^(a[335] & b[241])^(a[334] & b[242])^(a[333] & b[243])^(a[332] & b[244])^(a[331] & b[245])^(a[330] & b[246])^(a[329] & b[247])^(a[328] & b[248])^(a[327] & b[249])^(a[326] & b[250])^(a[325] & b[251])^(a[324] & b[252])^(a[323] & b[253])^(a[322] & b[254])^(a[321] & b[255])^(a[320] & b[256])^(a[319] & b[257])^(a[318] & b[258])^(a[317] & b[259])^(a[316] & b[260])^(a[315] & b[261])^(a[314] & b[262])^(a[313] & b[263])^(a[312] & b[264])^(a[311] & b[265])^(a[310] & b[266])^(a[309] & b[267])^(a[308] & b[268])^(a[307] & b[269])^(a[306] & b[270])^(a[305] & b[271])^(a[304] & b[272])^(a[303] & b[273])^(a[302] & b[274])^(a[301] & b[275])^(a[300] & b[276])^(a[299] & b[277])^(a[298] & b[278])^(a[297] & b[279])^(a[296] & b[280])^(a[295] & b[281])^(a[294] & b[282])^(a[293] & b[283])^(a[292] & b[284])^(a[291] & b[285])^(a[290] & b[286])^(a[289] & b[287])^(a[288] & b[288])^(a[287] & b[289])^(a[286] & b[290])^(a[285] & b[291])^(a[284] & b[292])^(a[283] & b[293])^(a[282] & b[294])^(a[281] & b[295])^(a[280] & b[296])^(a[279] & b[297])^(a[278] & b[298])^(a[277] & b[299])^(a[276] & b[300])^(a[275] & b[301])^(a[274] & b[302])^(a[273] & b[303])^(a[272] & b[304])^(a[271] & b[305])^(a[270] & b[306])^(a[269] & b[307])^(a[268] & b[308])^(a[267] & b[309])^(a[266] & b[310])^(a[265] & b[311])^(a[264] & b[312])^(a[263] & b[313])^(a[262] & b[314])^(a[261] & b[315])^(a[260] & b[316])^(a[259] & b[317])^(a[258] & b[318])^(a[257] & b[319])^(a[256] & b[320])^(a[255] & b[321])^(a[254] & b[322])^(a[253] & b[323])^(a[252] & b[324])^(a[251] & b[325])^(a[250] & b[326])^(a[249] & b[327])^(a[248] & b[328])^(a[247] & b[329])^(a[246] & b[330])^(a[245] & b[331])^(a[244] & b[332])^(a[243] & b[333])^(a[242] & b[334])^(a[241] & b[335])^(a[240] & b[336])^(a[239] & b[337])^(a[238] & b[338])^(a[237] & b[339])^(a[236] & b[340])^(a[235] & b[341])^(a[234] & b[342])^(a[233] & b[343])^(a[232] & b[344])^(a[231] & b[345])^(a[230] & b[346])^(a[229] & b[347])^(a[228] & b[348])^(a[227] & b[349])^(a[226] & b[350])^(a[225] & b[351])^(a[224] & b[352])^(a[223] & b[353])^(a[222] & b[354])^(a[221] & b[355])^(a[220] & b[356])^(a[219] & b[357])^(a[218] & b[358])^(a[217] & b[359])^(a[216] & b[360])^(a[215] & b[361])^(a[214] & b[362])^(a[213] & b[363])^(a[212] & b[364])^(a[211] & b[365])^(a[210] & b[366])^(a[209] & b[367])^(a[208] & b[368])^(a[207] & b[369])^(a[206] & b[370])^(a[205] & b[371])^(a[204] & b[372])^(a[203] & b[373])^(a[202] & b[374])^(a[201] & b[375])^(a[200] & b[376])^(a[199] & b[377])^(a[198] & b[378])^(a[197] & b[379])^(a[196] & b[380])^(a[195] & b[381])^(a[194] & b[382])^(a[193] & b[383])^(a[192] & b[384])^(a[191] & b[385])^(a[190] & b[386])^(a[189] & b[387])^(a[188] & b[388])^(a[187] & b[389])^(a[186] & b[390])^(a[185] & b[391])^(a[184] & b[392])^(a[183] & b[393])^(a[182] & b[394])^(a[181] & b[395])^(a[180] & b[396])^(a[179] & b[397])^(a[178] & b[398])^(a[177] & b[399])^(a[176] & b[400])^(a[175] & b[401])^(a[174] & b[402])^(a[173] & b[403])^(a[172] & b[404])^(a[171] & b[405])^(a[170] & b[406])^(a[169] & b[407])^(a[168] & b[408]);
assign y[577] = (a[408] & b[169])^(a[407] & b[170])^(a[406] & b[171])^(a[405] & b[172])^(a[404] & b[173])^(a[403] & b[174])^(a[402] & b[175])^(a[401] & b[176])^(a[400] & b[177])^(a[399] & b[178])^(a[398] & b[179])^(a[397] & b[180])^(a[396] & b[181])^(a[395] & b[182])^(a[394] & b[183])^(a[393] & b[184])^(a[392] & b[185])^(a[391] & b[186])^(a[390] & b[187])^(a[389] & b[188])^(a[388] & b[189])^(a[387] & b[190])^(a[386] & b[191])^(a[385] & b[192])^(a[384] & b[193])^(a[383] & b[194])^(a[382] & b[195])^(a[381] & b[196])^(a[380] & b[197])^(a[379] & b[198])^(a[378] & b[199])^(a[377] & b[200])^(a[376] & b[201])^(a[375] & b[202])^(a[374] & b[203])^(a[373] & b[204])^(a[372] & b[205])^(a[371] & b[206])^(a[370] & b[207])^(a[369] & b[208])^(a[368] & b[209])^(a[367] & b[210])^(a[366] & b[211])^(a[365] & b[212])^(a[364] & b[213])^(a[363] & b[214])^(a[362] & b[215])^(a[361] & b[216])^(a[360] & b[217])^(a[359] & b[218])^(a[358] & b[219])^(a[357] & b[220])^(a[356] & b[221])^(a[355] & b[222])^(a[354] & b[223])^(a[353] & b[224])^(a[352] & b[225])^(a[351] & b[226])^(a[350] & b[227])^(a[349] & b[228])^(a[348] & b[229])^(a[347] & b[230])^(a[346] & b[231])^(a[345] & b[232])^(a[344] & b[233])^(a[343] & b[234])^(a[342] & b[235])^(a[341] & b[236])^(a[340] & b[237])^(a[339] & b[238])^(a[338] & b[239])^(a[337] & b[240])^(a[336] & b[241])^(a[335] & b[242])^(a[334] & b[243])^(a[333] & b[244])^(a[332] & b[245])^(a[331] & b[246])^(a[330] & b[247])^(a[329] & b[248])^(a[328] & b[249])^(a[327] & b[250])^(a[326] & b[251])^(a[325] & b[252])^(a[324] & b[253])^(a[323] & b[254])^(a[322] & b[255])^(a[321] & b[256])^(a[320] & b[257])^(a[319] & b[258])^(a[318] & b[259])^(a[317] & b[260])^(a[316] & b[261])^(a[315] & b[262])^(a[314] & b[263])^(a[313] & b[264])^(a[312] & b[265])^(a[311] & b[266])^(a[310] & b[267])^(a[309] & b[268])^(a[308] & b[269])^(a[307] & b[270])^(a[306] & b[271])^(a[305] & b[272])^(a[304] & b[273])^(a[303] & b[274])^(a[302] & b[275])^(a[301] & b[276])^(a[300] & b[277])^(a[299] & b[278])^(a[298] & b[279])^(a[297] & b[280])^(a[296] & b[281])^(a[295] & b[282])^(a[294] & b[283])^(a[293] & b[284])^(a[292] & b[285])^(a[291] & b[286])^(a[290] & b[287])^(a[289] & b[288])^(a[288] & b[289])^(a[287] & b[290])^(a[286] & b[291])^(a[285] & b[292])^(a[284] & b[293])^(a[283] & b[294])^(a[282] & b[295])^(a[281] & b[296])^(a[280] & b[297])^(a[279] & b[298])^(a[278] & b[299])^(a[277] & b[300])^(a[276] & b[301])^(a[275] & b[302])^(a[274] & b[303])^(a[273] & b[304])^(a[272] & b[305])^(a[271] & b[306])^(a[270] & b[307])^(a[269] & b[308])^(a[268] & b[309])^(a[267] & b[310])^(a[266] & b[311])^(a[265] & b[312])^(a[264] & b[313])^(a[263] & b[314])^(a[262] & b[315])^(a[261] & b[316])^(a[260] & b[317])^(a[259] & b[318])^(a[258] & b[319])^(a[257] & b[320])^(a[256] & b[321])^(a[255] & b[322])^(a[254] & b[323])^(a[253] & b[324])^(a[252] & b[325])^(a[251] & b[326])^(a[250] & b[327])^(a[249] & b[328])^(a[248] & b[329])^(a[247] & b[330])^(a[246] & b[331])^(a[245] & b[332])^(a[244] & b[333])^(a[243] & b[334])^(a[242] & b[335])^(a[241] & b[336])^(a[240] & b[337])^(a[239] & b[338])^(a[238] & b[339])^(a[237] & b[340])^(a[236] & b[341])^(a[235] & b[342])^(a[234] & b[343])^(a[233] & b[344])^(a[232] & b[345])^(a[231] & b[346])^(a[230] & b[347])^(a[229] & b[348])^(a[228] & b[349])^(a[227] & b[350])^(a[226] & b[351])^(a[225] & b[352])^(a[224] & b[353])^(a[223] & b[354])^(a[222] & b[355])^(a[221] & b[356])^(a[220] & b[357])^(a[219] & b[358])^(a[218] & b[359])^(a[217] & b[360])^(a[216] & b[361])^(a[215] & b[362])^(a[214] & b[363])^(a[213] & b[364])^(a[212] & b[365])^(a[211] & b[366])^(a[210] & b[367])^(a[209] & b[368])^(a[208] & b[369])^(a[207] & b[370])^(a[206] & b[371])^(a[205] & b[372])^(a[204] & b[373])^(a[203] & b[374])^(a[202] & b[375])^(a[201] & b[376])^(a[200] & b[377])^(a[199] & b[378])^(a[198] & b[379])^(a[197] & b[380])^(a[196] & b[381])^(a[195] & b[382])^(a[194] & b[383])^(a[193] & b[384])^(a[192] & b[385])^(a[191] & b[386])^(a[190] & b[387])^(a[189] & b[388])^(a[188] & b[389])^(a[187] & b[390])^(a[186] & b[391])^(a[185] & b[392])^(a[184] & b[393])^(a[183] & b[394])^(a[182] & b[395])^(a[181] & b[396])^(a[180] & b[397])^(a[179] & b[398])^(a[178] & b[399])^(a[177] & b[400])^(a[176] & b[401])^(a[175] & b[402])^(a[174] & b[403])^(a[173] & b[404])^(a[172] & b[405])^(a[171] & b[406])^(a[170] & b[407])^(a[169] & b[408]);
assign y[578] = (a[408] & b[170])^(a[407] & b[171])^(a[406] & b[172])^(a[405] & b[173])^(a[404] & b[174])^(a[403] & b[175])^(a[402] & b[176])^(a[401] & b[177])^(a[400] & b[178])^(a[399] & b[179])^(a[398] & b[180])^(a[397] & b[181])^(a[396] & b[182])^(a[395] & b[183])^(a[394] & b[184])^(a[393] & b[185])^(a[392] & b[186])^(a[391] & b[187])^(a[390] & b[188])^(a[389] & b[189])^(a[388] & b[190])^(a[387] & b[191])^(a[386] & b[192])^(a[385] & b[193])^(a[384] & b[194])^(a[383] & b[195])^(a[382] & b[196])^(a[381] & b[197])^(a[380] & b[198])^(a[379] & b[199])^(a[378] & b[200])^(a[377] & b[201])^(a[376] & b[202])^(a[375] & b[203])^(a[374] & b[204])^(a[373] & b[205])^(a[372] & b[206])^(a[371] & b[207])^(a[370] & b[208])^(a[369] & b[209])^(a[368] & b[210])^(a[367] & b[211])^(a[366] & b[212])^(a[365] & b[213])^(a[364] & b[214])^(a[363] & b[215])^(a[362] & b[216])^(a[361] & b[217])^(a[360] & b[218])^(a[359] & b[219])^(a[358] & b[220])^(a[357] & b[221])^(a[356] & b[222])^(a[355] & b[223])^(a[354] & b[224])^(a[353] & b[225])^(a[352] & b[226])^(a[351] & b[227])^(a[350] & b[228])^(a[349] & b[229])^(a[348] & b[230])^(a[347] & b[231])^(a[346] & b[232])^(a[345] & b[233])^(a[344] & b[234])^(a[343] & b[235])^(a[342] & b[236])^(a[341] & b[237])^(a[340] & b[238])^(a[339] & b[239])^(a[338] & b[240])^(a[337] & b[241])^(a[336] & b[242])^(a[335] & b[243])^(a[334] & b[244])^(a[333] & b[245])^(a[332] & b[246])^(a[331] & b[247])^(a[330] & b[248])^(a[329] & b[249])^(a[328] & b[250])^(a[327] & b[251])^(a[326] & b[252])^(a[325] & b[253])^(a[324] & b[254])^(a[323] & b[255])^(a[322] & b[256])^(a[321] & b[257])^(a[320] & b[258])^(a[319] & b[259])^(a[318] & b[260])^(a[317] & b[261])^(a[316] & b[262])^(a[315] & b[263])^(a[314] & b[264])^(a[313] & b[265])^(a[312] & b[266])^(a[311] & b[267])^(a[310] & b[268])^(a[309] & b[269])^(a[308] & b[270])^(a[307] & b[271])^(a[306] & b[272])^(a[305] & b[273])^(a[304] & b[274])^(a[303] & b[275])^(a[302] & b[276])^(a[301] & b[277])^(a[300] & b[278])^(a[299] & b[279])^(a[298] & b[280])^(a[297] & b[281])^(a[296] & b[282])^(a[295] & b[283])^(a[294] & b[284])^(a[293] & b[285])^(a[292] & b[286])^(a[291] & b[287])^(a[290] & b[288])^(a[289] & b[289])^(a[288] & b[290])^(a[287] & b[291])^(a[286] & b[292])^(a[285] & b[293])^(a[284] & b[294])^(a[283] & b[295])^(a[282] & b[296])^(a[281] & b[297])^(a[280] & b[298])^(a[279] & b[299])^(a[278] & b[300])^(a[277] & b[301])^(a[276] & b[302])^(a[275] & b[303])^(a[274] & b[304])^(a[273] & b[305])^(a[272] & b[306])^(a[271] & b[307])^(a[270] & b[308])^(a[269] & b[309])^(a[268] & b[310])^(a[267] & b[311])^(a[266] & b[312])^(a[265] & b[313])^(a[264] & b[314])^(a[263] & b[315])^(a[262] & b[316])^(a[261] & b[317])^(a[260] & b[318])^(a[259] & b[319])^(a[258] & b[320])^(a[257] & b[321])^(a[256] & b[322])^(a[255] & b[323])^(a[254] & b[324])^(a[253] & b[325])^(a[252] & b[326])^(a[251] & b[327])^(a[250] & b[328])^(a[249] & b[329])^(a[248] & b[330])^(a[247] & b[331])^(a[246] & b[332])^(a[245] & b[333])^(a[244] & b[334])^(a[243] & b[335])^(a[242] & b[336])^(a[241] & b[337])^(a[240] & b[338])^(a[239] & b[339])^(a[238] & b[340])^(a[237] & b[341])^(a[236] & b[342])^(a[235] & b[343])^(a[234] & b[344])^(a[233] & b[345])^(a[232] & b[346])^(a[231] & b[347])^(a[230] & b[348])^(a[229] & b[349])^(a[228] & b[350])^(a[227] & b[351])^(a[226] & b[352])^(a[225] & b[353])^(a[224] & b[354])^(a[223] & b[355])^(a[222] & b[356])^(a[221] & b[357])^(a[220] & b[358])^(a[219] & b[359])^(a[218] & b[360])^(a[217] & b[361])^(a[216] & b[362])^(a[215] & b[363])^(a[214] & b[364])^(a[213] & b[365])^(a[212] & b[366])^(a[211] & b[367])^(a[210] & b[368])^(a[209] & b[369])^(a[208] & b[370])^(a[207] & b[371])^(a[206] & b[372])^(a[205] & b[373])^(a[204] & b[374])^(a[203] & b[375])^(a[202] & b[376])^(a[201] & b[377])^(a[200] & b[378])^(a[199] & b[379])^(a[198] & b[380])^(a[197] & b[381])^(a[196] & b[382])^(a[195] & b[383])^(a[194] & b[384])^(a[193] & b[385])^(a[192] & b[386])^(a[191] & b[387])^(a[190] & b[388])^(a[189] & b[389])^(a[188] & b[390])^(a[187] & b[391])^(a[186] & b[392])^(a[185] & b[393])^(a[184] & b[394])^(a[183] & b[395])^(a[182] & b[396])^(a[181] & b[397])^(a[180] & b[398])^(a[179] & b[399])^(a[178] & b[400])^(a[177] & b[401])^(a[176] & b[402])^(a[175] & b[403])^(a[174] & b[404])^(a[173] & b[405])^(a[172] & b[406])^(a[171] & b[407])^(a[170] & b[408]);
assign y[579] = (a[408] & b[171])^(a[407] & b[172])^(a[406] & b[173])^(a[405] & b[174])^(a[404] & b[175])^(a[403] & b[176])^(a[402] & b[177])^(a[401] & b[178])^(a[400] & b[179])^(a[399] & b[180])^(a[398] & b[181])^(a[397] & b[182])^(a[396] & b[183])^(a[395] & b[184])^(a[394] & b[185])^(a[393] & b[186])^(a[392] & b[187])^(a[391] & b[188])^(a[390] & b[189])^(a[389] & b[190])^(a[388] & b[191])^(a[387] & b[192])^(a[386] & b[193])^(a[385] & b[194])^(a[384] & b[195])^(a[383] & b[196])^(a[382] & b[197])^(a[381] & b[198])^(a[380] & b[199])^(a[379] & b[200])^(a[378] & b[201])^(a[377] & b[202])^(a[376] & b[203])^(a[375] & b[204])^(a[374] & b[205])^(a[373] & b[206])^(a[372] & b[207])^(a[371] & b[208])^(a[370] & b[209])^(a[369] & b[210])^(a[368] & b[211])^(a[367] & b[212])^(a[366] & b[213])^(a[365] & b[214])^(a[364] & b[215])^(a[363] & b[216])^(a[362] & b[217])^(a[361] & b[218])^(a[360] & b[219])^(a[359] & b[220])^(a[358] & b[221])^(a[357] & b[222])^(a[356] & b[223])^(a[355] & b[224])^(a[354] & b[225])^(a[353] & b[226])^(a[352] & b[227])^(a[351] & b[228])^(a[350] & b[229])^(a[349] & b[230])^(a[348] & b[231])^(a[347] & b[232])^(a[346] & b[233])^(a[345] & b[234])^(a[344] & b[235])^(a[343] & b[236])^(a[342] & b[237])^(a[341] & b[238])^(a[340] & b[239])^(a[339] & b[240])^(a[338] & b[241])^(a[337] & b[242])^(a[336] & b[243])^(a[335] & b[244])^(a[334] & b[245])^(a[333] & b[246])^(a[332] & b[247])^(a[331] & b[248])^(a[330] & b[249])^(a[329] & b[250])^(a[328] & b[251])^(a[327] & b[252])^(a[326] & b[253])^(a[325] & b[254])^(a[324] & b[255])^(a[323] & b[256])^(a[322] & b[257])^(a[321] & b[258])^(a[320] & b[259])^(a[319] & b[260])^(a[318] & b[261])^(a[317] & b[262])^(a[316] & b[263])^(a[315] & b[264])^(a[314] & b[265])^(a[313] & b[266])^(a[312] & b[267])^(a[311] & b[268])^(a[310] & b[269])^(a[309] & b[270])^(a[308] & b[271])^(a[307] & b[272])^(a[306] & b[273])^(a[305] & b[274])^(a[304] & b[275])^(a[303] & b[276])^(a[302] & b[277])^(a[301] & b[278])^(a[300] & b[279])^(a[299] & b[280])^(a[298] & b[281])^(a[297] & b[282])^(a[296] & b[283])^(a[295] & b[284])^(a[294] & b[285])^(a[293] & b[286])^(a[292] & b[287])^(a[291] & b[288])^(a[290] & b[289])^(a[289] & b[290])^(a[288] & b[291])^(a[287] & b[292])^(a[286] & b[293])^(a[285] & b[294])^(a[284] & b[295])^(a[283] & b[296])^(a[282] & b[297])^(a[281] & b[298])^(a[280] & b[299])^(a[279] & b[300])^(a[278] & b[301])^(a[277] & b[302])^(a[276] & b[303])^(a[275] & b[304])^(a[274] & b[305])^(a[273] & b[306])^(a[272] & b[307])^(a[271] & b[308])^(a[270] & b[309])^(a[269] & b[310])^(a[268] & b[311])^(a[267] & b[312])^(a[266] & b[313])^(a[265] & b[314])^(a[264] & b[315])^(a[263] & b[316])^(a[262] & b[317])^(a[261] & b[318])^(a[260] & b[319])^(a[259] & b[320])^(a[258] & b[321])^(a[257] & b[322])^(a[256] & b[323])^(a[255] & b[324])^(a[254] & b[325])^(a[253] & b[326])^(a[252] & b[327])^(a[251] & b[328])^(a[250] & b[329])^(a[249] & b[330])^(a[248] & b[331])^(a[247] & b[332])^(a[246] & b[333])^(a[245] & b[334])^(a[244] & b[335])^(a[243] & b[336])^(a[242] & b[337])^(a[241] & b[338])^(a[240] & b[339])^(a[239] & b[340])^(a[238] & b[341])^(a[237] & b[342])^(a[236] & b[343])^(a[235] & b[344])^(a[234] & b[345])^(a[233] & b[346])^(a[232] & b[347])^(a[231] & b[348])^(a[230] & b[349])^(a[229] & b[350])^(a[228] & b[351])^(a[227] & b[352])^(a[226] & b[353])^(a[225] & b[354])^(a[224] & b[355])^(a[223] & b[356])^(a[222] & b[357])^(a[221] & b[358])^(a[220] & b[359])^(a[219] & b[360])^(a[218] & b[361])^(a[217] & b[362])^(a[216] & b[363])^(a[215] & b[364])^(a[214] & b[365])^(a[213] & b[366])^(a[212] & b[367])^(a[211] & b[368])^(a[210] & b[369])^(a[209] & b[370])^(a[208] & b[371])^(a[207] & b[372])^(a[206] & b[373])^(a[205] & b[374])^(a[204] & b[375])^(a[203] & b[376])^(a[202] & b[377])^(a[201] & b[378])^(a[200] & b[379])^(a[199] & b[380])^(a[198] & b[381])^(a[197] & b[382])^(a[196] & b[383])^(a[195] & b[384])^(a[194] & b[385])^(a[193] & b[386])^(a[192] & b[387])^(a[191] & b[388])^(a[190] & b[389])^(a[189] & b[390])^(a[188] & b[391])^(a[187] & b[392])^(a[186] & b[393])^(a[185] & b[394])^(a[184] & b[395])^(a[183] & b[396])^(a[182] & b[397])^(a[181] & b[398])^(a[180] & b[399])^(a[179] & b[400])^(a[178] & b[401])^(a[177] & b[402])^(a[176] & b[403])^(a[175] & b[404])^(a[174] & b[405])^(a[173] & b[406])^(a[172] & b[407])^(a[171] & b[408]);
assign y[580] = (a[408] & b[172])^(a[407] & b[173])^(a[406] & b[174])^(a[405] & b[175])^(a[404] & b[176])^(a[403] & b[177])^(a[402] & b[178])^(a[401] & b[179])^(a[400] & b[180])^(a[399] & b[181])^(a[398] & b[182])^(a[397] & b[183])^(a[396] & b[184])^(a[395] & b[185])^(a[394] & b[186])^(a[393] & b[187])^(a[392] & b[188])^(a[391] & b[189])^(a[390] & b[190])^(a[389] & b[191])^(a[388] & b[192])^(a[387] & b[193])^(a[386] & b[194])^(a[385] & b[195])^(a[384] & b[196])^(a[383] & b[197])^(a[382] & b[198])^(a[381] & b[199])^(a[380] & b[200])^(a[379] & b[201])^(a[378] & b[202])^(a[377] & b[203])^(a[376] & b[204])^(a[375] & b[205])^(a[374] & b[206])^(a[373] & b[207])^(a[372] & b[208])^(a[371] & b[209])^(a[370] & b[210])^(a[369] & b[211])^(a[368] & b[212])^(a[367] & b[213])^(a[366] & b[214])^(a[365] & b[215])^(a[364] & b[216])^(a[363] & b[217])^(a[362] & b[218])^(a[361] & b[219])^(a[360] & b[220])^(a[359] & b[221])^(a[358] & b[222])^(a[357] & b[223])^(a[356] & b[224])^(a[355] & b[225])^(a[354] & b[226])^(a[353] & b[227])^(a[352] & b[228])^(a[351] & b[229])^(a[350] & b[230])^(a[349] & b[231])^(a[348] & b[232])^(a[347] & b[233])^(a[346] & b[234])^(a[345] & b[235])^(a[344] & b[236])^(a[343] & b[237])^(a[342] & b[238])^(a[341] & b[239])^(a[340] & b[240])^(a[339] & b[241])^(a[338] & b[242])^(a[337] & b[243])^(a[336] & b[244])^(a[335] & b[245])^(a[334] & b[246])^(a[333] & b[247])^(a[332] & b[248])^(a[331] & b[249])^(a[330] & b[250])^(a[329] & b[251])^(a[328] & b[252])^(a[327] & b[253])^(a[326] & b[254])^(a[325] & b[255])^(a[324] & b[256])^(a[323] & b[257])^(a[322] & b[258])^(a[321] & b[259])^(a[320] & b[260])^(a[319] & b[261])^(a[318] & b[262])^(a[317] & b[263])^(a[316] & b[264])^(a[315] & b[265])^(a[314] & b[266])^(a[313] & b[267])^(a[312] & b[268])^(a[311] & b[269])^(a[310] & b[270])^(a[309] & b[271])^(a[308] & b[272])^(a[307] & b[273])^(a[306] & b[274])^(a[305] & b[275])^(a[304] & b[276])^(a[303] & b[277])^(a[302] & b[278])^(a[301] & b[279])^(a[300] & b[280])^(a[299] & b[281])^(a[298] & b[282])^(a[297] & b[283])^(a[296] & b[284])^(a[295] & b[285])^(a[294] & b[286])^(a[293] & b[287])^(a[292] & b[288])^(a[291] & b[289])^(a[290] & b[290])^(a[289] & b[291])^(a[288] & b[292])^(a[287] & b[293])^(a[286] & b[294])^(a[285] & b[295])^(a[284] & b[296])^(a[283] & b[297])^(a[282] & b[298])^(a[281] & b[299])^(a[280] & b[300])^(a[279] & b[301])^(a[278] & b[302])^(a[277] & b[303])^(a[276] & b[304])^(a[275] & b[305])^(a[274] & b[306])^(a[273] & b[307])^(a[272] & b[308])^(a[271] & b[309])^(a[270] & b[310])^(a[269] & b[311])^(a[268] & b[312])^(a[267] & b[313])^(a[266] & b[314])^(a[265] & b[315])^(a[264] & b[316])^(a[263] & b[317])^(a[262] & b[318])^(a[261] & b[319])^(a[260] & b[320])^(a[259] & b[321])^(a[258] & b[322])^(a[257] & b[323])^(a[256] & b[324])^(a[255] & b[325])^(a[254] & b[326])^(a[253] & b[327])^(a[252] & b[328])^(a[251] & b[329])^(a[250] & b[330])^(a[249] & b[331])^(a[248] & b[332])^(a[247] & b[333])^(a[246] & b[334])^(a[245] & b[335])^(a[244] & b[336])^(a[243] & b[337])^(a[242] & b[338])^(a[241] & b[339])^(a[240] & b[340])^(a[239] & b[341])^(a[238] & b[342])^(a[237] & b[343])^(a[236] & b[344])^(a[235] & b[345])^(a[234] & b[346])^(a[233] & b[347])^(a[232] & b[348])^(a[231] & b[349])^(a[230] & b[350])^(a[229] & b[351])^(a[228] & b[352])^(a[227] & b[353])^(a[226] & b[354])^(a[225] & b[355])^(a[224] & b[356])^(a[223] & b[357])^(a[222] & b[358])^(a[221] & b[359])^(a[220] & b[360])^(a[219] & b[361])^(a[218] & b[362])^(a[217] & b[363])^(a[216] & b[364])^(a[215] & b[365])^(a[214] & b[366])^(a[213] & b[367])^(a[212] & b[368])^(a[211] & b[369])^(a[210] & b[370])^(a[209] & b[371])^(a[208] & b[372])^(a[207] & b[373])^(a[206] & b[374])^(a[205] & b[375])^(a[204] & b[376])^(a[203] & b[377])^(a[202] & b[378])^(a[201] & b[379])^(a[200] & b[380])^(a[199] & b[381])^(a[198] & b[382])^(a[197] & b[383])^(a[196] & b[384])^(a[195] & b[385])^(a[194] & b[386])^(a[193] & b[387])^(a[192] & b[388])^(a[191] & b[389])^(a[190] & b[390])^(a[189] & b[391])^(a[188] & b[392])^(a[187] & b[393])^(a[186] & b[394])^(a[185] & b[395])^(a[184] & b[396])^(a[183] & b[397])^(a[182] & b[398])^(a[181] & b[399])^(a[180] & b[400])^(a[179] & b[401])^(a[178] & b[402])^(a[177] & b[403])^(a[176] & b[404])^(a[175] & b[405])^(a[174] & b[406])^(a[173] & b[407])^(a[172] & b[408]);
assign y[581] = (a[408] & b[173])^(a[407] & b[174])^(a[406] & b[175])^(a[405] & b[176])^(a[404] & b[177])^(a[403] & b[178])^(a[402] & b[179])^(a[401] & b[180])^(a[400] & b[181])^(a[399] & b[182])^(a[398] & b[183])^(a[397] & b[184])^(a[396] & b[185])^(a[395] & b[186])^(a[394] & b[187])^(a[393] & b[188])^(a[392] & b[189])^(a[391] & b[190])^(a[390] & b[191])^(a[389] & b[192])^(a[388] & b[193])^(a[387] & b[194])^(a[386] & b[195])^(a[385] & b[196])^(a[384] & b[197])^(a[383] & b[198])^(a[382] & b[199])^(a[381] & b[200])^(a[380] & b[201])^(a[379] & b[202])^(a[378] & b[203])^(a[377] & b[204])^(a[376] & b[205])^(a[375] & b[206])^(a[374] & b[207])^(a[373] & b[208])^(a[372] & b[209])^(a[371] & b[210])^(a[370] & b[211])^(a[369] & b[212])^(a[368] & b[213])^(a[367] & b[214])^(a[366] & b[215])^(a[365] & b[216])^(a[364] & b[217])^(a[363] & b[218])^(a[362] & b[219])^(a[361] & b[220])^(a[360] & b[221])^(a[359] & b[222])^(a[358] & b[223])^(a[357] & b[224])^(a[356] & b[225])^(a[355] & b[226])^(a[354] & b[227])^(a[353] & b[228])^(a[352] & b[229])^(a[351] & b[230])^(a[350] & b[231])^(a[349] & b[232])^(a[348] & b[233])^(a[347] & b[234])^(a[346] & b[235])^(a[345] & b[236])^(a[344] & b[237])^(a[343] & b[238])^(a[342] & b[239])^(a[341] & b[240])^(a[340] & b[241])^(a[339] & b[242])^(a[338] & b[243])^(a[337] & b[244])^(a[336] & b[245])^(a[335] & b[246])^(a[334] & b[247])^(a[333] & b[248])^(a[332] & b[249])^(a[331] & b[250])^(a[330] & b[251])^(a[329] & b[252])^(a[328] & b[253])^(a[327] & b[254])^(a[326] & b[255])^(a[325] & b[256])^(a[324] & b[257])^(a[323] & b[258])^(a[322] & b[259])^(a[321] & b[260])^(a[320] & b[261])^(a[319] & b[262])^(a[318] & b[263])^(a[317] & b[264])^(a[316] & b[265])^(a[315] & b[266])^(a[314] & b[267])^(a[313] & b[268])^(a[312] & b[269])^(a[311] & b[270])^(a[310] & b[271])^(a[309] & b[272])^(a[308] & b[273])^(a[307] & b[274])^(a[306] & b[275])^(a[305] & b[276])^(a[304] & b[277])^(a[303] & b[278])^(a[302] & b[279])^(a[301] & b[280])^(a[300] & b[281])^(a[299] & b[282])^(a[298] & b[283])^(a[297] & b[284])^(a[296] & b[285])^(a[295] & b[286])^(a[294] & b[287])^(a[293] & b[288])^(a[292] & b[289])^(a[291] & b[290])^(a[290] & b[291])^(a[289] & b[292])^(a[288] & b[293])^(a[287] & b[294])^(a[286] & b[295])^(a[285] & b[296])^(a[284] & b[297])^(a[283] & b[298])^(a[282] & b[299])^(a[281] & b[300])^(a[280] & b[301])^(a[279] & b[302])^(a[278] & b[303])^(a[277] & b[304])^(a[276] & b[305])^(a[275] & b[306])^(a[274] & b[307])^(a[273] & b[308])^(a[272] & b[309])^(a[271] & b[310])^(a[270] & b[311])^(a[269] & b[312])^(a[268] & b[313])^(a[267] & b[314])^(a[266] & b[315])^(a[265] & b[316])^(a[264] & b[317])^(a[263] & b[318])^(a[262] & b[319])^(a[261] & b[320])^(a[260] & b[321])^(a[259] & b[322])^(a[258] & b[323])^(a[257] & b[324])^(a[256] & b[325])^(a[255] & b[326])^(a[254] & b[327])^(a[253] & b[328])^(a[252] & b[329])^(a[251] & b[330])^(a[250] & b[331])^(a[249] & b[332])^(a[248] & b[333])^(a[247] & b[334])^(a[246] & b[335])^(a[245] & b[336])^(a[244] & b[337])^(a[243] & b[338])^(a[242] & b[339])^(a[241] & b[340])^(a[240] & b[341])^(a[239] & b[342])^(a[238] & b[343])^(a[237] & b[344])^(a[236] & b[345])^(a[235] & b[346])^(a[234] & b[347])^(a[233] & b[348])^(a[232] & b[349])^(a[231] & b[350])^(a[230] & b[351])^(a[229] & b[352])^(a[228] & b[353])^(a[227] & b[354])^(a[226] & b[355])^(a[225] & b[356])^(a[224] & b[357])^(a[223] & b[358])^(a[222] & b[359])^(a[221] & b[360])^(a[220] & b[361])^(a[219] & b[362])^(a[218] & b[363])^(a[217] & b[364])^(a[216] & b[365])^(a[215] & b[366])^(a[214] & b[367])^(a[213] & b[368])^(a[212] & b[369])^(a[211] & b[370])^(a[210] & b[371])^(a[209] & b[372])^(a[208] & b[373])^(a[207] & b[374])^(a[206] & b[375])^(a[205] & b[376])^(a[204] & b[377])^(a[203] & b[378])^(a[202] & b[379])^(a[201] & b[380])^(a[200] & b[381])^(a[199] & b[382])^(a[198] & b[383])^(a[197] & b[384])^(a[196] & b[385])^(a[195] & b[386])^(a[194] & b[387])^(a[193] & b[388])^(a[192] & b[389])^(a[191] & b[390])^(a[190] & b[391])^(a[189] & b[392])^(a[188] & b[393])^(a[187] & b[394])^(a[186] & b[395])^(a[185] & b[396])^(a[184] & b[397])^(a[183] & b[398])^(a[182] & b[399])^(a[181] & b[400])^(a[180] & b[401])^(a[179] & b[402])^(a[178] & b[403])^(a[177] & b[404])^(a[176] & b[405])^(a[175] & b[406])^(a[174] & b[407])^(a[173] & b[408]);
assign y[582] = (a[408] & b[174])^(a[407] & b[175])^(a[406] & b[176])^(a[405] & b[177])^(a[404] & b[178])^(a[403] & b[179])^(a[402] & b[180])^(a[401] & b[181])^(a[400] & b[182])^(a[399] & b[183])^(a[398] & b[184])^(a[397] & b[185])^(a[396] & b[186])^(a[395] & b[187])^(a[394] & b[188])^(a[393] & b[189])^(a[392] & b[190])^(a[391] & b[191])^(a[390] & b[192])^(a[389] & b[193])^(a[388] & b[194])^(a[387] & b[195])^(a[386] & b[196])^(a[385] & b[197])^(a[384] & b[198])^(a[383] & b[199])^(a[382] & b[200])^(a[381] & b[201])^(a[380] & b[202])^(a[379] & b[203])^(a[378] & b[204])^(a[377] & b[205])^(a[376] & b[206])^(a[375] & b[207])^(a[374] & b[208])^(a[373] & b[209])^(a[372] & b[210])^(a[371] & b[211])^(a[370] & b[212])^(a[369] & b[213])^(a[368] & b[214])^(a[367] & b[215])^(a[366] & b[216])^(a[365] & b[217])^(a[364] & b[218])^(a[363] & b[219])^(a[362] & b[220])^(a[361] & b[221])^(a[360] & b[222])^(a[359] & b[223])^(a[358] & b[224])^(a[357] & b[225])^(a[356] & b[226])^(a[355] & b[227])^(a[354] & b[228])^(a[353] & b[229])^(a[352] & b[230])^(a[351] & b[231])^(a[350] & b[232])^(a[349] & b[233])^(a[348] & b[234])^(a[347] & b[235])^(a[346] & b[236])^(a[345] & b[237])^(a[344] & b[238])^(a[343] & b[239])^(a[342] & b[240])^(a[341] & b[241])^(a[340] & b[242])^(a[339] & b[243])^(a[338] & b[244])^(a[337] & b[245])^(a[336] & b[246])^(a[335] & b[247])^(a[334] & b[248])^(a[333] & b[249])^(a[332] & b[250])^(a[331] & b[251])^(a[330] & b[252])^(a[329] & b[253])^(a[328] & b[254])^(a[327] & b[255])^(a[326] & b[256])^(a[325] & b[257])^(a[324] & b[258])^(a[323] & b[259])^(a[322] & b[260])^(a[321] & b[261])^(a[320] & b[262])^(a[319] & b[263])^(a[318] & b[264])^(a[317] & b[265])^(a[316] & b[266])^(a[315] & b[267])^(a[314] & b[268])^(a[313] & b[269])^(a[312] & b[270])^(a[311] & b[271])^(a[310] & b[272])^(a[309] & b[273])^(a[308] & b[274])^(a[307] & b[275])^(a[306] & b[276])^(a[305] & b[277])^(a[304] & b[278])^(a[303] & b[279])^(a[302] & b[280])^(a[301] & b[281])^(a[300] & b[282])^(a[299] & b[283])^(a[298] & b[284])^(a[297] & b[285])^(a[296] & b[286])^(a[295] & b[287])^(a[294] & b[288])^(a[293] & b[289])^(a[292] & b[290])^(a[291] & b[291])^(a[290] & b[292])^(a[289] & b[293])^(a[288] & b[294])^(a[287] & b[295])^(a[286] & b[296])^(a[285] & b[297])^(a[284] & b[298])^(a[283] & b[299])^(a[282] & b[300])^(a[281] & b[301])^(a[280] & b[302])^(a[279] & b[303])^(a[278] & b[304])^(a[277] & b[305])^(a[276] & b[306])^(a[275] & b[307])^(a[274] & b[308])^(a[273] & b[309])^(a[272] & b[310])^(a[271] & b[311])^(a[270] & b[312])^(a[269] & b[313])^(a[268] & b[314])^(a[267] & b[315])^(a[266] & b[316])^(a[265] & b[317])^(a[264] & b[318])^(a[263] & b[319])^(a[262] & b[320])^(a[261] & b[321])^(a[260] & b[322])^(a[259] & b[323])^(a[258] & b[324])^(a[257] & b[325])^(a[256] & b[326])^(a[255] & b[327])^(a[254] & b[328])^(a[253] & b[329])^(a[252] & b[330])^(a[251] & b[331])^(a[250] & b[332])^(a[249] & b[333])^(a[248] & b[334])^(a[247] & b[335])^(a[246] & b[336])^(a[245] & b[337])^(a[244] & b[338])^(a[243] & b[339])^(a[242] & b[340])^(a[241] & b[341])^(a[240] & b[342])^(a[239] & b[343])^(a[238] & b[344])^(a[237] & b[345])^(a[236] & b[346])^(a[235] & b[347])^(a[234] & b[348])^(a[233] & b[349])^(a[232] & b[350])^(a[231] & b[351])^(a[230] & b[352])^(a[229] & b[353])^(a[228] & b[354])^(a[227] & b[355])^(a[226] & b[356])^(a[225] & b[357])^(a[224] & b[358])^(a[223] & b[359])^(a[222] & b[360])^(a[221] & b[361])^(a[220] & b[362])^(a[219] & b[363])^(a[218] & b[364])^(a[217] & b[365])^(a[216] & b[366])^(a[215] & b[367])^(a[214] & b[368])^(a[213] & b[369])^(a[212] & b[370])^(a[211] & b[371])^(a[210] & b[372])^(a[209] & b[373])^(a[208] & b[374])^(a[207] & b[375])^(a[206] & b[376])^(a[205] & b[377])^(a[204] & b[378])^(a[203] & b[379])^(a[202] & b[380])^(a[201] & b[381])^(a[200] & b[382])^(a[199] & b[383])^(a[198] & b[384])^(a[197] & b[385])^(a[196] & b[386])^(a[195] & b[387])^(a[194] & b[388])^(a[193] & b[389])^(a[192] & b[390])^(a[191] & b[391])^(a[190] & b[392])^(a[189] & b[393])^(a[188] & b[394])^(a[187] & b[395])^(a[186] & b[396])^(a[185] & b[397])^(a[184] & b[398])^(a[183] & b[399])^(a[182] & b[400])^(a[181] & b[401])^(a[180] & b[402])^(a[179] & b[403])^(a[178] & b[404])^(a[177] & b[405])^(a[176] & b[406])^(a[175] & b[407])^(a[174] & b[408]);
assign y[583] = (a[408] & b[175])^(a[407] & b[176])^(a[406] & b[177])^(a[405] & b[178])^(a[404] & b[179])^(a[403] & b[180])^(a[402] & b[181])^(a[401] & b[182])^(a[400] & b[183])^(a[399] & b[184])^(a[398] & b[185])^(a[397] & b[186])^(a[396] & b[187])^(a[395] & b[188])^(a[394] & b[189])^(a[393] & b[190])^(a[392] & b[191])^(a[391] & b[192])^(a[390] & b[193])^(a[389] & b[194])^(a[388] & b[195])^(a[387] & b[196])^(a[386] & b[197])^(a[385] & b[198])^(a[384] & b[199])^(a[383] & b[200])^(a[382] & b[201])^(a[381] & b[202])^(a[380] & b[203])^(a[379] & b[204])^(a[378] & b[205])^(a[377] & b[206])^(a[376] & b[207])^(a[375] & b[208])^(a[374] & b[209])^(a[373] & b[210])^(a[372] & b[211])^(a[371] & b[212])^(a[370] & b[213])^(a[369] & b[214])^(a[368] & b[215])^(a[367] & b[216])^(a[366] & b[217])^(a[365] & b[218])^(a[364] & b[219])^(a[363] & b[220])^(a[362] & b[221])^(a[361] & b[222])^(a[360] & b[223])^(a[359] & b[224])^(a[358] & b[225])^(a[357] & b[226])^(a[356] & b[227])^(a[355] & b[228])^(a[354] & b[229])^(a[353] & b[230])^(a[352] & b[231])^(a[351] & b[232])^(a[350] & b[233])^(a[349] & b[234])^(a[348] & b[235])^(a[347] & b[236])^(a[346] & b[237])^(a[345] & b[238])^(a[344] & b[239])^(a[343] & b[240])^(a[342] & b[241])^(a[341] & b[242])^(a[340] & b[243])^(a[339] & b[244])^(a[338] & b[245])^(a[337] & b[246])^(a[336] & b[247])^(a[335] & b[248])^(a[334] & b[249])^(a[333] & b[250])^(a[332] & b[251])^(a[331] & b[252])^(a[330] & b[253])^(a[329] & b[254])^(a[328] & b[255])^(a[327] & b[256])^(a[326] & b[257])^(a[325] & b[258])^(a[324] & b[259])^(a[323] & b[260])^(a[322] & b[261])^(a[321] & b[262])^(a[320] & b[263])^(a[319] & b[264])^(a[318] & b[265])^(a[317] & b[266])^(a[316] & b[267])^(a[315] & b[268])^(a[314] & b[269])^(a[313] & b[270])^(a[312] & b[271])^(a[311] & b[272])^(a[310] & b[273])^(a[309] & b[274])^(a[308] & b[275])^(a[307] & b[276])^(a[306] & b[277])^(a[305] & b[278])^(a[304] & b[279])^(a[303] & b[280])^(a[302] & b[281])^(a[301] & b[282])^(a[300] & b[283])^(a[299] & b[284])^(a[298] & b[285])^(a[297] & b[286])^(a[296] & b[287])^(a[295] & b[288])^(a[294] & b[289])^(a[293] & b[290])^(a[292] & b[291])^(a[291] & b[292])^(a[290] & b[293])^(a[289] & b[294])^(a[288] & b[295])^(a[287] & b[296])^(a[286] & b[297])^(a[285] & b[298])^(a[284] & b[299])^(a[283] & b[300])^(a[282] & b[301])^(a[281] & b[302])^(a[280] & b[303])^(a[279] & b[304])^(a[278] & b[305])^(a[277] & b[306])^(a[276] & b[307])^(a[275] & b[308])^(a[274] & b[309])^(a[273] & b[310])^(a[272] & b[311])^(a[271] & b[312])^(a[270] & b[313])^(a[269] & b[314])^(a[268] & b[315])^(a[267] & b[316])^(a[266] & b[317])^(a[265] & b[318])^(a[264] & b[319])^(a[263] & b[320])^(a[262] & b[321])^(a[261] & b[322])^(a[260] & b[323])^(a[259] & b[324])^(a[258] & b[325])^(a[257] & b[326])^(a[256] & b[327])^(a[255] & b[328])^(a[254] & b[329])^(a[253] & b[330])^(a[252] & b[331])^(a[251] & b[332])^(a[250] & b[333])^(a[249] & b[334])^(a[248] & b[335])^(a[247] & b[336])^(a[246] & b[337])^(a[245] & b[338])^(a[244] & b[339])^(a[243] & b[340])^(a[242] & b[341])^(a[241] & b[342])^(a[240] & b[343])^(a[239] & b[344])^(a[238] & b[345])^(a[237] & b[346])^(a[236] & b[347])^(a[235] & b[348])^(a[234] & b[349])^(a[233] & b[350])^(a[232] & b[351])^(a[231] & b[352])^(a[230] & b[353])^(a[229] & b[354])^(a[228] & b[355])^(a[227] & b[356])^(a[226] & b[357])^(a[225] & b[358])^(a[224] & b[359])^(a[223] & b[360])^(a[222] & b[361])^(a[221] & b[362])^(a[220] & b[363])^(a[219] & b[364])^(a[218] & b[365])^(a[217] & b[366])^(a[216] & b[367])^(a[215] & b[368])^(a[214] & b[369])^(a[213] & b[370])^(a[212] & b[371])^(a[211] & b[372])^(a[210] & b[373])^(a[209] & b[374])^(a[208] & b[375])^(a[207] & b[376])^(a[206] & b[377])^(a[205] & b[378])^(a[204] & b[379])^(a[203] & b[380])^(a[202] & b[381])^(a[201] & b[382])^(a[200] & b[383])^(a[199] & b[384])^(a[198] & b[385])^(a[197] & b[386])^(a[196] & b[387])^(a[195] & b[388])^(a[194] & b[389])^(a[193] & b[390])^(a[192] & b[391])^(a[191] & b[392])^(a[190] & b[393])^(a[189] & b[394])^(a[188] & b[395])^(a[187] & b[396])^(a[186] & b[397])^(a[185] & b[398])^(a[184] & b[399])^(a[183] & b[400])^(a[182] & b[401])^(a[181] & b[402])^(a[180] & b[403])^(a[179] & b[404])^(a[178] & b[405])^(a[177] & b[406])^(a[176] & b[407])^(a[175] & b[408]);
assign y[584] = (a[408] & b[176])^(a[407] & b[177])^(a[406] & b[178])^(a[405] & b[179])^(a[404] & b[180])^(a[403] & b[181])^(a[402] & b[182])^(a[401] & b[183])^(a[400] & b[184])^(a[399] & b[185])^(a[398] & b[186])^(a[397] & b[187])^(a[396] & b[188])^(a[395] & b[189])^(a[394] & b[190])^(a[393] & b[191])^(a[392] & b[192])^(a[391] & b[193])^(a[390] & b[194])^(a[389] & b[195])^(a[388] & b[196])^(a[387] & b[197])^(a[386] & b[198])^(a[385] & b[199])^(a[384] & b[200])^(a[383] & b[201])^(a[382] & b[202])^(a[381] & b[203])^(a[380] & b[204])^(a[379] & b[205])^(a[378] & b[206])^(a[377] & b[207])^(a[376] & b[208])^(a[375] & b[209])^(a[374] & b[210])^(a[373] & b[211])^(a[372] & b[212])^(a[371] & b[213])^(a[370] & b[214])^(a[369] & b[215])^(a[368] & b[216])^(a[367] & b[217])^(a[366] & b[218])^(a[365] & b[219])^(a[364] & b[220])^(a[363] & b[221])^(a[362] & b[222])^(a[361] & b[223])^(a[360] & b[224])^(a[359] & b[225])^(a[358] & b[226])^(a[357] & b[227])^(a[356] & b[228])^(a[355] & b[229])^(a[354] & b[230])^(a[353] & b[231])^(a[352] & b[232])^(a[351] & b[233])^(a[350] & b[234])^(a[349] & b[235])^(a[348] & b[236])^(a[347] & b[237])^(a[346] & b[238])^(a[345] & b[239])^(a[344] & b[240])^(a[343] & b[241])^(a[342] & b[242])^(a[341] & b[243])^(a[340] & b[244])^(a[339] & b[245])^(a[338] & b[246])^(a[337] & b[247])^(a[336] & b[248])^(a[335] & b[249])^(a[334] & b[250])^(a[333] & b[251])^(a[332] & b[252])^(a[331] & b[253])^(a[330] & b[254])^(a[329] & b[255])^(a[328] & b[256])^(a[327] & b[257])^(a[326] & b[258])^(a[325] & b[259])^(a[324] & b[260])^(a[323] & b[261])^(a[322] & b[262])^(a[321] & b[263])^(a[320] & b[264])^(a[319] & b[265])^(a[318] & b[266])^(a[317] & b[267])^(a[316] & b[268])^(a[315] & b[269])^(a[314] & b[270])^(a[313] & b[271])^(a[312] & b[272])^(a[311] & b[273])^(a[310] & b[274])^(a[309] & b[275])^(a[308] & b[276])^(a[307] & b[277])^(a[306] & b[278])^(a[305] & b[279])^(a[304] & b[280])^(a[303] & b[281])^(a[302] & b[282])^(a[301] & b[283])^(a[300] & b[284])^(a[299] & b[285])^(a[298] & b[286])^(a[297] & b[287])^(a[296] & b[288])^(a[295] & b[289])^(a[294] & b[290])^(a[293] & b[291])^(a[292] & b[292])^(a[291] & b[293])^(a[290] & b[294])^(a[289] & b[295])^(a[288] & b[296])^(a[287] & b[297])^(a[286] & b[298])^(a[285] & b[299])^(a[284] & b[300])^(a[283] & b[301])^(a[282] & b[302])^(a[281] & b[303])^(a[280] & b[304])^(a[279] & b[305])^(a[278] & b[306])^(a[277] & b[307])^(a[276] & b[308])^(a[275] & b[309])^(a[274] & b[310])^(a[273] & b[311])^(a[272] & b[312])^(a[271] & b[313])^(a[270] & b[314])^(a[269] & b[315])^(a[268] & b[316])^(a[267] & b[317])^(a[266] & b[318])^(a[265] & b[319])^(a[264] & b[320])^(a[263] & b[321])^(a[262] & b[322])^(a[261] & b[323])^(a[260] & b[324])^(a[259] & b[325])^(a[258] & b[326])^(a[257] & b[327])^(a[256] & b[328])^(a[255] & b[329])^(a[254] & b[330])^(a[253] & b[331])^(a[252] & b[332])^(a[251] & b[333])^(a[250] & b[334])^(a[249] & b[335])^(a[248] & b[336])^(a[247] & b[337])^(a[246] & b[338])^(a[245] & b[339])^(a[244] & b[340])^(a[243] & b[341])^(a[242] & b[342])^(a[241] & b[343])^(a[240] & b[344])^(a[239] & b[345])^(a[238] & b[346])^(a[237] & b[347])^(a[236] & b[348])^(a[235] & b[349])^(a[234] & b[350])^(a[233] & b[351])^(a[232] & b[352])^(a[231] & b[353])^(a[230] & b[354])^(a[229] & b[355])^(a[228] & b[356])^(a[227] & b[357])^(a[226] & b[358])^(a[225] & b[359])^(a[224] & b[360])^(a[223] & b[361])^(a[222] & b[362])^(a[221] & b[363])^(a[220] & b[364])^(a[219] & b[365])^(a[218] & b[366])^(a[217] & b[367])^(a[216] & b[368])^(a[215] & b[369])^(a[214] & b[370])^(a[213] & b[371])^(a[212] & b[372])^(a[211] & b[373])^(a[210] & b[374])^(a[209] & b[375])^(a[208] & b[376])^(a[207] & b[377])^(a[206] & b[378])^(a[205] & b[379])^(a[204] & b[380])^(a[203] & b[381])^(a[202] & b[382])^(a[201] & b[383])^(a[200] & b[384])^(a[199] & b[385])^(a[198] & b[386])^(a[197] & b[387])^(a[196] & b[388])^(a[195] & b[389])^(a[194] & b[390])^(a[193] & b[391])^(a[192] & b[392])^(a[191] & b[393])^(a[190] & b[394])^(a[189] & b[395])^(a[188] & b[396])^(a[187] & b[397])^(a[186] & b[398])^(a[185] & b[399])^(a[184] & b[400])^(a[183] & b[401])^(a[182] & b[402])^(a[181] & b[403])^(a[180] & b[404])^(a[179] & b[405])^(a[178] & b[406])^(a[177] & b[407])^(a[176] & b[408]);
assign y[585] = (a[408] & b[177])^(a[407] & b[178])^(a[406] & b[179])^(a[405] & b[180])^(a[404] & b[181])^(a[403] & b[182])^(a[402] & b[183])^(a[401] & b[184])^(a[400] & b[185])^(a[399] & b[186])^(a[398] & b[187])^(a[397] & b[188])^(a[396] & b[189])^(a[395] & b[190])^(a[394] & b[191])^(a[393] & b[192])^(a[392] & b[193])^(a[391] & b[194])^(a[390] & b[195])^(a[389] & b[196])^(a[388] & b[197])^(a[387] & b[198])^(a[386] & b[199])^(a[385] & b[200])^(a[384] & b[201])^(a[383] & b[202])^(a[382] & b[203])^(a[381] & b[204])^(a[380] & b[205])^(a[379] & b[206])^(a[378] & b[207])^(a[377] & b[208])^(a[376] & b[209])^(a[375] & b[210])^(a[374] & b[211])^(a[373] & b[212])^(a[372] & b[213])^(a[371] & b[214])^(a[370] & b[215])^(a[369] & b[216])^(a[368] & b[217])^(a[367] & b[218])^(a[366] & b[219])^(a[365] & b[220])^(a[364] & b[221])^(a[363] & b[222])^(a[362] & b[223])^(a[361] & b[224])^(a[360] & b[225])^(a[359] & b[226])^(a[358] & b[227])^(a[357] & b[228])^(a[356] & b[229])^(a[355] & b[230])^(a[354] & b[231])^(a[353] & b[232])^(a[352] & b[233])^(a[351] & b[234])^(a[350] & b[235])^(a[349] & b[236])^(a[348] & b[237])^(a[347] & b[238])^(a[346] & b[239])^(a[345] & b[240])^(a[344] & b[241])^(a[343] & b[242])^(a[342] & b[243])^(a[341] & b[244])^(a[340] & b[245])^(a[339] & b[246])^(a[338] & b[247])^(a[337] & b[248])^(a[336] & b[249])^(a[335] & b[250])^(a[334] & b[251])^(a[333] & b[252])^(a[332] & b[253])^(a[331] & b[254])^(a[330] & b[255])^(a[329] & b[256])^(a[328] & b[257])^(a[327] & b[258])^(a[326] & b[259])^(a[325] & b[260])^(a[324] & b[261])^(a[323] & b[262])^(a[322] & b[263])^(a[321] & b[264])^(a[320] & b[265])^(a[319] & b[266])^(a[318] & b[267])^(a[317] & b[268])^(a[316] & b[269])^(a[315] & b[270])^(a[314] & b[271])^(a[313] & b[272])^(a[312] & b[273])^(a[311] & b[274])^(a[310] & b[275])^(a[309] & b[276])^(a[308] & b[277])^(a[307] & b[278])^(a[306] & b[279])^(a[305] & b[280])^(a[304] & b[281])^(a[303] & b[282])^(a[302] & b[283])^(a[301] & b[284])^(a[300] & b[285])^(a[299] & b[286])^(a[298] & b[287])^(a[297] & b[288])^(a[296] & b[289])^(a[295] & b[290])^(a[294] & b[291])^(a[293] & b[292])^(a[292] & b[293])^(a[291] & b[294])^(a[290] & b[295])^(a[289] & b[296])^(a[288] & b[297])^(a[287] & b[298])^(a[286] & b[299])^(a[285] & b[300])^(a[284] & b[301])^(a[283] & b[302])^(a[282] & b[303])^(a[281] & b[304])^(a[280] & b[305])^(a[279] & b[306])^(a[278] & b[307])^(a[277] & b[308])^(a[276] & b[309])^(a[275] & b[310])^(a[274] & b[311])^(a[273] & b[312])^(a[272] & b[313])^(a[271] & b[314])^(a[270] & b[315])^(a[269] & b[316])^(a[268] & b[317])^(a[267] & b[318])^(a[266] & b[319])^(a[265] & b[320])^(a[264] & b[321])^(a[263] & b[322])^(a[262] & b[323])^(a[261] & b[324])^(a[260] & b[325])^(a[259] & b[326])^(a[258] & b[327])^(a[257] & b[328])^(a[256] & b[329])^(a[255] & b[330])^(a[254] & b[331])^(a[253] & b[332])^(a[252] & b[333])^(a[251] & b[334])^(a[250] & b[335])^(a[249] & b[336])^(a[248] & b[337])^(a[247] & b[338])^(a[246] & b[339])^(a[245] & b[340])^(a[244] & b[341])^(a[243] & b[342])^(a[242] & b[343])^(a[241] & b[344])^(a[240] & b[345])^(a[239] & b[346])^(a[238] & b[347])^(a[237] & b[348])^(a[236] & b[349])^(a[235] & b[350])^(a[234] & b[351])^(a[233] & b[352])^(a[232] & b[353])^(a[231] & b[354])^(a[230] & b[355])^(a[229] & b[356])^(a[228] & b[357])^(a[227] & b[358])^(a[226] & b[359])^(a[225] & b[360])^(a[224] & b[361])^(a[223] & b[362])^(a[222] & b[363])^(a[221] & b[364])^(a[220] & b[365])^(a[219] & b[366])^(a[218] & b[367])^(a[217] & b[368])^(a[216] & b[369])^(a[215] & b[370])^(a[214] & b[371])^(a[213] & b[372])^(a[212] & b[373])^(a[211] & b[374])^(a[210] & b[375])^(a[209] & b[376])^(a[208] & b[377])^(a[207] & b[378])^(a[206] & b[379])^(a[205] & b[380])^(a[204] & b[381])^(a[203] & b[382])^(a[202] & b[383])^(a[201] & b[384])^(a[200] & b[385])^(a[199] & b[386])^(a[198] & b[387])^(a[197] & b[388])^(a[196] & b[389])^(a[195] & b[390])^(a[194] & b[391])^(a[193] & b[392])^(a[192] & b[393])^(a[191] & b[394])^(a[190] & b[395])^(a[189] & b[396])^(a[188] & b[397])^(a[187] & b[398])^(a[186] & b[399])^(a[185] & b[400])^(a[184] & b[401])^(a[183] & b[402])^(a[182] & b[403])^(a[181] & b[404])^(a[180] & b[405])^(a[179] & b[406])^(a[178] & b[407])^(a[177] & b[408]);
assign y[586] = (a[408] & b[178])^(a[407] & b[179])^(a[406] & b[180])^(a[405] & b[181])^(a[404] & b[182])^(a[403] & b[183])^(a[402] & b[184])^(a[401] & b[185])^(a[400] & b[186])^(a[399] & b[187])^(a[398] & b[188])^(a[397] & b[189])^(a[396] & b[190])^(a[395] & b[191])^(a[394] & b[192])^(a[393] & b[193])^(a[392] & b[194])^(a[391] & b[195])^(a[390] & b[196])^(a[389] & b[197])^(a[388] & b[198])^(a[387] & b[199])^(a[386] & b[200])^(a[385] & b[201])^(a[384] & b[202])^(a[383] & b[203])^(a[382] & b[204])^(a[381] & b[205])^(a[380] & b[206])^(a[379] & b[207])^(a[378] & b[208])^(a[377] & b[209])^(a[376] & b[210])^(a[375] & b[211])^(a[374] & b[212])^(a[373] & b[213])^(a[372] & b[214])^(a[371] & b[215])^(a[370] & b[216])^(a[369] & b[217])^(a[368] & b[218])^(a[367] & b[219])^(a[366] & b[220])^(a[365] & b[221])^(a[364] & b[222])^(a[363] & b[223])^(a[362] & b[224])^(a[361] & b[225])^(a[360] & b[226])^(a[359] & b[227])^(a[358] & b[228])^(a[357] & b[229])^(a[356] & b[230])^(a[355] & b[231])^(a[354] & b[232])^(a[353] & b[233])^(a[352] & b[234])^(a[351] & b[235])^(a[350] & b[236])^(a[349] & b[237])^(a[348] & b[238])^(a[347] & b[239])^(a[346] & b[240])^(a[345] & b[241])^(a[344] & b[242])^(a[343] & b[243])^(a[342] & b[244])^(a[341] & b[245])^(a[340] & b[246])^(a[339] & b[247])^(a[338] & b[248])^(a[337] & b[249])^(a[336] & b[250])^(a[335] & b[251])^(a[334] & b[252])^(a[333] & b[253])^(a[332] & b[254])^(a[331] & b[255])^(a[330] & b[256])^(a[329] & b[257])^(a[328] & b[258])^(a[327] & b[259])^(a[326] & b[260])^(a[325] & b[261])^(a[324] & b[262])^(a[323] & b[263])^(a[322] & b[264])^(a[321] & b[265])^(a[320] & b[266])^(a[319] & b[267])^(a[318] & b[268])^(a[317] & b[269])^(a[316] & b[270])^(a[315] & b[271])^(a[314] & b[272])^(a[313] & b[273])^(a[312] & b[274])^(a[311] & b[275])^(a[310] & b[276])^(a[309] & b[277])^(a[308] & b[278])^(a[307] & b[279])^(a[306] & b[280])^(a[305] & b[281])^(a[304] & b[282])^(a[303] & b[283])^(a[302] & b[284])^(a[301] & b[285])^(a[300] & b[286])^(a[299] & b[287])^(a[298] & b[288])^(a[297] & b[289])^(a[296] & b[290])^(a[295] & b[291])^(a[294] & b[292])^(a[293] & b[293])^(a[292] & b[294])^(a[291] & b[295])^(a[290] & b[296])^(a[289] & b[297])^(a[288] & b[298])^(a[287] & b[299])^(a[286] & b[300])^(a[285] & b[301])^(a[284] & b[302])^(a[283] & b[303])^(a[282] & b[304])^(a[281] & b[305])^(a[280] & b[306])^(a[279] & b[307])^(a[278] & b[308])^(a[277] & b[309])^(a[276] & b[310])^(a[275] & b[311])^(a[274] & b[312])^(a[273] & b[313])^(a[272] & b[314])^(a[271] & b[315])^(a[270] & b[316])^(a[269] & b[317])^(a[268] & b[318])^(a[267] & b[319])^(a[266] & b[320])^(a[265] & b[321])^(a[264] & b[322])^(a[263] & b[323])^(a[262] & b[324])^(a[261] & b[325])^(a[260] & b[326])^(a[259] & b[327])^(a[258] & b[328])^(a[257] & b[329])^(a[256] & b[330])^(a[255] & b[331])^(a[254] & b[332])^(a[253] & b[333])^(a[252] & b[334])^(a[251] & b[335])^(a[250] & b[336])^(a[249] & b[337])^(a[248] & b[338])^(a[247] & b[339])^(a[246] & b[340])^(a[245] & b[341])^(a[244] & b[342])^(a[243] & b[343])^(a[242] & b[344])^(a[241] & b[345])^(a[240] & b[346])^(a[239] & b[347])^(a[238] & b[348])^(a[237] & b[349])^(a[236] & b[350])^(a[235] & b[351])^(a[234] & b[352])^(a[233] & b[353])^(a[232] & b[354])^(a[231] & b[355])^(a[230] & b[356])^(a[229] & b[357])^(a[228] & b[358])^(a[227] & b[359])^(a[226] & b[360])^(a[225] & b[361])^(a[224] & b[362])^(a[223] & b[363])^(a[222] & b[364])^(a[221] & b[365])^(a[220] & b[366])^(a[219] & b[367])^(a[218] & b[368])^(a[217] & b[369])^(a[216] & b[370])^(a[215] & b[371])^(a[214] & b[372])^(a[213] & b[373])^(a[212] & b[374])^(a[211] & b[375])^(a[210] & b[376])^(a[209] & b[377])^(a[208] & b[378])^(a[207] & b[379])^(a[206] & b[380])^(a[205] & b[381])^(a[204] & b[382])^(a[203] & b[383])^(a[202] & b[384])^(a[201] & b[385])^(a[200] & b[386])^(a[199] & b[387])^(a[198] & b[388])^(a[197] & b[389])^(a[196] & b[390])^(a[195] & b[391])^(a[194] & b[392])^(a[193] & b[393])^(a[192] & b[394])^(a[191] & b[395])^(a[190] & b[396])^(a[189] & b[397])^(a[188] & b[398])^(a[187] & b[399])^(a[186] & b[400])^(a[185] & b[401])^(a[184] & b[402])^(a[183] & b[403])^(a[182] & b[404])^(a[181] & b[405])^(a[180] & b[406])^(a[179] & b[407])^(a[178] & b[408]);
assign y[587] = (a[408] & b[179])^(a[407] & b[180])^(a[406] & b[181])^(a[405] & b[182])^(a[404] & b[183])^(a[403] & b[184])^(a[402] & b[185])^(a[401] & b[186])^(a[400] & b[187])^(a[399] & b[188])^(a[398] & b[189])^(a[397] & b[190])^(a[396] & b[191])^(a[395] & b[192])^(a[394] & b[193])^(a[393] & b[194])^(a[392] & b[195])^(a[391] & b[196])^(a[390] & b[197])^(a[389] & b[198])^(a[388] & b[199])^(a[387] & b[200])^(a[386] & b[201])^(a[385] & b[202])^(a[384] & b[203])^(a[383] & b[204])^(a[382] & b[205])^(a[381] & b[206])^(a[380] & b[207])^(a[379] & b[208])^(a[378] & b[209])^(a[377] & b[210])^(a[376] & b[211])^(a[375] & b[212])^(a[374] & b[213])^(a[373] & b[214])^(a[372] & b[215])^(a[371] & b[216])^(a[370] & b[217])^(a[369] & b[218])^(a[368] & b[219])^(a[367] & b[220])^(a[366] & b[221])^(a[365] & b[222])^(a[364] & b[223])^(a[363] & b[224])^(a[362] & b[225])^(a[361] & b[226])^(a[360] & b[227])^(a[359] & b[228])^(a[358] & b[229])^(a[357] & b[230])^(a[356] & b[231])^(a[355] & b[232])^(a[354] & b[233])^(a[353] & b[234])^(a[352] & b[235])^(a[351] & b[236])^(a[350] & b[237])^(a[349] & b[238])^(a[348] & b[239])^(a[347] & b[240])^(a[346] & b[241])^(a[345] & b[242])^(a[344] & b[243])^(a[343] & b[244])^(a[342] & b[245])^(a[341] & b[246])^(a[340] & b[247])^(a[339] & b[248])^(a[338] & b[249])^(a[337] & b[250])^(a[336] & b[251])^(a[335] & b[252])^(a[334] & b[253])^(a[333] & b[254])^(a[332] & b[255])^(a[331] & b[256])^(a[330] & b[257])^(a[329] & b[258])^(a[328] & b[259])^(a[327] & b[260])^(a[326] & b[261])^(a[325] & b[262])^(a[324] & b[263])^(a[323] & b[264])^(a[322] & b[265])^(a[321] & b[266])^(a[320] & b[267])^(a[319] & b[268])^(a[318] & b[269])^(a[317] & b[270])^(a[316] & b[271])^(a[315] & b[272])^(a[314] & b[273])^(a[313] & b[274])^(a[312] & b[275])^(a[311] & b[276])^(a[310] & b[277])^(a[309] & b[278])^(a[308] & b[279])^(a[307] & b[280])^(a[306] & b[281])^(a[305] & b[282])^(a[304] & b[283])^(a[303] & b[284])^(a[302] & b[285])^(a[301] & b[286])^(a[300] & b[287])^(a[299] & b[288])^(a[298] & b[289])^(a[297] & b[290])^(a[296] & b[291])^(a[295] & b[292])^(a[294] & b[293])^(a[293] & b[294])^(a[292] & b[295])^(a[291] & b[296])^(a[290] & b[297])^(a[289] & b[298])^(a[288] & b[299])^(a[287] & b[300])^(a[286] & b[301])^(a[285] & b[302])^(a[284] & b[303])^(a[283] & b[304])^(a[282] & b[305])^(a[281] & b[306])^(a[280] & b[307])^(a[279] & b[308])^(a[278] & b[309])^(a[277] & b[310])^(a[276] & b[311])^(a[275] & b[312])^(a[274] & b[313])^(a[273] & b[314])^(a[272] & b[315])^(a[271] & b[316])^(a[270] & b[317])^(a[269] & b[318])^(a[268] & b[319])^(a[267] & b[320])^(a[266] & b[321])^(a[265] & b[322])^(a[264] & b[323])^(a[263] & b[324])^(a[262] & b[325])^(a[261] & b[326])^(a[260] & b[327])^(a[259] & b[328])^(a[258] & b[329])^(a[257] & b[330])^(a[256] & b[331])^(a[255] & b[332])^(a[254] & b[333])^(a[253] & b[334])^(a[252] & b[335])^(a[251] & b[336])^(a[250] & b[337])^(a[249] & b[338])^(a[248] & b[339])^(a[247] & b[340])^(a[246] & b[341])^(a[245] & b[342])^(a[244] & b[343])^(a[243] & b[344])^(a[242] & b[345])^(a[241] & b[346])^(a[240] & b[347])^(a[239] & b[348])^(a[238] & b[349])^(a[237] & b[350])^(a[236] & b[351])^(a[235] & b[352])^(a[234] & b[353])^(a[233] & b[354])^(a[232] & b[355])^(a[231] & b[356])^(a[230] & b[357])^(a[229] & b[358])^(a[228] & b[359])^(a[227] & b[360])^(a[226] & b[361])^(a[225] & b[362])^(a[224] & b[363])^(a[223] & b[364])^(a[222] & b[365])^(a[221] & b[366])^(a[220] & b[367])^(a[219] & b[368])^(a[218] & b[369])^(a[217] & b[370])^(a[216] & b[371])^(a[215] & b[372])^(a[214] & b[373])^(a[213] & b[374])^(a[212] & b[375])^(a[211] & b[376])^(a[210] & b[377])^(a[209] & b[378])^(a[208] & b[379])^(a[207] & b[380])^(a[206] & b[381])^(a[205] & b[382])^(a[204] & b[383])^(a[203] & b[384])^(a[202] & b[385])^(a[201] & b[386])^(a[200] & b[387])^(a[199] & b[388])^(a[198] & b[389])^(a[197] & b[390])^(a[196] & b[391])^(a[195] & b[392])^(a[194] & b[393])^(a[193] & b[394])^(a[192] & b[395])^(a[191] & b[396])^(a[190] & b[397])^(a[189] & b[398])^(a[188] & b[399])^(a[187] & b[400])^(a[186] & b[401])^(a[185] & b[402])^(a[184] & b[403])^(a[183] & b[404])^(a[182] & b[405])^(a[181] & b[406])^(a[180] & b[407])^(a[179] & b[408]);
assign y[588] = (a[408] & b[180])^(a[407] & b[181])^(a[406] & b[182])^(a[405] & b[183])^(a[404] & b[184])^(a[403] & b[185])^(a[402] & b[186])^(a[401] & b[187])^(a[400] & b[188])^(a[399] & b[189])^(a[398] & b[190])^(a[397] & b[191])^(a[396] & b[192])^(a[395] & b[193])^(a[394] & b[194])^(a[393] & b[195])^(a[392] & b[196])^(a[391] & b[197])^(a[390] & b[198])^(a[389] & b[199])^(a[388] & b[200])^(a[387] & b[201])^(a[386] & b[202])^(a[385] & b[203])^(a[384] & b[204])^(a[383] & b[205])^(a[382] & b[206])^(a[381] & b[207])^(a[380] & b[208])^(a[379] & b[209])^(a[378] & b[210])^(a[377] & b[211])^(a[376] & b[212])^(a[375] & b[213])^(a[374] & b[214])^(a[373] & b[215])^(a[372] & b[216])^(a[371] & b[217])^(a[370] & b[218])^(a[369] & b[219])^(a[368] & b[220])^(a[367] & b[221])^(a[366] & b[222])^(a[365] & b[223])^(a[364] & b[224])^(a[363] & b[225])^(a[362] & b[226])^(a[361] & b[227])^(a[360] & b[228])^(a[359] & b[229])^(a[358] & b[230])^(a[357] & b[231])^(a[356] & b[232])^(a[355] & b[233])^(a[354] & b[234])^(a[353] & b[235])^(a[352] & b[236])^(a[351] & b[237])^(a[350] & b[238])^(a[349] & b[239])^(a[348] & b[240])^(a[347] & b[241])^(a[346] & b[242])^(a[345] & b[243])^(a[344] & b[244])^(a[343] & b[245])^(a[342] & b[246])^(a[341] & b[247])^(a[340] & b[248])^(a[339] & b[249])^(a[338] & b[250])^(a[337] & b[251])^(a[336] & b[252])^(a[335] & b[253])^(a[334] & b[254])^(a[333] & b[255])^(a[332] & b[256])^(a[331] & b[257])^(a[330] & b[258])^(a[329] & b[259])^(a[328] & b[260])^(a[327] & b[261])^(a[326] & b[262])^(a[325] & b[263])^(a[324] & b[264])^(a[323] & b[265])^(a[322] & b[266])^(a[321] & b[267])^(a[320] & b[268])^(a[319] & b[269])^(a[318] & b[270])^(a[317] & b[271])^(a[316] & b[272])^(a[315] & b[273])^(a[314] & b[274])^(a[313] & b[275])^(a[312] & b[276])^(a[311] & b[277])^(a[310] & b[278])^(a[309] & b[279])^(a[308] & b[280])^(a[307] & b[281])^(a[306] & b[282])^(a[305] & b[283])^(a[304] & b[284])^(a[303] & b[285])^(a[302] & b[286])^(a[301] & b[287])^(a[300] & b[288])^(a[299] & b[289])^(a[298] & b[290])^(a[297] & b[291])^(a[296] & b[292])^(a[295] & b[293])^(a[294] & b[294])^(a[293] & b[295])^(a[292] & b[296])^(a[291] & b[297])^(a[290] & b[298])^(a[289] & b[299])^(a[288] & b[300])^(a[287] & b[301])^(a[286] & b[302])^(a[285] & b[303])^(a[284] & b[304])^(a[283] & b[305])^(a[282] & b[306])^(a[281] & b[307])^(a[280] & b[308])^(a[279] & b[309])^(a[278] & b[310])^(a[277] & b[311])^(a[276] & b[312])^(a[275] & b[313])^(a[274] & b[314])^(a[273] & b[315])^(a[272] & b[316])^(a[271] & b[317])^(a[270] & b[318])^(a[269] & b[319])^(a[268] & b[320])^(a[267] & b[321])^(a[266] & b[322])^(a[265] & b[323])^(a[264] & b[324])^(a[263] & b[325])^(a[262] & b[326])^(a[261] & b[327])^(a[260] & b[328])^(a[259] & b[329])^(a[258] & b[330])^(a[257] & b[331])^(a[256] & b[332])^(a[255] & b[333])^(a[254] & b[334])^(a[253] & b[335])^(a[252] & b[336])^(a[251] & b[337])^(a[250] & b[338])^(a[249] & b[339])^(a[248] & b[340])^(a[247] & b[341])^(a[246] & b[342])^(a[245] & b[343])^(a[244] & b[344])^(a[243] & b[345])^(a[242] & b[346])^(a[241] & b[347])^(a[240] & b[348])^(a[239] & b[349])^(a[238] & b[350])^(a[237] & b[351])^(a[236] & b[352])^(a[235] & b[353])^(a[234] & b[354])^(a[233] & b[355])^(a[232] & b[356])^(a[231] & b[357])^(a[230] & b[358])^(a[229] & b[359])^(a[228] & b[360])^(a[227] & b[361])^(a[226] & b[362])^(a[225] & b[363])^(a[224] & b[364])^(a[223] & b[365])^(a[222] & b[366])^(a[221] & b[367])^(a[220] & b[368])^(a[219] & b[369])^(a[218] & b[370])^(a[217] & b[371])^(a[216] & b[372])^(a[215] & b[373])^(a[214] & b[374])^(a[213] & b[375])^(a[212] & b[376])^(a[211] & b[377])^(a[210] & b[378])^(a[209] & b[379])^(a[208] & b[380])^(a[207] & b[381])^(a[206] & b[382])^(a[205] & b[383])^(a[204] & b[384])^(a[203] & b[385])^(a[202] & b[386])^(a[201] & b[387])^(a[200] & b[388])^(a[199] & b[389])^(a[198] & b[390])^(a[197] & b[391])^(a[196] & b[392])^(a[195] & b[393])^(a[194] & b[394])^(a[193] & b[395])^(a[192] & b[396])^(a[191] & b[397])^(a[190] & b[398])^(a[189] & b[399])^(a[188] & b[400])^(a[187] & b[401])^(a[186] & b[402])^(a[185] & b[403])^(a[184] & b[404])^(a[183] & b[405])^(a[182] & b[406])^(a[181] & b[407])^(a[180] & b[408]);
assign y[589] = (a[408] & b[181])^(a[407] & b[182])^(a[406] & b[183])^(a[405] & b[184])^(a[404] & b[185])^(a[403] & b[186])^(a[402] & b[187])^(a[401] & b[188])^(a[400] & b[189])^(a[399] & b[190])^(a[398] & b[191])^(a[397] & b[192])^(a[396] & b[193])^(a[395] & b[194])^(a[394] & b[195])^(a[393] & b[196])^(a[392] & b[197])^(a[391] & b[198])^(a[390] & b[199])^(a[389] & b[200])^(a[388] & b[201])^(a[387] & b[202])^(a[386] & b[203])^(a[385] & b[204])^(a[384] & b[205])^(a[383] & b[206])^(a[382] & b[207])^(a[381] & b[208])^(a[380] & b[209])^(a[379] & b[210])^(a[378] & b[211])^(a[377] & b[212])^(a[376] & b[213])^(a[375] & b[214])^(a[374] & b[215])^(a[373] & b[216])^(a[372] & b[217])^(a[371] & b[218])^(a[370] & b[219])^(a[369] & b[220])^(a[368] & b[221])^(a[367] & b[222])^(a[366] & b[223])^(a[365] & b[224])^(a[364] & b[225])^(a[363] & b[226])^(a[362] & b[227])^(a[361] & b[228])^(a[360] & b[229])^(a[359] & b[230])^(a[358] & b[231])^(a[357] & b[232])^(a[356] & b[233])^(a[355] & b[234])^(a[354] & b[235])^(a[353] & b[236])^(a[352] & b[237])^(a[351] & b[238])^(a[350] & b[239])^(a[349] & b[240])^(a[348] & b[241])^(a[347] & b[242])^(a[346] & b[243])^(a[345] & b[244])^(a[344] & b[245])^(a[343] & b[246])^(a[342] & b[247])^(a[341] & b[248])^(a[340] & b[249])^(a[339] & b[250])^(a[338] & b[251])^(a[337] & b[252])^(a[336] & b[253])^(a[335] & b[254])^(a[334] & b[255])^(a[333] & b[256])^(a[332] & b[257])^(a[331] & b[258])^(a[330] & b[259])^(a[329] & b[260])^(a[328] & b[261])^(a[327] & b[262])^(a[326] & b[263])^(a[325] & b[264])^(a[324] & b[265])^(a[323] & b[266])^(a[322] & b[267])^(a[321] & b[268])^(a[320] & b[269])^(a[319] & b[270])^(a[318] & b[271])^(a[317] & b[272])^(a[316] & b[273])^(a[315] & b[274])^(a[314] & b[275])^(a[313] & b[276])^(a[312] & b[277])^(a[311] & b[278])^(a[310] & b[279])^(a[309] & b[280])^(a[308] & b[281])^(a[307] & b[282])^(a[306] & b[283])^(a[305] & b[284])^(a[304] & b[285])^(a[303] & b[286])^(a[302] & b[287])^(a[301] & b[288])^(a[300] & b[289])^(a[299] & b[290])^(a[298] & b[291])^(a[297] & b[292])^(a[296] & b[293])^(a[295] & b[294])^(a[294] & b[295])^(a[293] & b[296])^(a[292] & b[297])^(a[291] & b[298])^(a[290] & b[299])^(a[289] & b[300])^(a[288] & b[301])^(a[287] & b[302])^(a[286] & b[303])^(a[285] & b[304])^(a[284] & b[305])^(a[283] & b[306])^(a[282] & b[307])^(a[281] & b[308])^(a[280] & b[309])^(a[279] & b[310])^(a[278] & b[311])^(a[277] & b[312])^(a[276] & b[313])^(a[275] & b[314])^(a[274] & b[315])^(a[273] & b[316])^(a[272] & b[317])^(a[271] & b[318])^(a[270] & b[319])^(a[269] & b[320])^(a[268] & b[321])^(a[267] & b[322])^(a[266] & b[323])^(a[265] & b[324])^(a[264] & b[325])^(a[263] & b[326])^(a[262] & b[327])^(a[261] & b[328])^(a[260] & b[329])^(a[259] & b[330])^(a[258] & b[331])^(a[257] & b[332])^(a[256] & b[333])^(a[255] & b[334])^(a[254] & b[335])^(a[253] & b[336])^(a[252] & b[337])^(a[251] & b[338])^(a[250] & b[339])^(a[249] & b[340])^(a[248] & b[341])^(a[247] & b[342])^(a[246] & b[343])^(a[245] & b[344])^(a[244] & b[345])^(a[243] & b[346])^(a[242] & b[347])^(a[241] & b[348])^(a[240] & b[349])^(a[239] & b[350])^(a[238] & b[351])^(a[237] & b[352])^(a[236] & b[353])^(a[235] & b[354])^(a[234] & b[355])^(a[233] & b[356])^(a[232] & b[357])^(a[231] & b[358])^(a[230] & b[359])^(a[229] & b[360])^(a[228] & b[361])^(a[227] & b[362])^(a[226] & b[363])^(a[225] & b[364])^(a[224] & b[365])^(a[223] & b[366])^(a[222] & b[367])^(a[221] & b[368])^(a[220] & b[369])^(a[219] & b[370])^(a[218] & b[371])^(a[217] & b[372])^(a[216] & b[373])^(a[215] & b[374])^(a[214] & b[375])^(a[213] & b[376])^(a[212] & b[377])^(a[211] & b[378])^(a[210] & b[379])^(a[209] & b[380])^(a[208] & b[381])^(a[207] & b[382])^(a[206] & b[383])^(a[205] & b[384])^(a[204] & b[385])^(a[203] & b[386])^(a[202] & b[387])^(a[201] & b[388])^(a[200] & b[389])^(a[199] & b[390])^(a[198] & b[391])^(a[197] & b[392])^(a[196] & b[393])^(a[195] & b[394])^(a[194] & b[395])^(a[193] & b[396])^(a[192] & b[397])^(a[191] & b[398])^(a[190] & b[399])^(a[189] & b[400])^(a[188] & b[401])^(a[187] & b[402])^(a[186] & b[403])^(a[185] & b[404])^(a[184] & b[405])^(a[183] & b[406])^(a[182] & b[407])^(a[181] & b[408]);
assign y[590] = (a[408] & b[182])^(a[407] & b[183])^(a[406] & b[184])^(a[405] & b[185])^(a[404] & b[186])^(a[403] & b[187])^(a[402] & b[188])^(a[401] & b[189])^(a[400] & b[190])^(a[399] & b[191])^(a[398] & b[192])^(a[397] & b[193])^(a[396] & b[194])^(a[395] & b[195])^(a[394] & b[196])^(a[393] & b[197])^(a[392] & b[198])^(a[391] & b[199])^(a[390] & b[200])^(a[389] & b[201])^(a[388] & b[202])^(a[387] & b[203])^(a[386] & b[204])^(a[385] & b[205])^(a[384] & b[206])^(a[383] & b[207])^(a[382] & b[208])^(a[381] & b[209])^(a[380] & b[210])^(a[379] & b[211])^(a[378] & b[212])^(a[377] & b[213])^(a[376] & b[214])^(a[375] & b[215])^(a[374] & b[216])^(a[373] & b[217])^(a[372] & b[218])^(a[371] & b[219])^(a[370] & b[220])^(a[369] & b[221])^(a[368] & b[222])^(a[367] & b[223])^(a[366] & b[224])^(a[365] & b[225])^(a[364] & b[226])^(a[363] & b[227])^(a[362] & b[228])^(a[361] & b[229])^(a[360] & b[230])^(a[359] & b[231])^(a[358] & b[232])^(a[357] & b[233])^(a[356] & b[234])^(a[355] & b[235])^(a[354] & b[236])^(a[353] & b[237])^(a[352] & b[238])^(a[351] & b[239])^(a[350] & b[240])^(a[349] & b[241])^(a[348] & b[242])^(a[347] & b[243])^(a[346] & b[244])^(a[345] & b[245])^(a[344] & b[246])^(a[343] & b[247])^(a[342] & b[248])^(a[341] & b[249])^(a[340] & b[250])^(a[339] & b[251])^(a[338] & b[252])^(a[337] & b[253])^(a[336] & b[254])^(a[335] & b[255])^(a[334] & b[256])^(a[333] & b[257])^(a[332] & b[258])^(a[331] & b[259])^(a[330] & b[260])^(a[329] & b[261])^(a[328] & b[262])^(a[327] & b[263])^(a[326] & b[264])^(a[325] & b[265])^(a[324] & b[266])^(a[323] & b[267])^(a[322] & b[268])^(a[321] & b[269])^(a[320] & b[270])^(a[319] & b[271])^(a[318] & b[272])^(a[317] & b[273])^(a[316] & b[274])^(a[315] & b[275])^(a[314] & b[276])^(a[313] & b[277])^(a[312] & b[278])^(a[311] & b[279])^(a[310] & b[280])^(a[309] & b[281])^(a[308] & b[282])^(a[307] & b[283])^(a[306] & b[284])^(a[305] & b[285])^(a[304] & b[286])^(a[303] & b[287])^(a[302] & b[288])^(a[301] & b[289])^(a[300] & b[290])^(a[299] & b[291])^(a[298] & b[292])^(a[297] & b[293])^(a[296] & b[294])^(a[295] & b[295])^(a[294] & b[296])^(a[293] & b[297])^(a[292] & b[298])^(a[291] & b[299])^(a[290] & b[300])^(a[289] & b[301])^(a[288] & b[302])^(a[287] & b[303])^(a[286] & b[304])^(a[285] & b[305])^(a[284] & b[306])^(a[283] & b[307])^(a[282] & b[308])^(a[281] & b[309])^(a[280] & b[310])^(a[279] & b[311])^(a[278] & b[312])^(a[277] & b[313])^(a[276] & b[314])^(a[275] & b[315])^(a[274] & b[316])^(a[273] & b[317])^(a[272] & b[318])^(a[271] & b[319])^(a[270] & b[320])^(a[269] & b[321])^(a[268] & b[322])^(a[267] & b[323])^(a[266] & b[324])^(a[265] & b[325])^(a[264] & b[326])^(a[263] & b[327])^(a[262] & b[328])^(a[261] & b[329])^(a[260] & b[330])^(a[259] & b[331])^(a[258] & b[332])^(a[257] & b[333])^(a[256] & b[334])^(a[255] & b[335])^(a[254] & b[336])^(a[253] & b[337])^(a[252] & b[338])^(a[251] & b[339])^(a[250] & b[340])^(a[249] & b[341])^(a[248] & b[342])^(a[247] & b[343])^(a[246] & b[344])^(a[245] & b[345])^(a[244] & b[346])^(a[243] & b[347])^(a[242] & b[348])^(a[241] & b[349])^(a[240] & b[350])^(a[239] & b[351])^(a[238] & b[352])^(a[237] & b[353])^(a[236] & b[354])^(a[235] & b[355])^(a[234] & b[356])^(a[233] & b[357])^(a[232] & b[358])^(a[231] & b[359])^(a[230] & b[360])^(a[229] & b[361])^(a[228] & b[362])^(a[227] & b[363])^(a[226] & b[364])^(a[225] & b[365])^(a[224] & b[366])^(a[223] & b[367])^(a[222] & b[368])^(a[221] & b[369])^(a[220] & b[370])^(a[219] & b[371])^(a[218] & b[372])^(a[217] & b[373])^(a[216] & b[374])^(a[215] & b[375])^(a[214] & b[376])^(a[213] & b[377])^(a[212] & b[378])^(a[211] & b[379])^(a[210] & b[380])^(a[209] & b[381])^(a[208] & b[382])^(a[207] & b[383])^(a[206] & b[384])^(a[205] & b[385])^(a[204] & b[386])^(a[203] & b[387])^(a[202] & b[388])^(a[201] & b[389])^(a[200] & b[390])^(a[199] & b[391])^(a[198] & b[392])^(a[197] & b[393])^(a[196] & b[394])^(a[195] & b[395])^(a[194] & b[396])^(a[193] & b[397])^(a[192] & b[398])^(a[191] & b[399])^(a[190] & b[400])^(a[189] & b[401])^(a[188] & b[402])^(a[187] & b[403])^(a[186] & b[404])^(a[185] & b[405])^(a[184] & b[406])^(a[183] & b[407])^(a[182] & b[408]);
assign y[591] = (a[408] & b[183])^(a[407] & b[184])^(a[406] & b[185])^(a[405] & b[186])^(a[404] & b[187])^(a[403] & b[188])^(a[402] & b[189])^(a[401] & b[190])^(a[400] & b[191])^(a[399] & b[192])^(a[398] & b[193])^(a[397] & b[194])^(a[396] & b[195])^(a[395] & b[196])^(a[394] & b[197])^(a[393] & b[198])^(a[392] & b[199])^(a[391] & b[200])^(a[390] & b[201])^(a[389] & b[202])^(a[388] & b[203])^(a[387] & b[204])^(a[386] & b[205])^(a[385] & b[206])^(a[384] & b[207])^(a[383] & b[208])^(a[382] & b[209])^(a[381] & b[210])^(a[380] & b[211])^(a[379] & b[212])^(a[378] & b[213])^(a[377] & b[214])^(a[376] & b[215])^(a[375] & b[216])^(a[374] & b[217])^(a[373] & b[218])^(a[372] & b[219])^(a[371] & b[220])^(a[370] & b[221])^(a[369] & b[222])^(a[368] & b[223])^(a[367] & b[224])^(a[366] & b[225])^(a[365] & b[226])^(a[364] & b[227])^(a[363] & b[228])^(a[362] & b[229])^(a[361] & b[230])^(a[360] & b[231])^(a[359] & b[232])^(a[358] & b[233])^(a[357] & b[234])^(a[356] & b[235])^(a[355] & b[236])^(a[354] & b[237])^(a[353] & b[238])^(a[352] & b[239])^(a[351] & b[240])^(a[350] & b[241])^(a[349] & b[242])^(a[348] & b[243])^(a[347] & b[244])^(a[346] & b[245])^(a[345] & b[246])^(a[344] & b[247])^(a[343] & b[248])^(a[342] & b[249])^(a[341] & b[250])^(a[340] & b[251])^(a[339] & b[252])^(a[338] & b[253])^(a[337] & b[254])^(a[336] & b[255])^(a[335] & b[256])^(a[334] & b[257])^(a[333] & b[258])^(a[332] & b[259])^(a[331] & b[260])^(a[330] & b[261])^(a[329] & b[262])^(a[328] & b[263])^(a[327] & b[264])^(a[326] & b[265])^(a[325] & b[266])^(a[324] & b[267])^(a[323] & b[268])^(a[322] & b[269])^(a[321] & b[270])^(a[320] & b[271])^(a[319] & b[272])^(a[318] & b[273])^(a[317] & b[274])^(a[316] & b[275])^(a[315] & b[276])^(a[314] & b[277])^(a[313] & b[278])^(a[312] & b[279])^(a[311] & b[280])^(a[310] & b[281])^(a[309] & b[282])^(a[308] & b[283])^(a[307] & b[284])^(a[306] & b[285])^(a[305] & b[286])^(a[304] & b[287])^(a[303] & b[288])^(a[302] & b[289])^(a[301] & b[290])^(a[300] & b[291])^(a[299] & b[292])^(a[298] & b[293])^(a[297] & b[294])^(a[296] & b[295])^(a[295] & b[296])^(a[294] & b[297])^(a[293] & b[298])^(a[292] & b[299])^(a[291] & b[300])^(a[290] & b[301])^(a[289] & b[302])^(a[288] & b[303])^(a[287] & b[304])^(a[286] & b[305])^(a[285] & b[306])^(a[284] & b[307])^(a[283] & b[308])^(a[282] & b[309])^(a[281] & b[310])^(a[280] & b[311])^(a[279] & b[312])^(a[278] & b[313])^(a[277] & b[314])^(a[276] & b[315])^(a[275] & b[316])^(a[274] & b[317])^(a[273] & b[318])^(a[272] & b[319])^(a[271] & b[320])^(a[270] & b[321])^(a[269] & b[322])^(a[268] & b[323])^(a[267] & b[324])^(a[266] & b[325])^(a[265] & b[326])^(a[264] & b[327])^(a[263] & b[328])^(a[262] & b[329])^(a[261] & b[330])^(a[260] & b[331])^(a[259] & b[332])^(a[258] & b[333])^(a[257] & b[334])^(a[256] & b[335])^(a[255] & b[336])^(a[254] & b[337])^(a[253] & b[338])^(a[252] & b[339])^(a[251] & b[340])^(a[250] & b[341])^(a[249] & b[342])^(a[248] & b[343])^(a[247] & b[344])^(a[246] & b[345])^(a[245] & b[346])^(a[244] & b[347])^(a[243] & b[348])^(a[242] & b[349])^(a[241] & b[350])^(a[240] & b[351])^(a[239] & b[352])^(a[238] & b[353])^(a[237] & b[354])^(a[236] & b[355])^(a[235] & b[356])^(a[234] & b[357])^(a[233] & b[358])^(a[232] & b[359])^(a[231] & b[360])^(a[230] & b[361])^(a[229] & b[362])^(a[228] & b[363])^(a[227] & b[364])^(a[226] & b[365])^(a[225] & b[366])^(a[224] & b[367])^(a[223] & b[368])^(a[222] & b[369])^(a[221] & b[370])^(a[220] & b[371])^(a[219] & b[372])^(a[218] & b[373])^(a[217] & b[374])^(a[216] & b[375])^(a[215] & b[376])^(a[214] & b[377])^(a[213] & b[378])^(a[212] & b[379])^(a[211] & b[380])^(a[210] & b[381])^(a[209] & b[382])^(a[208] & b[383])^(a[207] & b[384])^(a[206] & b[385])^(a[205] & b[386])^(a[204] & b[387])^(a[203] & b[388])^(a[202] & b[389])^(a[201] & b[390])^(a[200] & b[391])^(a[199] & b[392])^(a[198] & b[393])^(a[197] & b[394])^(a[196] & b[395])^(a[195] & b[396])^(a[194] & b[397])^(a[193] & b[398])^(a[192] & b[399])^(a[191] & b[400])^(a[190] & b[401])^(a[189] & b[402])^(a[188] & b[403])^(a[187] & b[404])^(a[186] & b[405])^(a[185] & b[406])^(a[184] & b[407])^(a[183] & b[408]);
assign y[592] = (a[408] & b[184])^(a[407] & b[185])^(a[406] & b[186])^(a[405] & b[187])^(a[404] & b[188])^(a[403] & b[189])^(a[402] & b[190])^(a[401] & b[191])^(a[400] & b[192])^(a[399] & b[193])^(a[398] & b[194])^(a[397] & b[195])^(a[396] & b[196])^(a[395] & b[197])^(a[394] & b[198])^(a[393] & b[199])^(a[392] & b[200])^(a[391] & b[201])^(a[390] & b[202])^(a[389] & b[203])^(a[388] & b[204])^(a[387] & b[205])^(a[386] & b[206])^(a[385] & b[207])^(a[384] & b[208])^(a[383] & b[209])^(a[382] & b[210])^(a[381] & b[211])^(a[380] & b[212])^(a[379] & b[213])^(a[378] & b[214])^(a[377] & b[215])^(a[376] & b[216])^(a[375] & b[217])^(a[374] & b[218])^(a[373] & b[219])^(a[372] & b[220])^(a[371] & b[221])^(a[370] & b[222])^(a[369] & b[223])^(a[368] & b[224])^(a[367] & b[225])^(a[366] & b[226])^(a[365] & b[227])^(a[364] & b[228])^(a[363] & b[229])^(a[362] & b[230])^(a[361] & b[231])^(a[360] & b[232])^(a[359] & b[233])^(a[358] & b[234])^(a[357] & b[235])^(a[356] & b[236])^(a[355] & b[237])^(a[354] & b[238])^(a[353] & b[239])^(a[352] & b[240])^(a[351] & b[241])^(a[350] & b[242])^(a[349] & b[243])^(a[348] & b[244])^(a[347] & b[245])^(a[346] & b[246])^(a[345] & b[247])^(a[344] & b[248])^(a[343] & b[249])^(a[342] & b[250])^(a[341] & b[251])^(a[340] & b[252])^(a[339] & b[253])^(a[338] & b[254])^(a[337] & b[255])^(a[336] & b[256])^(a[335] & b[257])^(a[334] & b[258])^(a[333] & b[259])^(a[332] & b[260])^(a[331] & b[261])^(a[330] & b[262])^(a[329] & b[263])^(a[328] & b[264])^(a[327] & b[265])^(a[326] & b[266])^(a[325] & b[267])^(a[324] & b[268])^(a[323] & b[269])^(a[322] & b[270])^(a[321] & b[271])^(a[320] & b[272])^(a[319] & b[273])^(a[318] & b[274])^(a[317] & b[275])^(a[316] & b[276])^(a[315] & b[277])^(a[314] & b[278])^(a[313] & b[279])^(a[312] & b[280])^(a[311] & b[281])^(a[310] & b[282])^(a[309] & b[283])^(a[308] & b[284])^(a[307] & b[285])^(a[306] & b[286])^(a[305] & b[287])^(a[304] & b[288])^(a[303] & b[289])^(a[302] & b[290])^(a[301] & b[291])^(a[300] & b[292])^(a[299] & b[293])^(a[298] & b[294])^(a[297] & b[295])^(a[296] & b[296])^(a[295] & b[297])^(a[294] & b[298])^(a[293] & b[299])^(a[292] & b[300])^(a[291] & b[301])^(a[290] & b[302])^(a[289] & b[303])^(a[288] & b[304])^(a[287] & b[305])^(a[286] & b[306])^(a[285] & b[307])^(a[284] & b[308])^(a[283] & b[309])^(a[282] & b[310])^(a[281] & b[311])^(a[280] & b[312])^(a[279] & b[313])^(a[278] & b[314])^(a[277] & b[315])^(a[276] & b[316])^(a[275] & b[317])^(a[274] & b[318])^(a[273] & b[319])^(a[272] & b[320])^(a[271] & b[321])^(a[270] & b[322])^(a[269] & b[323])^(a[268] & b[324])^(a[267] & b[325])^(a[266] & b[326])^(a[265] & b[327])^(a[264] & b[328])^(a[263] & b[329])^(a[262] & b[330])^(a[261] & b[331])^(a[260] & b[332])^(a[259] & b[333])^(a[258] & b[334])^(a[257] & b[335])^(a[256] & b[336])^(a[255] & b[337])^(a[254] & b[338])^(a[253] & b[339])^(a[252] & b[340])^(a[251] & b[341])^(a[250] & b[342])^(a[249] & b[343])^(a[248] & b[344])^(a[247] & b[345])^(a[246] & b[346])^(a[245] & b[347])^(a[244] & b[348])^(a[243] & b[349])^(a[242] & b[350])^(a[241] & b[351])^(a[240] & b[352])^(a[239] & b[353])^(a[238] & b[354])^(a[237] & b[355])^(a[236] & b[356])^(a[235] & b[357])^(a[234] & b[358])^(a[233] & b[359])^(a[232] & b[360])^(a[231] & b[361])^(a[230] & b[362])^(a[229] & b[363])^(a[228] & b[364])^(a[227] & b[365])^(a[226] & b[366])^(a[225] & b[367])^(a[224] & b[368])^(a[223] & b[369])^(a[222] & b[370])^(a[221] & b[371])^(a[220] & b[372])^(a[219] & b[373])^(a[218] & b[374])^(a[217] & b[375])^(a[216] & b[376])^(a[215] & b[377])^(a[214] & b[378])^(a[213] & b[379])^(a[212] & b[380])^(a[211] & b[381])^(a[210] & b[382])^(a[209] & b[383])^(a[208] & b[384])^(a[207] & b[385])^(a[206] & b[386])^(a[205] & b[387])^(a[204] & b[388])^(a[203] & b[389])^(a[202] & b[390])^(a[201] & b[391])^(a[200] & b[392])^(a[199] & b[393])^(a[198] & b[394])^(a[197] & b[395])^(a[196] & b[396])^(a[195] & b[397])^(a[194] & b[398])^(a[193] & b[399])^(a[192] & b[400])^(a[191] & b[401])^(a[190] & b[402])^(a[189] & b[403])^(a[188] & b[404])^(a[187] & b[405])^(a[186] & b[406])^(a[185] & b[407])^(a[184] & b[408]);
assign y[593] = (a[408] & b[185])^(a[407] & b[186])^(a[406] & b[187])^(a[405] & b[188])^(a[404] & b[189])^(a[403] & b[190])^(a[402] & b[191])^(a[401] & b[192])^(a[400] & b[193])^(a[399] & b[194])^(a[398] & b[195])^(a[397] & b[196])^(a[396] & b[197])^(a[395] & b[198])^(a[394] & b[199])^(a[393] & b[200])^(a[392] & b[201])^(a[391] & b[202])^(a[390] & b[203])^(a[389] & b[204])^(a[388] & b[205])^(a[387] & b[206])^(a[386] & b[207])^(a[385] & b[208])^(a[384] & b[209])^(a[383] & b[210])^(a[382] & b[211])^(a[381] & b[212])^(a[380] & b[213])^(a[379] & b[214])^(a[378] & b[215])^(a[377] & b[216])^(a[376] & b[217])^(a[375] & b[218])^(a[374] & b[219])^(a[373] & b[220])^(a[372] & b[221])^(a[371] & b[222])^(a[370] & b[223])^(a[369] & b[224])^(a[368] & b[225])^(a[367] & b[226])^(a[366] & b[227])^(a[365] & b[228])^(a[364] & b[229])^(a[363] & b[230])^(a[362] & b[231])^(a[361] & b[232])^(a[360] & b[233])^(a[359] & b[234])^(a[358] & b[235])^(a[357] & b[236])^(a[356] & b[237])^(a[355] & b[238])^(a[354] & b[239])^(a[353] & b[240])^(a[352] & b[241])^(a[351] & b[242])^(a[350] & b[243])^(a[349] & b[244])^(a[348] & b[245])^(a[347] & b[246])^(a[346] & b[247])^(a[345] & b[248])^(a[344] & b[249])^(a[343] & b[250])^(a[342] & b[251])^(a[341] & b[252])^(a[340] & b[253])^(a[339] & b[254])^(a[338] & b[255])^(a[337] & b[256])^(a[336] & b[257])^(a[335] & b[258])^(a[334] & b[259])^(a[333] & b[260])^(a[332] & b[261])^(a[331] & b[262])^(a[330] & b[263])^(a[329] & b[264])^(a[328] & b[265])^(a[327] & b[266])^(a[326] & b[267])^(a[325] & b[268])^(a[324] & b[269])^(a[323] & b[270])^(a[322] & b[271])^(a[321] & b[272])^(a[320] & b[273])^(a[319] & b[274])^(a[318] & b[275])^(a[317] & b[276])^(a[316] & b[277])^(a[315] & b[278])^(a[314] & b[279])^(a[313] & b[280])^(a[312] & b[281])^(a[311] & b[282])^(a[310] & b[283])^(a[309] & b[284])^(a[308] & b[285])^(a[307] & b[286])^(a[306] & b[287])^(a[305] & b[288])^(a[304] & b[289])^(a[303] & b[290])^(a[302] & b[291])^(a[301] & b[292])^(a[300] & b[293])^(a[299] & b[294])^(a[298] & b[295])^(a[297] & b[296])^(a[296] & b[297])^(a[295] & b[298])^(a[294] & b[299])^(a[293] & b[300])^(a[292] & b[301])^(a[291] & b[302])^(a[290] & b[303])^(a[289] & b[304])^(a[288] & b[305])^(a[287] & b[306])^(a[286] & b[307])^(a[285] & b[308])^(a[284] & b[309])^(a[283] & b[310])^(a[282] & b[311])^(a[281] & b[312])^(a[280] & b[313])^(a[279] & b[314])^(a[278] & b[315])^(a[277] & b[316])^(a[276] & b[317])^(a[275] & b[318])^(a[274] & b[319])^(a[273] & b[320])^(a[272] & b[321])^(a[271] & b[322])^(a[270] & b[323])^(a[269] & b[324])^(a[268] & b[325])^(a[267] & b[326])^(a[266] & b[327])^(a[265] & b[328])^(a[264] & b[329])^(a[263] & b[330])^(a[262] & b[331])^(a[261] & b[332])^(a[260] & b[333])^(a[259] & b[334])^(a[258] & b[335])^(a[257] & b[336])^(a[256] & b[337])^(a[255] & b[338])^(a[254] & b[339])^(a[253] & b[340])^(a[252] & b[341])^(a[251] & b[342])^(a[250] & b[343])^(a[249] & b[344])^(a[248] & b[345])^(a[247] & b[346])^(a[246] & b[347])^(a[245] & b[348])^(a[244] & b[349])^(a[243] & b[350])^(a[242] & b[351])^(a[241] & b[352])^(a[240] & b[353])^(a[239] & b[354])^(a[238] & b[355])^(a[237] & b[356])^(a[236] & b[357])^(a[235] & b[358])^(a[234] & b[359])^(a[233] & b[360])^(a[232] & b[361])^(a[231] & b[362])^(a[230] & b[363])^(a[229] & b[364])^(a[228] & b[365])^(a[227] & b[366])^(a[226] & b[367])^(a[225] & b[368])^(a[224] & b[369])^(a[223] & b[370])^(a[222] & b[371])^(a[221] & b[372])^(a[220] & b[373])^(a[219] & b[374])^(a[218] & b[375])^(a[217] & b[376])^(a[216] & b[377])^(a[215] & b[378])^(a[214] & b[379])^(a[213] & b[380])^(a[212] & b[381])^(a[211] & b[382])^(a[210] & b[383])^(a[209] & b[384])^(a[208] & b[385])^(a[207] & b[386])^(a[206] & b[387])^(a[205] & b[388])^(a[204] & b[389])^(a[203] & b[390])^(a[202] & b[391])^(a[201] & b[392])^(a[200] & b[393])^(a[199] & b[394])^(a[198] & b[395])^(a[197] & b[396])^(a[196] & b[397])^(a[195] & b[398])^(a[194] & b[399])^(a[193] & b[400])^(a[192] & b[401])^(a[191] & b[402])^(a[190] & b[403])^(a[189] & b[404])^(a[188] & b[405])^(a[187] & b[406])^(a[186] & b[407])^(a[185] & b[408]);
assign y[594] = (a[408] & b[186])^(a[407] & b[187])^(a[406] & b[188])^(a[405] & b[189])^(a[404] & b[190])^(a[403] & b[191])^(a[402] & b[192])^(a[401] & b[193])^(a[400] & b[194])^(a[399] & b[195])^(a[398] & b[196])^(a[397] & b[197])^(a[396] & b[198])^(a[395] & b[199])^(a[394] & b[200])^(a[393] & b[201])^(a[392] & b[202])^(a[391] & b[203])^(a[390] & b[204])^(a[389] & b[205])^(a[388] & b[206])^(a[387] & b[207])^(a[386] & b[208])^(a[385] & b[209])^(a[384] & b[210])^(a[383] & b[211])^(a[382] & b[212])^(a[381] & b[213])^(a[380] & b[214])^(a[379] & b[215])^(a[378] & b[216])^(a[377] & b[217])^(a[376] & b[218])^(a[375] & b[219])^(a[374] & b[220])^(a[373] & b[221])^(a[372] & b[222])^(a[371] & b[223])^(a[370] & b[224])^(a[369] & b[225])^(a[368] & b[226])^(a[367] & b[227])^(a[366] & b[228])^(a[365] & b[229])^(a[364] & b[230])^(a[363] & b[231])^(a[362] & b[232])^(a[361] & b[233])^(a[360] & b[234])^(a[359] & b[235])^(a[358] & b[236])^(a[357] & b[237])^(a[356] & b[238])^(a[355] & b[239])^(a[354] & b[240])^(a[353] & b[241])^(a[352] & b[242])^(a[351] & b[243])^(a[350] & b[244])^(a[349] & b[245])^(a[348] & b[246])^(a[347] & b[247])^(a[346] & b[248])^(a[345] & b[249])^(a[344] & b[250])^(a[343] & b[251])^(a[342] & b[252])^(a[341] & b[253])^(a[340] & b[254])^(a[339] & b[255])^(a[338] & b[256])^(a[337] & b[257])^(a[336] & b[258])^(a[335] & b[259])^(a[334] & b[260])^(a[333] & b[261])^(a[332] & b[262])^(a[331] & b[263])^(a[330] & b[264])^(a[329] & b[265])^(a[328] & b[266])^(a[327] & b[267])^(a[326] & b[268])^(a[325] & b[269])^(a[324] & b[270])^(a[323] & b[271])^(a[322] & b[272])^(a[321] & b[273])^(a[320] & b[274])^(a[319] & b[275])^(a[318] & b[276])^(a[317] & b[277])^(a[316] & b[278])^(a[315] & b[279])^(a[314] & b[280])^(a[313] & b[281])^(a[312] & b[282])^(a[311] & b[283])^(a[310] & b[284])^(a[309] & b[285])^(a[308] & b[286])^(a[307] & b[287])^(a[306] & b[288])^(a[305] & b[289])^(a[304] & b[290])^(a[303] & b[291])^(a[302] & b[292])^(a[301] & b[293])^(a[300] & b[294])^(a[299] & b[295])^(a[298] & b[296])^(a[297] & b[297])^(a[296] & b[298])^(a[295] & b[299])^(a[294] & b[300])^(a[293] & b[301])^(a[292] & b[302])^(a[291] & b[303])^(a[290] & b[304])^(a[289] & b[305])^(a[288] & b[306])^(a[287] & b[307])^(a[286] & b[308])^(a[285] & b[309])^(a[284] & b[310])^(a[283] & b[311])^(a[282] & b[312])^(a[281] & b[313])^(a[280] & b[314])^(a[279] & b[315])^(a[278] & b[316])^(a[277] & b[317])^(a[276] & b[318])^(a[275] & b[319])^(a[274] & b[320])^(a[273] & b[321])^(a[272] & b[322])^(a[271] & b[323])^(a[270] & b[324])^(a[269] & b[325])^(a[268] & b[326])^(a[267] & b[327])^(a[266] & b[328])^(a[265] & b[329])^(a[264] & b[330])^(a[263] & b[331])^(a[262] & b[332])^(a[261] & b[333])^(a[260] & b[334])^(a[259] & b[335])^(a[258] & b[336])^(a[257] & b[337])^(a[256] & b[338])^(a[255] & b[339])^(a[254] & b[340])^(a[253] & b[341])^(a[252] & b[342])^(a[251] & b[343])^(a[250] & b[344])^(a[249] & b[345])^(a[248] & b[346])^(a[247] & b[347])^(a[246] & b[348])^(a[245] & b[349])^(a[244] & b[350])^(a[243] & b[351])^(a[242] & b[352])^(a[241] & b[353])^(a[240] & b[354])^(a[239] & b[355])^(a[238] & b[356])^(a[237] & b[357])^(a[236] & b[358])^(a[235] & b[359])^(a[234] & b[360])^(a[233] & b[361])^(a[232] & b[362])^(a[231] & b[363])^(a[230] & b[364])^(a[229] & b[365])^(a[228] & b[366])^(a[227] & b[367])^(a[226] & b[368])^(a[225] & b[369])^(a[224] & b[370])^(a[223] & b[371])^(a[222] & b[372])^(a[221] & b[373])^(a[220] & b[374])^(a[219] & b[375])^(a[218] & b[376])^(a[217] & b[377])^(a[216] & b[378])^(a[215] & b[379])^(a[214] & b[380])^(a[213] & b[381])^(a[212] & b[382])^(a[211] & b[383])^(a[210] & b[384])^(a[209] & b[385])^(a[208] & b[386])^(a[207] & b[387])^(a[206] & b[388])^(a[205] & b[389])^(a[204] & b[390])^(a[203] & b[391])^(a[202] & b[392])^(a[201] & b[393])^(a[200] & b[394])^(a[199] & b[395])^(a[198] & b[396])^(a[197] & b[397])^(a[196] & b[398])^(a[195] & b[399])^(a[194] & b[400])^(a[193] & b[401])^(a[192] & b[402])^(a[191] & b[403])^(a[190] & b[404])^(a[189] & b[405])^(a[188] & b[406])^(a[187] & b[407])^(a[186] & b[408]);
assign y[595] = (a[408] & b[187])^(a[407] & b[188])^(a[406] & b[189])^(a[405] & b[190])^(a[404] & b[191])^(a[403] & b[192])^(a[402] & b[193])^(a[401] & b[194])^(a[400] & b[195])^(a[399] & b[196])^(a[398] & b[197])^(a[397] & b[198])^(a[396] & b[199])^(a[395] & b[200])^(a[394] & b[201])^(a[393] & b[202])^(a[392] & b[203])^(a[391] & b[204])^(a[390] & b[205])^(a[389] & b[206])^(a[388] & b[207])^(a[387] & b[208])^(a[386] & b[209])^(a[385] & b[210])^(a[384] & b[211])^(a[383] & b[212])^(a[382] & b[213])^(a[381] & b[214])^(a[380] & b[215])^(a[379] & b[216])^(a[378] & b[217])^(a[377] & b[218])^(a[376] & b[219])^(a[375] & b[220])^(a[374] & b[221])^(a[373] & b[222])^(a[372] & b[223])^(a[371] & b[224])^(a[370] & b[225])^(a[369] & b[226])^(a[368] & b[227])^(a[367] & b[228])^(a[366] & b[229])^(a[365] & b[230])^(a[364] & b[231])^(a[363] & b[232])^(a[362] & b[233])^(a[361] & b[234])^(a[360] & b[235])^(a[359] & b[236])^(a[358] & b[237])^(a[357] & b[238])^(a[356] & b[239])^(a[355] & b[240])^(a[354] & b[241])^(a[353] & b[242])^(a[352] & b[243])^(a[351] & b[244])^(a[350] & b[245])^(a[349] & b[246])^(a[348] & b[247])^(a[347] & b[248])^(a[346] & b[249])^(a[345] & b[250])^(a[344] & b[251])^(a[343] & b[252])^(a[342] & b[253])^(a[341] & b[254])^(a[340] & b[255])^(a[339] & b[256])^(a[338] & b[257])^(a[337] & b[258])^(a[336] & b[259])^(a[335] & b[260])^(a[334] & b[261])^(a[333] & b[262])^(a[332] & b[263])^(a[331] & b[264])^(a[330] & b[265])^(a[329] & b[266])^(a[328] & b[267])^(a[327] & b[268])^(a[326] & b[269])^(a[325] & b[270])^(a[324] & b[271])^(a[323] & b[272])^(a[322] & b[273])^(a[321] & b[274])^(a[320] & b[275])^(a[319] & b[276])^(a[318] & b[277])^(a[317] & b[278])^(a[316] & b[279])^(a[315] & b[280])^(a[314] & b[281])^(a[313] & b[282])^(a[312] & b[283])^(a[311] & b[284])^(a[310] & b[285])^(a[309] & b[286])^(a[308] & b[287])^(a[307] & b[288])^(a[306] & b[289])^(a[305] & b[290])^(a[304] & b[291])^(a[303] & b[292])^(a[302] & b[293])^(a[301] & b[294])^(a[300] & b[295])^(a[299] & b[296])^(a[298] & b[297])^(a[297] & b[298])^(a[296] & b[299])^(a[295] & b[300])^(a[294] & b[301])^(a[293] & b[302])^(a[292] & b[303])^(a[291] & b[304])^(a[290] & b[305])^(a[289] & b[306])^(a[288] & b[307])^(a[287] & b[308])^(a[286] & b[309])^(a[285] & b[310])^(a[284] & b[311])^(a[283] & b[312])^(a[282] & b[313])^(a[281] & b[314])^(a[280] & b[315])^(a[279] & b[316])^(a[278] & b[317])^(a[277] & b[318])^(a[276] & b[319])^(a[275] & b[320])^(a[274] & b[321])^(a[273] & b[322])^(a[272] & b[323])^(a[271] & b[324])^(a[270] & b[325])^(a[269] & b[326])^(a[268] & b[327])^(a[267] & b[328])^(a[266] & b[329])^(a[265] & b[330])^(a[264] & b[331])^(a[263] & b[332])^(a[262] & b[333])^(a[261] & b[334])^(a[260] & b[335])^(a[259] & b[336])^(a[258] & b[337])^(a[257] & b[338])^(a[256] & b[339])^(a[255] & b[340])^(a[254] & b[341])^(a[253] & b[342])^(a[252] & b[343])^(a[251] & b[344])^(a[250] & b[345])^(a[249] & b[346])^(a[248] & b[347])^(a[247] & b[348])^(a[246] & b[349])^(a[245] & b[350])^(a[244] & b[351])^(a[243] & b[352])^(a[242] & b[353])^(a[241] & b[354])^(a[240] & b[355])^(a[239] & b[356])^(a[238] & b[357])^(a[237] & b[358])^(a[236] & b[359])^(a[235] & b[360])^(a[234] & b[361])^(a[233] & b[362])^(a[232] & b[363])^(a[231] & b[364])^(a[230] & b[365])^(a[229] & b[366])^(a[228] & b[367])^(a[227] & b[368])^(a[226] & b[369])^(a[225] & b[370])^(a[224] & b[371])^(a[223] & b[372])^(a[222] & b[373])^(a[221] & b[374])^(a[220] & b[375])^(a[219] & b[376])^(a[218] & b[377])^(a[217] & b[378])^(a[216] & b[379])^(a[215] & b[380])^(a[214] & b[381])^(a[213] & b[382])^(a[212] & b[383])^(a[211] & b[384])^(a[210] & b[385])^(a[209] & b[386])^(a[208] & b[387])^(a[207] & b[388])^(a[206] & b[389])^(a[205] & b[390])^(a[204] & b[391])^(a[203] & b[392])^(a[202] & b[393])^(a[201] & b[394])^(a[200] & b[395])^(a[199] & b[396])^(a[198] & b[397])^(a[197] & b[398])^(a[196] & b[399])^(a[195] & b[400])^(a[194] & b[401])^(a[193] & b[402])^(a[192] & b[403])^(a[191] & b[404])^(a[190] & b[405])^(a[189] & b[406])^(a[188] & b[407])^(a[187] & b[408]);
assign y[596] = (a[408] & b[188])^(a[407] & b[189])^(a[406] & b[190])^(a[405] & b[191])^(a[404] & b[192])^(a[403] & b[193])^(a[402] & b[194])^(a[401] & b[195])^(a[400] & b[196])^(a[399] & b[197])^(a[398] & b[198])^(a[397] & b[199])^(a[396] & b[200])^(a[395] & b[201])^(a[394] & b[202])^(a[393] & b[203])^(a[392] & b[204])^(a[391] & b[205])^(a[390] & b[206])^(a[389] & b[207])^(a[388] & b[208])^(a[387] & b[209])^(a[386] & b[210])^(a[385] & b[211])^(a[384] & b[212])^(a[383] & b[213])^(a[382] & b[214])^(a[381] & b[215])^(a[380] & b[216])^(a[379] & b[217])^(a[378] & b[218])^(a[377] & b[219])^(a[376] & b[220])^(a[375] & b[221])^(a[374] & b[222])^(a[373] & b[223])^(a[372] & b[224])^(a[371] & b[225])^(a[370] & b[226])^(a[369] & b[227])^(a[368] & b[228])^(a[367] & b[229])^(a[366] & b[230])^(a[365] & b[231])^(a[364] & b[232])^(a[363] & b[233])^(a[362] & b[234])^(a[361] & b[235])^(a[360] & b[236])^(a[359] & b[237])^(a[358] & b[238])^(a[357] & b[239])^(a[356] & b[240])^(a[355] & b[241])^(a[354] & b[242])^(a[353] & b[243])^(a[352] & b[244])^(a[351] & b[245])^(a[350] & b[246])^(a[349] & b[247])^(a[348] & b[248])^(a[347] & b[249])^(a[346] & b[250])^(a[345] & b[251])^(a[344] & b[252])^(a[343] & b[253])^(a[342] & b[254])^(a[341] & b[255])^(a[340] & b[256])^(a[339] & b[257])^(a[338] & b[258])^(a[337] & b[259])^(a[336] & b[260])^(a[335] & b[261])^(a[334] & b[262])^(a[333] & b[263])^(a[332] & b[264])^(a[331] & b[265])^(a[330] & b[266])^(a[329] & b[267])^(a[328] & b[268])^(a[327] & b[269])^(a[326] & b[270])^(a[325] & b[271])^(a[324] & b[272])^(a[323] & b[273])^(a[322] & b[274])^(a[321] & b[275])^(a[320] & b[276])^(a[319] & b[277])^(a[318] & b[278])^(a[317] & b[279])^(a[316] & b[280])^(a[315] & b[281])^(a[314] & b[282])^(a[313] & b[283])^(a[312] & b[284])^(a[311] & b[285])^(a[310] & b[286])^(a[309] & b[287])^(a[308] & b[288])^(a[307] & b[289])^(a[306] & b[290])^(a[305] & b[291])^(a[304] & b[292])^(a[303] & b[293])^(a[302] & b[294])^(a[301] & b[295])^(a[300] & b[296])^(a[299] & b[297])^(a[298] & b[298])^(a[297] & b[299])^(a[296] & b[300])^(a[295] & b[301])^(a[294] & b[302])^(a[293] & b[303])^(a[292] & b[304])^(a[291] & b[305])^(a[290] & b[306])^(a[289] & b[307])^(a[288] & b[308])^(a[287] & b[309])^(a[286] & b[310])^(a[285] & b[311])^(a[284] & b[312])^(a[283] & b[313])^(a[282] & b[314])^(a[281] & b[315])^(a[280] & b[316])^(a[279] & b[317])^(a[278] & b[318])^(a[277] & b[319])^(a[276] & b[320])^(a[275] & b[321])^(a[274] & b[322])^(a[273] & b[323])^(a[272] & b[324])^(a[271] & b[325])^(a[270] & b[326])^(a[269] & b[327])^(a[268] & b[328])^(a[267] & b[329])^(a[266] & b[330])^(a[265] & b[331])^(a[264] & b[332])^(a[263] & b[333])^(a[262] & b[334])^(a[261] & b[335])^(a[260] & b[336])^(a[259] & b[337])^(a[258] & b[338])^(a[257] & b[339])^(a[256] & b[340])^(a[255] & b[341])^(a[254] & b[342])^(a[253] & b[343])^(a[252] & b[344])^(a[251] & b[345])^(a[250] & b[346])^(a[249] & b[347])^(a[248] & b[348])^(a[247] & b[349])^(a[246] & b[350])^(a[245] & b[351])^(a[244] & b[352])^(a[243] & b[353])^(a[242] & b[354])^(a[241] & b[355])^(a[240] & b[356])^(a[239] & b[357])^(a[238] & b[358])^(a[237] & b[359])^(a[236] & b[360])^(a[235] & b[361])^(a[234] & b[362])^(a[233] & b[363])^(a[232] & b[364])^(a[231] & b[365])^(a[230] & b[366])^(a[229] & b[367])^(a[228] & b[368])^(a[227] & b[369])^(a[226] & b[370])^(a[225] & b[371])^(a[224] & b[372])^(a[223] & b[373])^(a[222] & b[374])^(a[221] & b[375])^(a[220] & b[376])^(a[219] & b[377])^(a[218] & b[378])^(a[217] & b[379])^(a[216] & b[380])^(a[215] & b[381])^(a[214] & b[382])^(a[213] & b[383])^(a[212] & b[384])^(a[211] & b[385])^(a[210] & b[386])^(a[209] & b[387])^(a[208] & b[388])^(a[207] & b[389])^(a[206] & b[390])^(a[205] & b[391])^(a[204] & b[392])^(a[203] & b[393])^(a[202] & b[394])^(a[201] & b[395])^(a[200] & b[396])^(a[199] & b[397])^(a[198] & b[398])^(a[197] & b[399])^(a[196] & b[400])^(a[195] & b[401])^(a[194] & b[402])^(a[193] & b[403])^(a[192] & b[404])^(a[191] & b[405])^(a[190] & b[406])^(a[189] & b[407])^(a[188] & b[408]);
assign y[597] = (a[408] & b[189])^(a[407] & b[190])^(a[406] & b[191])^(a[405] & b[192])^(a[404] & b[193])^(a[403] & b[194])^(a[402] & b[195])^(a[401] & b[196])^(a[400] & b[197])^(a[399] & b[198])^(a[398] & b[199])^(a[397] & b[200])^(a[396] & b[201])^(a[395] & b[202])^(a[394] & b[203])^(a[393] & b[204])^(a[392] & b[205])^(a[391] & b[206])^(a[390] & b[207])^(a[389] & b[208])^(a[388] & b[209])^(a[387] & b[210])^(a[386] & b[211])^(a[385] & b[212])^(a[384] & b[213])^(a[383] & b[214])^(a[382] & b[215])^(a[381] & b[216])^(a[380] & b[217])^(a[379] & b[218])^(a[378] & b[219])^(a[377] & b[220])^(a[376] & b[221])^(a[375] & b[222])^(a[374] & b[223])^(a[373] & b[224])^(a[372] & b[225])^(a[371] & b[226])^(a[370] & b[227])^(a[369] & b[228])^(a[368] & b[229])^(a[367] & b[230])^(a[366] & b[231])^(a[365] & b[232])^(a[364] & b[233])^(a[363] & b[234])^(a[362] & b[235])^(a[361] & b[236])^(a[360] & b[237])^(a[359] & b[238])^(a[358] & b[239])^(a[357] & b[240])^(a[356] & b[241])^(a[355] & b[242])^(a[354] & b[243])^(a[353] & b[244])^(a[352] & b[245])^(a[351] & b[246])^(a[350] & b[247])^(a[349] & b[248])^(a[348] & b[249])^(a[347] & b[250])^(a[346] & b[251])^(a[345] & b[252])^(a[344] & b[253])^(a[343] & b[254])^(a[342] & b[255])^(a[341] & b[256])^(a[340] & b[257])^(a[339] & b[258])^(a[338] & b[259])^(a[337] & b[260])^(a[336] & b[261])^(a[335] & b[262])^(a[334] & b[263])^(a[333] & b[264])^(a[332] & b[265])^(a[331] & b[266])^(a[330] & b[267])^(a[329] & b[268])^(a[328] & b[269])^(a[327] & b[270])^(a[326] & b[271])^(a[325] & b[272])^(a[324] & b[273])^(a[323] & b[274])^(a[322] & b[275])^(a[321] & b[276])^(a[320] & b[277])^(a[319] & b[278])^(a[318] & b[279])^(a[317] & b[280])^(a[316] & b[281])^(a[315] & b[282])^(a[314] & b[283])^(a[313] & b[284])^(a[312] & b[285])^(a[311] & b[286])^(a[310] & b[287])^(a[309] & b[288])^(a[308] & b[289])^(a[307] & b[290])^(a[306] & b[291])^(a[305] & b[292])^(a[304] & b[293])^(a[303] & b[294])^(a[302] & b[295])^(a[301] & b[296])^(a[300] & b[297])^(a[299] & b[298])^(a[298] & b[299])^(a[297] & b[300])^(a[296] & b[301])^(a[295] & b[302])^(a[294] & b[303])^(a[293] & b[304])^(a[292] & b[305])^(a[291] & b[306])^(a[290] & b[307])^(a[289] & b[308])^(a[288] & b[309])^(a[287] & b[310])^(a[286] & b[311])^(a[285] & b[312])^(a[284] & b[313])^(a[283] & b[314])^(a[282] & b[315])^(a[281] & b[316])^(a[280] & b[317])^(a[279] & b[318])^(a[278] & b[319])^(a[277] & b[320])^(a[276] & b[321])^(a[275] & b[322])^(a[274] & b[323])^(a[273] & b[324])^(a[272] & b[325])^(a[271] & b[326])^(a[270] & b[327])^(a[269] & b[328])^(a[268] & b[329])^(a[267] & b[330])^(a[266] & b[331])^(a[265] & b[332])^(a[264] & b[333])^(a[263] & b[334])^(a[262] & b[335])^(a[261] & b[336])^(a[260] & b[337])^(a[259] & b[338])^(a[258] & b[339])^(a[257] & b[340])^(a[256] & b[341])^(a[255] & b[342])^(a[254] & b[343])^(a[253] & b[344])^(a[252] & b[345])^(a[251] & b[346])^(a[250] & b[347])^(a[249] & b[348])^(a[248] & b[349])^(a[247] & b[350])^(a[246] & b[351])^(a[245] & b[352])^(a[244] & b[353])^(a[243] & b[354])^(a[242] & b[355])^(a[241] & b[356])^(a[240] & b[357])^(a[239] & b[358])^(a[238] & b[359])^(a[237] & b[360])^(a[236] & b[361])^(a[235] & b[362])^(a[234] & b[363])^(a[233] & b[364])^(a[232] & b[365])^(a[231] & b[366])^(a[230] & b[367])^(a[229] & b[368])^(a[228] & b[369])^(a[227] & b[370])^(a[226] & b[371])^(a[225] & b[372])^(a[224] & b[373])^(a[223] & b[374])^(a[222] & b[375])^(a[221] & b[376])^(a[220] & b[377])^(a[219] & b[378])^(a[218] & b[379])^(a[217] & b[380])^(a[216] & b[381])^(a[215] & b[382])^(a[214] & b[383])^(a[213] & b[384])^(a[212] & b[385])^(a[211] & b[386])^(a[210] & b[387])^(a[209] & b[388])^(a[208] & b[389])^(a[207] & b[390])^(a[206] & b[391])^(a[205] & b[392])^(a[204] & b[393])^(a[203] & b[394])^(a[202] & b[395])^(a[201] & b[396])^(a[200] & b[397])^(a[199] & b[398])^(a[198] & b[399])^(a[197] & b[400])^(a[196] & b[401])^(a[195] & b[402])^(a[194] & b[403])^(a[193] & b[404])^(a[192] & b[405])^(a[191] & b[406])^(a[190] & b[407])^(a[189] & b[408]);
assign y[598] = (a[408] & b[190])^(a[407] & b[191])^(a[406] & b[192])^(a[405] & b[193])^(a[404] & b[194])^(a[403] & b[195])^(a[402] & b[196])^(a[401] & b[197])^(a[400] & b[198])^(a[399] & b[199])^(a[398] & b[200])^(a[397] & b[201])^(a[396] & b[202])^(a[395] & b[203])^(a[394] & b[204])^(a[393] & b[205])^(a[392] & b[206])^(a[391] & b[207])^(a[390] & b[208])^(a[389] & b[209])^(a[388] & b[210])^(a[387] & b[211])^(a[386] & b[212])^(a[385] & b[213])^(a[384] & b[214])^(a[383] & b[215])^(a[382] & b[216])^(a[381] & b[217])^(a[380] & b[218])^(a[379] & b[219])^(a[378] & b[220])^(a[377] & b[221])^(a[376] & b[222])^(a[375] & b[223])^(a[374] & b[224])^(a[373] & b[225])^(a[372] & b[226])^(a[371] & b[227])^(a[370] & b[228])^(a[369] & b[229])^(a[368] & b[230])^(a[367] & b[231])^(a[366] & b[232])^(a[365] & b[233])^(a[364] & b[234])^(a[363] & b[235])^(a[362] & b[236])^(a[361] & b[237])^(a[360] & b[238])^(a[359] & b[239])^(a[358] & b[240])^(a[357] & b[241])^(a[356] & b[242])^(a[355] & b[243])^(a[354] & b[244])^(a[353] & b[245])^(a[352] & b[246])^(a[351] & b[247])^(a[350] & b[248])^(a[349] & b[249])^(a[348] & b[250])^(a[347] & b[251])^(a[346] & b[252])^(a[345] & b[253])^(a[344] & b[254])^(a[343] & b[255])^(a[342] & b[256])^(a[341] & b[257])^(a[340] & b[258])^(a[339] & b[259])^(a[338] & b[260])^(a[337] & b[261])^(a[336] & b[262])^(a[335] & b[263])^(a[334] & b[264])^(a[333] & b[265])^(a[332] & b[266])^(a[331] & b[267])^(a[330] & b[268])^(a[329] & b[269])^(a[328] & b[270])^(a[327] & b[271])^(a[326] & b[272])^(a[325] & b[273])^(a[324] & b[274])^(a[323] & b[275])^(a[322] & b[276])^(a[321] & b[277])^(a[320] & b[278])^(a[319] & b[279])^(a[318] & b[280])^(a[317] & b[281])^(a[316] & b[282])^(a[315] & b[283])^(a[314] & b[284])^(a[313] & b[285])^(a[312] & b[286])^(a[311] & b[287])^(a[310] & b[288])^(a[309] & b[289])^(a[308] & b[290])^(a[307] & b[291])^(a[306] & b[292])^(a[305] & b[293])^(a[304] & b[294])^(a[303] & b[295])^(a[302] & b[296])^(a[301] & b[297])^(a[300] & b[298])^(a[299] & b[299])^(a[298] & b[300])^(a[297] & b[301])^(a[296] & b[302])^(a[295] & b[303])^(a[294] & b[304])^(a[293] & b[305])^(a[292] & b[306])^(a[291] & b[307])^(a[290] & b[308])^(a[289] & b[309])^(a[288] & b[310])^(a[287] & b[311])^(a[286] & b[312])^(a[285] & b[313])^(a[284] & b[314])^(a[283] & b[315])^(a[282] & b[316])^(a[281] & b[317])^(a[280] & b[318])^(a[279] & b[319])^(a[278] & b[320])^(a[277] & b[321])^(a[276] & b[322])^(a[275] & b[323])^(a[274] & b[324])^(a[273] & b[325])^(a[272] & b[326])^(a[271] & b[327])^(a[270] & b[328])^(a[269] & b[329])^(a[268] & b[330])^(a[267] & b[331])^(a[266] & b[332])^(a[265] & b[333])^(a[264] & b[334])^(a[263] & b[335])^(a[262] & b[336])^(a[261] & b[337])^(a[260] & b[338])^(a[259] & b[339])^(a[258] & b[340])^(a[257] & b[341])^(a[256] & b[342])^(a[255] & b[343])^(a[254] & b[344])^(a[253] & b[345])^(a[252] & b[346])^(a[251] & b[347])^(a[250] & b[348])^(a[249] & b[349])^(a[248] & b[350])^(a[247] & b[351])^(a[246] & b[352])^(a[245] & b[353])^(a[244] & b[354])^(a[243] & b[355])^(a[242] & b[356])^(a[241] & b[357])^(a[240] & b[358])^(a[239] & b[359])^(a[238] & b[360])^(a[237] & b[361])^(a[236] & b[362])^(a[235] & b[363])^(a[234] & b[364])^(a[233] & b[365])^(a[232] & b[366])^(a[231] & b[367])^(a[230] & b[368])^(a[229] & b[369])^(a[228] & b[370])^(a[227] & b[371])^(a[226] & b[372])^(a[225] & b[373])^(a[224] & b[374])^(a[223] & b[375])^(a[222] & b[376])^(a[221] & b[377])^(a[220] & b[378])^(a[219] & b[379])^(a[218] & b[380])^(a[217] & b[381])^(a[216] & b[382])^(a[215] & b[383])^(a[214] & b[384])^(a[213] & b[385])^(a[212] & b[386])^(a[211] & b[387])^(a[210] & b[388])^(a[209] & b[389])^(a[208] & b[390])^(a[207] & b[391])^(a[206] & b[392])^(a[205] & b[393])^(a[204] & b[394])^(a[203] & b[395])^(a[202] & b[396])^(a[201] & b[397])^(a[200] & b[398])^(a[199] & b[399])^(a[198] & b[400])^(a[197] & b[401])^(a[196] & b[402])^(a[195] & b[403])^(a[194] & b[404])^(a[193] & b[405])^(a[192] & b[406])^(a[191] & b[407])^(a[190] & b[408]);
assign y[599] = (a[408] & b[191])^(a[407] & b[192])^(a[406] & b[193])^(a[405] & b[194])^(a[404] & b[195])^(a[403] & b[196])^(a[402] & b[197])^(a[401] & b[198])^(a[400] & b[199])^(a[399] & b[200])^(a[398] & b[201])^(a[397] & b[202])^(a[396] & b[203])^(a[395] & b[204])^(a[394] & b[205])^(a[393] & b[206])^(a[392] & b[207])^(a[391] & b[208])^(a[390] & b[209])^(a[389] & b[210])^(a[388] & b[211])^(a[387] & b[212])^(a[386] & b[213])^(a[385] & b[214])^(a[384] & b[215])^(a[383] & b[216])^(a[382] & b[217])^(a[381] & b[218])^(a[380] & b[219])^(a[379] & b[220])^(a[378] & b[221])^(a[377] & b[222])^(a[376] & b[223])^(a[375] & b[224])^(a[374] & b[225])^(a[373] & b[226])^(a[372] & b[227])^(a[371] & b[228])^(a[370] & b[229])^(a[369] & b[230])^(a[368] & b[231])^(a[367] & b[232])^(a[366] & b[233])^(a[365] & b[234])^(a[364] & b[235])^(a[363] & b[236])^(a[362] & b[237])^(a[361] & b[238])^(a[360] & b[239])^(a[359] & b[240])^(a[358] & b[241])^(a[357] & b[242])^(a[356] & b[243])^(a[355] & b[244])^(a[354] & b[245])^(a[353] & b[246])^(a[352] & b[247])^(a[351] & b[248])^(a[350] & b[249])^(a[349] & b[250])^(a[348] & b[251])^(a[347] & b[252])^(a[346] & b[253])^(a[345] & b[254])^(a[344] & b[255])^(a[343] & b[256])^(a[342] & b[257])^(a[341] & b[258])^(a[340] & b[259])^(a[339] & b[260])^(a[338] & b[261])^(a[337] & b[262])^(a[336] & b[263])^(a[335] & b[264])^(a[334] & b[265])^(a[333] & b[266])^(a[332] & b[267])^(a[331] & b[268])^(a[330] & b[269])^(a[329] & b[270])^(a[328] & b[271])^(a[327] & b[272])^(a[326] & b[273])^(a[325] & b[274])^(a[324] & b[275])^(a[323] & b[276])^(a[322] & b[277])^(a[321] & b[278])^(a[320] & b[279])^(a[319] & b[280])^(a[318] & b[281])^(a[317] & b[282])^(a[316] & b[283])^(a[315] & b[284])^(a[314] & b[285])^(a[313] & b[286])^(a[312] & b[287])^(a[311] & b[288])^(a[310] & b[289])^(a[309] & b[290])^(a[308] & b[291])^(a[307] & b[292])^(a[306] & b[293])^(a[305] & b[294])^(a[304] & b[295])^(a[303] & b[296])^(a[302] & b[297])^(a[301] & b[298])^(a[300] & b[299])^(a[299] & b[300])^(a[298] & b[301])^(a[297] & b[302])^(a[296] & b[303])^(a[295] & b[304])^(a[294] & b[305])^(a[293] & b[306])^(a[292] & b[307])^(a[291] & b[308])^(a[290] & b[309])^(a[289] & b[310])^(a[288] & b[311])^(a[287] & b[312])^(a[286] & b[313])^(a[285] & b[314])^(a[284] & b[315])^(a[283] & b[316])^(a[282] & b[317])^(a[281] & b[318])^(a[280] & b[319])^(a[279] & b[320])^(a[278] & b[321])^(a[277] & b[322])^(a[276] & b[323])^(a[275] & b[324])^(a[274] & b[325])^(a[273] & b[326])^(a[272] & b[327])^(a[271] & b[328])^(a[270] & b[329])^(a[269] & b[330])^(a[268] & b[331])^(a[267] & b[332])^(a[266] & b[333])^(a[265] & b[334])^(a[264] & b[335])^(a[263] & b[336])^(a[262] & b[337])^(a[261] & b[338])^(a[260] & b[339])^(a[259] & b[340])^(a[258] & b[341])^(a[257] & b[342])^(a[256] & b[343])^(a[255] & b[344])^(a[254] & b[345])^(a[253] & b[346])^(a[252] & b[347])^(a[251] & b[348])^(a[250] & b[349])^(a[249] & b[350])^(a[248] & b[351])^(a[247] & b[352])^(a[246] & b[353])^(a[245] & b[354])^(a[244] & b[355])^(a[243] & b[356])^(a[242] & b[357])^(a[241] & b[358])^(a[240] & b[359])^(a[239] & b[360])^(a[238] & b[361])^(a[237] & b[362])^(a[236] & b[363])^(a[235] & b[364])^(a[234] & b[365])^(a[233] & b[366])^(a[232] & b[367])^(a[231] & b[368])^(a[230] & b[369])^(a[229] & b[370])^(a[228] & b[371])^(a[227] & b[372])^(a[226] & b[373])^(a[225] & b[374])^(a[224] & b[375])^(a[223] & b[376])^(a[222] & b[377])^(a[221] & b[378])^(a[220] & b[379])^(a[219] & b[380])^(a[218] & b[381])^(a[217] & b[382])^(a[216] & b[383])^(a[215] & b[384])^(a[214] & b[385])^(a[213] & b[386])^(a[212] & b[387])^(a[211] & b[388])^(a[210] & b[389])^(a[209] & b[390])^(a[208] & b[391])^(a[207] & b[392])^(a[206] & b[393])^(a[205] & b[394])^(a[204] & b[395])^(a[203] & b[396])^(a[202] & b[397])^(a[201] & b[398])^(a[200] & b[399])^(a[199] & b[400])^(a[198] & b[401])^(a[197] & b[402])^(a[196] & b[403])^(a[195] & b[404])^(a[194] & b[405])^(a[193] & b[406])^(a[192] & b[407])^(a[191] & b[408]);
assign y[600] = (a[408] & b[192])^(a[407] & b[193])^(a[406] & b[194])^(a[405] & b[195])^(a[404] & b[196])^(a[403] & b[197])^(a[402] & b[198])^(a[401] & b[199])^(a[400] & b[200])^(a[399] & b[201])^(a[398] & b[202])^(a[397] & b[203])^(a[396] & b[204])^(a[395] & b[205])^(a[394] & b[206])^(a[393] & b[207])^(a[392] & b[208])^(a[391] & b[209])^(a[390] & b[210])^(a[389] & b[211])^(a[388] & b[212])^(a[387] & b[213])^(a[386] & b[214])^(a[385] & b[215])^(a[384] & b[216])^(a[383] & b[217])^(a[382] & b[218])^(a[381] & b[219])^(a[380] & b[220])^(a[379] & b[221])^(a[378] & b[222])^(a[377] & b[223])^(a[376] & b[224])^(a[375] & b[225])^(a[374] & b[226])^(a[373] & b[227])^(a[372] & b[228])^(a[371] & b[229])^(a[370] & b[230])^(a[369] & b[231])^(a[368] & b[232])^(a[367] & b[233])^(a[366] & b[234])^(a[365] & b[235])^(a[364] & b[236])^(a[363] & b[237])^(a[362] & b[238])^(a[361] & b[239])^(a[360] & b[240])^(a[359] & b[241])^(a[358] & b[242])^(a[357] & b[243])^(a[356] & b[244])^(a[355] & b[245])^(a[354] & b[246])^(a[353] & b[247])^(a[352] & b[248])^(a[351] & b[249])^(a[350] & b[250])^(a[349] & b[251])^(a[348] & b[252])^(a[347] & b[253])^(a[346] & b[254])^(a[345] & b[255])^(a[344] & b[256])^(a[343] & b[257])^(a[342] & b[258])^(a[341] & b[259])^(a[340] & b[260])^(a[339] & b[261])^(a[338] & b[262])^(a[337] & b[263])^(a[336] & b[264])^(a[335] & b[265])^(a[334] & b[266])^(a[333] & b[267])^(a[332] & b[268])^(a[331] & b[269])^(a[330] & b[270])^(a[329] & b[271])^(a[328] & b[272])^(a[327] & b[273])^(a[326] & b[274])^(a[325] & b[275])^(a[324] & b[276])^(a[323] & b[277])^(a[322] & b[278])^(a[321] & b[279])^(a[320] & b[280])^(a[319] & b[281])^(a[318] & b[282])^(a[317] & b[283])^(a[316] & b[284])^(a[315] & b[285])^(a[314] & b[286])^(a[313] & b[287])^(a[312] & b[288])^(a[311] & b[289])^(a[310] & b[290])^(a[309] & b[291])^(a[308] & b[292])^(a[307] & b[293])^(a[306] & b[294])^(a[305] & b[295])^(a[304] & b[296])^(a[303] & b[297])^(a[302] & b[298])^(a[301] & b[299])^(a[300] & b[300])^(a[299] & b[301])^(a[298] & b[302])^(a[297] & b[303])^(a[296] & b[304])^(a[295] & b[305])^(a[294] & b[306])^(a[293] & b[307])^(a[292] & b[308])^(a[291] & b[309])^(a[290] & b[310])^(a[289] & b[311])^(a[288] & b[312])^(a[287] & b[313])^(a[286] & b[314])^(a[285] & b[315])^(a[284] & b[316])^(a[283] & b[317])^(a[282] & b[318])^(a[281] & b[319])^(a[280] & b[320])^(a[279] & b[321])^(a[278] & b[322])^(a[277] & b[323])^(a[276] & b[324])^(a[275] & b[325])^(a[274] & b[326])^(a[273] & b[327])^(a[272] & b[328])^(a[271] & b[329])^(a[270] & b[330])^(a[269] & b[331])^(a[268] & b[332])^(a[267] & b[333])^(a[266] & b[334])^(a[265] & b[335])^(a[264] & b[336])^(a[263] & b[337])^(a[262] & b[338])^(a[261] & b[339])^(a[260] & b[340])^(a[259] & b[341])^(a[258] & b[342])^(a[257] & b[343])^(a[256] & b[344])^(a[255] & b[345])^(a[254] & b[346])^(a[253] & b[347])^(a[252] & b[348])^(a[251] & b[349])^(a[250] & b[350])^(a[249] & b[351])^(a[248] & b[352])^(a[247] & b[353])^(a[246] & b[354])^(a[245] & b[355])^(a[244] & b[356])^(a[243] & b[357])^(a[242] & b[358])^(a[241] & b[359])^(a[240] & b[360])^(a[239] & b[361])^(a[238] & b[362])^(a[237] & b[363])^(a[236] & b[364])^(a[235] & b[365])^(a[234] & b[366])^(a[233] & b[367])^(a[232] & b[368])^(a[231] & b[369])^(a[230] & b[370])^(a[229] & b[371])^(a[228] & b[372])^(a[227] & b[373])^(a[226] & b[374])^(a[225] & b[375])^(a[224] & b[376])^(a[223] & b[377])^(a[222] & b[378])^(a[221] & b[379])^(a[220] & b[380])^(a[219] & b[381])^(a[218] & b[382])^(a[217] & b[383])^(a[216] & b[384])^(a[215] & b[385])^(a[214] & b[386])^(a[213] & b[387])^(a[212] & b[388])^(a[211] & b[389])^(a[210] & b[390])^(a[209] & b[391])^(a[208] & b[392])^(a[207] & b[393])^(a[206] & b[394])^(a[205] & b[395])^(a[204] & b[396])^(a[203] & b[397])^(a[202] & b[398])^(a[201] & b[399])^(a[200] & b[400])^(a[199] & b[401])^(a[198] & b[402])^(a[197] & b[403])^(a[196] & b[404])^(a[195] & b[405])^(a[194] & b[406])^(a[193] & b[407])^(a[192] & b[408]);
assign y[601] = (a[408] & b[193])^(a[407] & b[194])^(a[406] & b[195])^(a[405] & b[196])^(a[404] & b[197])^(a[403] & b[198])^(a[402] & b[199])^(a[401] & b[200])^(a[400] & b[201])^(a[399] & b[202])^(a[398] & b[203])^(a[397] & b[204])^(a[396] & b[205])^(a[395] & b[206])^(a[394] & b[207])^(a[393] & b[208])^(a[392] & b[209])^(a[391] & b[210])^(a[390] & b[211])^(a[389] & b[212])^(a[388] & b[213])^(a[387] & b[214])^(a[386] & b[215])^(a[385] & b[216])^(a[384] & b[217])^(a[383] & b[218])^(a[382] & b[219])^(a[381] & b[220])^(a[380] & b[221])^(a[379] & b[222])^(a[378] & b[223])^(a[377] & b[224])^(a[376] & b[225])^(a[375] & b[226])^(a[374] & b[227])^(a[373] & b[228])^(a[372] & b[229])^(a[371] & b[230])^(a[370] & b[231])^(a[369] & b[232])^(a[368] & b[233])^(a[367] & b[234])^(a[366] & b[235])^(a[365] & b[236])^(a[364] & b[237])^(a[363] & b[238])^(a[362] & b[239])^(a[361] & b[240])^(a[360] & b[241])^(a[359] & b[242])^(a[358] & b[243])^(a[357] & b[244])^(a[356] & b[245])^(a[355] & b[246])^(a[354] & b[247])^(a[353] & b[248])^(a[352] & b[249])^(a[351] & b[250])^(a[350] & b[251])^(a[349] & b[252])^(a[348] & b[253])^(a[347] & b[254])^(a[346] & b[255])^(a[345] & b[256])^(a[344] & b[257])^(a[343] & b[258])^(a[342] & b[259])^(a[341] & b[260])^(a[340] & b[261])^(a[339] & b[262])^(a[338] & b[263])^(a[337] & b[264])^(a[336] & b[265])^(a[335] & b[266])^(a[334] & b[267])^(a[333] & b[268])^(a[332] & b[269])^(a[331] & b[270])^(a[330] & b[271])^(a[329] & b[272])^(a[328] & b[273])^(a[327] & b[274])^(a[326] & b[275])^(a[325] & b[276])^(a[324] & b[277])^(a[323] & b[278])^(a[322] & b[279])^(a[321] & b[280])^(a[320] & b[281])^(a[319] & b[282])^(a[318] & b[283])^(a[317] & b[284])^(a[316] & b[285])^(a[315] & b[286])^(a[314] & b[287])^(a[313] & b[288])^(a[312] & b[289])^(a[311] & b[290])^(a[310] & b[291])^(a[309] & b[292])^(a[308] & b[293])^(a[307] & b[294])^(a[306] & b[295])^(a[305] & b[296])^(a[304] & b[297])^(a[303] & b[298])^(a[302] & b[299])^(a[301] & b[300])^(a[300] & b[301])^(a[299] & b[302])^(a[298] & b[303])^(a[297] & b[304])^(a[296] & b[305])^(a[295] & b[306])^(a[294] & b[307])^(a[293] & b[308])^(a[292] & b[309])^(a[291] & b[310])^(a[290] & b[311])^(a[289] & b[312])^(a[288] & b[313])^(a[287] & b[314])^(a[286] & b[315])^(a[285] & b[316])^(a[284] & b[317])^(a[283] & b[318])^(a[282] & b[319])^(a[281] & b[320])^(a[280] & b[321])^(a[279] & b[322])^(a[278] & b[323])^(a[277] & b[324])^(a[276] & b[325])^(a[275] & b[326])^(a[274] & b[327])^(a[273] & b[328])^(a[272] & b[329])^(a[271] & b[330])^(a[270] & b[331])^(a[269] & b[332])^(a[268] & b[333])^(a[267] & b[334])^(a[266] & b[335])^(a[265] & b[336])^(a[264] & b[337])^(a[263] & b[338])^(a[262] & b[339])^(a[261] & b[340])^(a[260] & b[341])^(a[259] & b[342])^(a[258] & b[343])^(a[257] & b[344])^(a[256] & b[345])^(a[255] & b[346])^(a[254] & b[347])^(a[253] & b[348])^(a[252] & b[349])^(a[251] & b[350])^(a[250] & b[351])^(a[249] & b[352])^(a[248] & b[353])^(a[247] & b[354])^(a[246] & b[355])^(a[245] & b[356])^(a[244] & b[357])^(a[243] & b[358])^(a[242] & b[359])^(a[241] & b[360])^(a[240] & b[361])^(a[239] & b[362])^(a[238] & b[363])^(a[237] & b[364])^(a[236] & b[365])^(a[235] & b[366])^(a[234] & b[367])^(a[233] & b[368])^(a[232] & b[369])^(a[231] & b[370])^(a[230] & b[371])^(a[229] & b[372])^(a[228] & b[373])^(a[227] & b[374])^(a[226] & b[375])^(a[225] & b[376])^(a[224] & b[377])^(a[223] & b[378])^(a[222] & b[379])^(a[221] & b[380])^(a[220] & b[381])^(a[219] & b[382])^(a[218] & b[383])^(a[217] & b[384])^(a[216] & b[385])^(a[215] & b[386])^(a[214] & b[387])^(a[213] & b[388])^(a[212] & b[389])^(a[211] & b[390])^(a[210] & b[391])^(a[209] & b[392])^(a[208] & b[393])^(a[207] & b[394])^(a[206] & b[395])^(a[205] & b[396])^(a[204] & b[397])^(a[203] & b[398])^(a[202] & b[399])^(a[201] & b[400])^(a[200] & b[401])^(a[199] & b[402])^(a[198] & b[403])^(a[197] & b[404])^(a[196] & b[405])^(a[195] & b[406])^(a[194] & b[407])^(a[193] & b[408]);
assign y[602] = (a[408] & b[194])^(a[407] & b[195])^(a[406] & b[196])^(a[405] & b[197])^(a[404] & b[198])^(a[403] & b[199])^(a[402] & b[200])^(a[401] & b[201])^(a[400] & b[202])^(a[399] & b[203])^(a[398] & b[204])^(a[397] & b[205])^(a[396] & b[206])^(a[395] & b[207])^(a[394] & b[208])^(a[393] & b[209])^(a[392] & b[210])^(a[391] & b[211])^(a[390] & b[212])^(a[389] & b[213])^(a[388] & b[214])^(a[387] & b[215])^(a[386] & b[216])^(a[385] & b[217])^(a[384] & b[218])^(a[383] & b[219])^(a[382] & b[220])^(a[381] & b[221])^(a[380] & b[222])^(a[379] & b[223])^(a[378] & b[224])^(a[377] & b[225])^(a[376] & b[226])^(a[375] & b[227])^(a[374] & b[228])^(a[373] & b[229])^(a[372] & b[230])^(a[371] & b[231])^(a[370] & b[232])^(a[369] & b[233])^(a[368] & b[234])^(a[367] & b[235])^(a[366] & b[236])^(a[365] & b[237])^(a[364] & b[238])^(a[363] & b[239])^(a[362] & b[240])^(a[361] & b[241])^(a[360] & b[242])^(a[359] & b[243])^(a[358] & b[244])^(a[357] & b[245])^(a[356] & b[246])^(a[355] & b[247])^(a[354] & b[248])^(a[353] & b[249])^(a[352] & b[250])^(a[351] & b[251])^(a[350] & b[252])^(a[349] & b[253])^(a[348] & b[254])^(a[347] & b[255])^(a[346] & b[256])^(a[345] & b[257])^(a[344] & b[258])^(a[343] & b[259])^(a[342] & b[260])^(a[341] & b[261])^(a[340] & b[262])^(a[339] & b[263])^(a[338] & b[264])^(a[337] & b[265])^(a[336] & b[266])^(a[335] & b[267])^(a[334] & b[268])^(a[333] & b[269])^(a[332] & b[270])^(a[331] & b[271])^(a[330] & b[272])^(a[329] & b[273])^(a[328] & b[274])^(a[327] & b[275])^(a[326] & b[276])^(a[325] & b[277])^(a[324] & b[278])^(a[323] & b[279])^(a[322] & b[280])^(a[321] & b[281])^(a[320] & b[282])^(a[319] & b[283])^(a[318] & b[284])^(a[317] & b[285])^(a[316] & b[286])^(a[315] & b[287])^(a[314] & b[288])^(a[313] & b[289])^(a[312] & b[290])^(a[311] & b[291])^(a[310] & b[292])^(a[309] & b[293])^(a[308] & b[294])^(a[307] & b[295])^(a[306] & b[296])^(a[305] & b[297])^(a[304] & b[298])^(a[303] & b[299])^(a[302] & b[300])^(a[301] & b[301])^(a[300] & b[302])^(a[299] & b[303])^(a[298] & b[304])^(a[297] & b[305])^(a[296] & b[306])^(a[295] & b[307])^(a[294] & b[308])^(a[293] & b[309])^(a[292] & b[310])^(a[291] & b[311])^(a[290] & b[312])^(a[289] & b[313])^(a[288] & b[314])^(a[287] & b[315])^(a[286] & b[316])^(a[285] & b[317])^(a[284] & b[318])^(a[283] & b[319])^(a[282] & b[320])^(a[281] & b[321])^(a[280] & b[322])^(a[279] & b[323])^(a[278] & b[324])^(a[277] & b[325])^(a[276] & b[326])^(a[275] & b[327])^(a[274] & b[328])^(a[273] & b[329])^(a[272] & b[330])^(a[271] & b[331])^(a[270] & b[332])^(a[269] & b[333])^(a[268] & b[334])^(a[267] & b[335])^(a[266] & b[336])^(a[265] & b[337])^(a[264] & b[338])^(a[263] & b[339])^(a[262] & b[340])^(a[261] & b[341])^(a[260] & b[342])^(a[259] & b[343])^(a[258] & b[344])^(a[257] & b[345])^(a[256] & b[346])^(a[255] & b[347])^(a[254] & b[348])^(a[253] & b[349])^(a[252] & b[350])^(a[251] & b[351])^(a[250] & b[352])^(a[249] & b[353])^(a[248] & b[354])^(a[247] & b[355])^(a[246] & b[356])^(a[245] & b[357])^(a[244] & b[358])^(a[243] & b[359])^(a[242] & b[360])^(a[241] & b[361])^(a[240] & b[362])^(a[239] & b[363])^(a[238] & b[364])^(a[237] & b[365])^(a[236] & b[366])^(a[235] & b[367])^(a[234] & b[368])^(a[233] & b[369])^(a[232] & b[370])^(a[231] & b[371])^(a[230] & b[372])^(a[229] & b[373])^(a[228] & b[374])^(a[227] & b[375])^(a[226] & b[376])^(a[225] & b[377])^(a[224] & b[378])^(a[223] & b[379])^(a[222] & b[380])^(a[221] & b[381])^(a[220] & b[382])^(a[219] & b[383])^(a[218] & b[384])^(a[217] & b[385])^(a[216] & b[386])^(a[215] & b[387])^(a[214] & b[388])^(a[213] & b[389])^(a[212] & b[390])^(a[211] & b[391])^(a[210] & b[392])^(a[209] & b[393])^(a[208] & b[394])^(a[207] & b[395])^(a[206] & b[396])^(a[205] & b[397])^(a[204] & b[398])^(a[203] & b[399])^(a[202] & b[400])^(a[201] & b[401])^(a[200] & b[402])^(a[199] & b[403])^(a[198] & b[404])^(a[197] & b[405])^(a[196] & b[406])^(a[195] & b[407])^(a[194] & b[408]);
assign y[603] = (a[408] & b[195])^(a[407] & b[196])^(a[406] & b[197])^(a[405] & b[198])^(a[404] & b[199])^(a[403] & b[200])^(a[402] & b[201])^(a[401] & b[202])^(a[400] & b[203])^(a[399] & b[204])^(a[398] & b[205])^(a[397] & b[206])^(a[396] & b[207])^(a[395] & b[208])^(a[394] & b[209])^(a[393] & b[210])^(a[392] & b[211])^(a[391] & b[212])^(a[390] & b[213])^(a[389] & b[214])^(a[388] & b[215])^(a[387] & b[216])^(a[386] & b[217])^(a[385] & b[218])^(a[384] & b[219])^(a[383] & b[220])^(a[382] & b[221])^(a[381] & b[222])^(a[380] & b[223])^(a[379] & b[224])^(a[378] & b[225])^(a[377] & b[226])^(a[376] & b[227])^(a[375] & b[228])^(a[374] & b[229])^(a[373] & b[230])^(a[372] & b[231])^(a[371] & b[232])^(a[370] & b[233])^(a[369] & b[234])^(a[368] & b[235])^(a[367] & b[236])^(a[366] & b[237])^(a[365] & b[238])^(a[364] & b[239])^(a[363] & b[240])^(a[362] & b[241])^(a[361] & b[242])^(a[360] & b[243])^(a[359] & b[244])^(a[358] & b[245])^(a[357] & b[246])^(a[356] & b[247])^(a[355] & b[248])^(a[354] & b[249])^(a[353] & b[250])^(a[352] & b[251])^(a[351] & b[252])^(a[350] & b[253])^(a[349] & b[254])^(a[348] & b[255])^(a[347] & b[256])^(a[346] & b[257])^(a[345] & b[258])^(a[344] & b[259])^(a[343] & b[260])^(a[342] & b[261])^(a[341] & b[262])^(a[340] & b[263])^(a[339] & b[264])^(a[338] & b[265])^(a[337] & b[266])^(a[336] & b[267])^(a[335] & b[268])^(a[334] & b[269])^(a[333] & b[270])^(a[332] & b[271])^(a[331] & b[272])^(a[330] & b[273])^(a[329] & b[274])^(a[328] & b[275])^(a[327] & b[276])^(a[326] & b[277])^(a[325] & b[278])^(a[324] & b[279])^(a[323] & b[280])^(a[322] & b[281])^(a[321] & b[282])^(a[320] & b[283])^(a[319] & b[284])^(a[318] & b[285])^(a[317] & b[286])^(a[316] & b[287])^(a[315] & b[288])^(a[314] & b[289])^(a[313] & b[290])^(a[312] & b[291])^(a[311] & b[292])^(a[310] & b[293])^(a[309] & b[294])^(a[308] & b[295])^(a[307] & b[296])^(a[306] & b[297])^(a[305] & b[298])^(a[304] & b[299])^(a[303] & b[300])^(a[302] & b[301])^(a[301] & b[302])^(a[300] & b[303])^(a[299] & b[304])^(a[298] & b[305])^(a[297] & b[306])^(a[296] & b[307])^(a[295] & b[308])^(a[294] & b[309])^(a[293] & b[310])^(a[292] & b[311])^(a[291] & b[312])^(a[290] & b[313])^(a[289] & b[314])^(a[288] & b[315])^(a[287] & b[316])^(a[286] & b[317])^(a[285] & b[318])^(a[284] & b[319])^(a[283] & b[320])^(a[282] & b[321])^(a[281] & b[322])^(a[280] & b[323])^(a[279] & b[324])^(a[278] & b[325])^(a[277] & b[326])^(a[276] & b[327])^(a[275] & b[328])^(a[274] & b[329])^(a[273] & b[330])^(a[272] & b[331])^(a[271] & b[332])^(a[270] & b[333])^(a[269] & b[334])^(a[268] & b[335])^(a[267] & b[336])^(a[266] & b[337])^(a[265] & b[338])^(a[264] & b[339])^(a[263] & b[340])^(a[262] & b[341])^(a[261] & b[342])^(a[260] & b[343])^(a[259] & b[344])^(a[258] & b[345])^(a[257] & b[346])^(a[256] & b[347])^(a[255] & b[348])^(a[254] & b[349])^(a[253] & b[350])^(a[252] & b[351])^(a[251] & b[352])^(a[250] & b[353])^(a[249] & b[354])^(a[248] & b[355])^(a[247] & b[356])^(a[246] & b[357])^(a[245] & b[358])^(a[244] & b[359])^(a[243] & b[360])^(a[242] & b[361])^(a[241] & b[362])^(a[240] & b[363])^(a[239] & b[364])^(a[238] & b[365])^(a[237] & b[366])^(a[236] & b[367])^(a[235] & b[368])^(a[234] & b[369])^(a[233] & b[370])^(a[232] & b[371])^(a[231] & b[372])^(a[230] & b[373])^(a[229] & b[374])^(a[228] & b[375])^(a[227] & b[376])^(a[226] & b[377])^(a[225] & b[378])^(a[224] & b[379])^(a[223] & b[380])^(a[222] & b[381])^(a[221] & b[382])^(a[220] & b[383])^(a[219] & b[384])^(a[218] & b[385])^(a[217] & b[386])^(a[216] & b[387])^(a[215] & b[388])^(a[214] & b[389])^(a[213] & b[390])^(a[212] & b[391])^(a[211] & b[392])^(a[210] & b[393])^(a[209] & b[394])^(a[208] & b[395])^(a[207] & b[396])^(a[206] & b[397])^(a[205] & b[398])^(a[204] & b[399])^(a[203] & b[400])^(a[202] & b[401])^(a[201] & b[402])^(a[200] & b[403])^(a[199] & b[404])^(a[198] & b[405])^(a[197] & b[406])^(a[196] & b[407])^(a[195] & b[408]);
assign y[604] = (a[408] & b[196])^(a[407] & b[197])^(a[406] & b[198])^(a[405] & b[199])^(a[404] & b[200])^(a[403] & b[201])^(a[402] & b[202])^(a[401] & b[203])^(a[400] & b[204])^(a[399] & b[205])^(a[398] & b[206])^(a[397] & b[207])^(a[396] & b[208])^(a[395] & b[209])^(a[394] & b[210])^(a[393] & b[211])^(a[392] & b[212])^(a[391] & b[213])^(a[390] & b[214])^(a[389] & b[215])^(a[388] & b[216])^(a[387] & b[217])^(a[386] & b[218])^(a[385] & b[219])^(a[384] & b[220])^(a[383] & b[221])^(a[382] & b[222])^(a[381] & b[223])^(a[380] & b[224])^(a[379] & b[225])^(a[378] & b[226])^(a[377] & b[227])^(a[376] & b[228])^(a[375] & b[229])^(a[374] & b[230])^(a[373] & b[231])^(a[372] & b[232])^(a[371] & b[233])^(a[370] & b[234])^(a[369] & b[235])^(a[368] & b[236])^(a[367] & b[237])^(a[366] & b[238])^(a[365] & b[239])^(a[364] & b[240])^(a[363] & b[241])^(a[362] & b[242])^(a[361] & b[243])^(a[360] & b[244])^(a[359] & b[245])^(a[358] & b[246])^(a[357] & b[247])^(a[356] & b[248])^(a[355] & b[249])^(a[354] & b[250])^(a[353] & b[251])^(a[352] & b[252])^(a[351] & b[253])^(a[350] & b[254])^(a[349] & b[255])^(a[348] & b[256])^(a[347] & b[257])^(a[346] & b[258])^(a[345] & b[259])^(a[344] & b[260])^(a[343] & b[261])^(a[342] & b[262])^(a[341] & b[263])^(a[340] & b[264])^(a[339] & b[265])^(a[338] & b[266])^(a[337] & b[267])^(a[336] & b[268])^(a[335] & b[269])^(a[334] & b[270])^(a[333] & b[271])^(a[332] & b[272])^(a[331] & b[273])^(a[330] & b[274])^(a[329] & b[275])^(a[328] & b[276])^(a[327] & b[277])^(a[326] & b[278])^(a[325] & b[279])^(a[324] & b[280])^(a[323] & b[281])^(a[322] & b[282])^(a[321] & b[283])^(a[320] & b[284])^(a[319] & b[285])^(a[318] & b[286])^(a[317] & b[287])^(a[316] & b[288])^(a[315] & b[289])^(a[314] & b[290])^(a[313] & b[291])^(a[312] & b[292])^(a[311] & b[293])^(a[310] & b[294])^(a[309] & b[295])^(a[308] & b[296])^(a[307] & b[297])^(a[306] & b[298])^(a[305] & b[299])^(a[304] & b[300])^(a[303] & b[301])^(a[302] & b[302])^(a[301] & b[303])^(a[300] & b[304])^(a[299] & b[305])^(a[298] & b[306])^(a[297] & b[307])^(a[296] & b[308])^(a[295] & b[309])^(a[294] & b[310])^(a[293] & b[311])^(a[292] & b[312])^(a[291] & b[313])^(a[290] & b[314])^(a[289] & b[315])^(a[288] & b[316])^(a[287] & b[317])^(a[286] & b[318])^(a[285] & b[319])^(a[284] & b[320])^(a[283] & b[321])^(a[282] & b[322])^(a[281] & b[323])^(a[280] & b[324])^(a[279] & b[325])^(a[278] & b[326])^(a[277] & b[327])^(a[276] & b[328])^(a[275] & b[329])^(a[274] & b[330])^(a[273] & b[331])^(a[272] & b[332])^(a[271] & b[333])^(a[270] & b[334])^(a[269] & b[335])^(a[268] & b[336])^(a[267] & b[337])^(a[266] & b[338])^(a[265] & b[339])^(a[264] & b[340])^(a[263] & b[341])^(a[262] & b[342])^(a[261] & b[343])^(a[260] & b[344])^(a[259] & b[345])^(a[258] & b[346])^(a[257] & b[347])^(a[256] & b[348])^(a[255] & b[349])^(a[254] & b[350])^(a[253] & b[351])^(a[252] & b[352])^(a[251] & b[353])^(a[250] & b[354])^(a[249] & b[355])^(a[248] & b[356])^(a[247] & b[357])^(a[246] & b[358])^(a[245] & b[359])^(a[244] & b[360])^(a[243] & b[361])^(a[242] & b[362])^(a[241] & b[363])^(a[240] & b[364])^(a[239] & b[365])^(a[238] & b[366])^(a[237] & b[367])^(a[236] & b[368])^(a[235] & b[369])^(a[234] & b[370])^(a[233] & b[371])^(a[232] & b[372])^(a[231] & b[373])^(a[230] & b[374])^(a[229] & b[375])^(a[228] & b[376])^(a[227] & b[377])^(a[226] & b[378])^(a[225] & b[379])^(a[224] & b[380])^(a[223] & b[381])^(a[222] & b[382])^(a[221] & b[383])^(a[220] & b[384])^(a[219] & b[385])^(a[218] & b[386])^(a[217] & b[387])^(a[216] & b[388])^(a[215] & b[389])^(a[214] & b[390])^(a[213] & b[391])^(a[212] & b[392])^(a[211] & b[393])^(a[210] & b[394])^(a[209] & b[395])^(a[208] & b[396])^(a[207] & b[397])^(a[206] & b[398])^(a[205] & b[399])^(a[204] & b[400])^(a[203] & b[401])^(a[202] & b[402])^(a[201] & b[403])^(a[200] & b[404])^(a[199] & b[405])^(a[198] & b[406])^(a[197] & b[407])^(a[196] & b[408]);
assign y[605] = (a[408] & b[197])^(a[407] & b[198])^(a[406] & b[199])^(a[405] & b[200])^(a[404] & b[201])^(a[403] & b[202])^(a[402] & b[203])^(a[401] & b[204])^(a[400] & b[205])^(a[399] & b[206])^(a[398] & b[207])^(a[397] & b[208])^(a[396] & b[209])^(a[395] & b[210])^(a[394] & b[211])^(a[393] & b[212])^(a[392] & b[213])^(a[391] & b[214])^(a[390] & b[215])^(a[389] & b[216])^(a[388] & b[217])^(a[387] & b[218])^(a[386] & b[219])^(a[385] & b[220])^(a[384] & b[221])^(a[383] & b[222])^(a[382] & b[223])^(a[381] & b[224])^(a[380] & b[225])^(a[379] & b[226])^(a[378] & b[227])^(a[377] & b[228])^(a[376] & b[229])^(a[375] & b[230])^(a[374] & b[231])^(a[373] & b[232])^(a[372] & b[233])^(a[371] & b[234])^(a[370] & b[235])^(a[369] & b[236])^(a[368] & b[237])^(a[367] & b[238])^(a[366] & b[239])^(a[365] & b[240])^(a[364] & b[241])^(a[363] & b[242])^(a[362] & b[243])^(a[361] & b[244])^(a[360] & b[245])^(a[359] & b[246])^(a[358] & b[247])^(a[357] & b[248])^(a[356] & b[249])^(a[355] & b[250])^(a[354] & b[251])^(a[353] & b[252])^(a[352] & b[253])^(a[351] & b[254])^(a[350] & b[255])^(a[349] & b[256])^(a[348] & b[257])^(a[347] & b[258])^(a[346] & b[259])^(a[345] & b[260])^(a[344] & b[261])^(a[343] & b[262])^(a[342] & b[263])^(a[341] & b[264])^(a[340] & b[265])^(a[339] & b[266])^(a[338] & b[267])^(a[337] & b[268])^(a[336] & b[269])^(a[335] & b[270])^(a[334] & b[271])^(a[333] & b[272])^(a[332] & b[273])^(a[331] & b[274])^(a[330] & b[275])^(a[329] & b[276])^(a[328] & b[277])^(a[327] & b[278])^(a[326] & b[279])^(a[325] & b[280])^(a[324] & b[281])^(a[323] & b[282])^(a[322] & b[283])^(a[321] & b[284])^(a[320] & b[285])^(a[319] & b[286])^(a[318] & b[287])^(a[317] & b[288])^(a[316] & b[289])^(a[315] & b[290])^(a[314] & b[291])^(a[313] & b[292])^(a[312] & b[293])^(a[311] & b[294])^(a[310] & b[295])^(a[309] & b[296])^(a[308] & b[297])^(a[307] & b[298])^(a[306] & b[299])^(a[305] & b[300])^(a[304] & b[301])^(a[303] & b[302])^(a[302] & b[303])^(a[301] & b[304])^(a[300] & b[305])^(a[299] & b[306])^(a[298] & b[307])^(a[297] & b[308])^(a[296] & b[309])^(a[295] & b[310])^(a[294] & b[311])^(a[293] & b[312])^(a[292] & b[313])^(a[291] & b[314])^(a[290] & b[315])^(a[289] & b[316])^(a[288] & b[317])^(a[287] & b[318])^(a[286] & b[319])^(a[285] & b[320])^(a[284] & b[321])^(a[283] & b[322])^(a[282] & b[323])^(a[281] & b[324])^(a[280] & b[325])^(a[279] & b[326])^(a[278] & b[327])^(a[277] & b[328])^(a[276] & b[329])^(a[275] & b[330])^(a[274] & b[331])^(a[273] & b[332])^(a[272] & b[333])^(a[271] & b[334])^(a[270] & b[335])^(a[269] & b[336])^(a[268] & b[337])^(a[267] & b[338])^(a[266] & b[339])^(a[265] & b[340])^(a[264] & b[341])^(a[263] & b[342])^(a[262] & b[343])^(a[261] & b[344])^(a[260] & b[345])^(a[259] & b[346])^(a[258] & b[347])^(a[257] & b[348])^(a[256] & b[349])^(a[255] & b[350])^(a[254] & b[351])^(a[253] & b[352])^(a[252] & b[353])^(a[251] & b[354])^(a[250] & b[355])^(a[249] & b[356])^(a[248] & b[357])^(a[247] & b[358])^(a[246] & b[359])^(a[245] & b[360])^(a[244] & b[361])^(a[243] & b[362])^(a[242] & b[363])^(a[241] & b[364])^(a[240] & b[365])^(a[239] & b[366])^(a[238] & b[367])^(a[237] & b[368])^(a[236] & b[369])^(a[235] & b[370])^(a[234] & b[371])^(a[233] & b[372])^(a[232] & b[373])^(a[231] & b[374])^(a[230] & b[375])^(a[229] & b[376])^(a[228] & b[377])^(a[227] & b[378])^(a[226] & b[379])^(a[225] & b[380])^(a[224] & b[381])^(a[223] & b[382])^(a[222] & b[383])^(a[221] & b[384])^(a[220] & b[385])^(a[219] & b[386])^(a[218] & b[387])^(a[217] & b[388])^(a[216] & b[389])^(a[215] & b[390])^(a[214] & b[391])^(a[213] & b[392])^(a[212] & b[393])^(a[211] & b[394])^(a[210] & b[395])^(a[209] & b[396])^(a[208] & b[397])^(a[207] & b[398])^(a[206] & b[399])^(a[205] & b[400])^(a[204] & b[401])^(a[203] & b[402])^(a[202] & b[403])^(a[201] & b[404])^(a[200] & b[405])^(a[199] & b[406])^(a[198] & b[407])^(a[197] & b[408]);
assign y[606] = (a[408] & b[198])^(a[407] & b[199])^(a[406] & b[200])^(a[405] & b[201])^(a[404] & b[202])^(a[403] & b[203])^(a[402] & b[204])^(a[401] & b[205])^(a[400] & b[206])^(a[399] & b[207])^(a[398] & b[208])^(a[397] & b[209])^(a[396] & b[210])^(a[395] & b[211])^(a[394] & b[212])^(a[393] & b[213])^(a[392] & b[214])^(a[391] & b[215])^(a[390] & b[216])^(a[389] & b[217])^(a[388] & b[218])^(a[387] & b[219])^(a[386] & b[220])^(a[385] & b[221])^(a[384] & b[222])^(a[383] & b[223])^(a[382] & b[224])^(a[381] & b[225])^(a[380] & b[226])^(a[379] & b[227])^(a[378] & b[228])^(a[377] & b[229])^(a[376] & b[230])^(a[375] & b[231])^(a[374] & b[232])^(a[373] & b[233])^(a[372] & b[234])^(a[371] & b[235])^(a[370] & b[236])^(a[369] & b[237])^(a[368] & b[238])^(a[367] & b[239])^(a[366] & b[240])^(a[365] & b[241])^(a[364] & b[242])^(a[363] & b[243])^(a[362] & b[244])^(a[361] & b[245])^(a[360] & b[246])^(a[359] & b[247])^(a[358] & b[248])^(a[357] & b[249])^(a[356] & b[250])^(a[355] & b[251])^(a[354] & b[252])^(a[353] & b[253])^(a[352] & b[254])^(a[351] & b[255])^(a[350] & b[256])^(a[349] & b[257])^(a[348] & b[258])^(a[347] & b[259])^(a[346] & b[260])^(a[345] & b[261])^(a[344] & b[262])^(a[343] & b[263])^(a[342] & b[264])^(a[341] & b[265])^(a[340] & b[266])^(a[339] & b[267])^(a[338] & b[268])^(a[337] & b[269])^(a[336] & b[270])^(a[335] & b[271])^(a[334] & b[272])^(a[333] & b[273])^(a[332] & b[274])^(a[331] & b[275])^(a[330] & b[276])^(a[329] & b[277])^(a[328] & b[278])^(a[327] & b[279])^(a[326] & b[280])^(a[325] & b[281])^(a[324] & b[282])^(a[323] & b[283])^(a[322] & b[284])^(a[321] & b[285])^(a[320] & b[286])^(a[319] & b[287])^(a[318] & b[288])^(a[317] & b[289])^(a[316] & b[290])^(a[315] & b[291])^(a[314] & b[292])^(a[313] & b[293])^(a[312] & b[294])^(a[311] & b[295])^(a[310] & b[296])^(a[309] & b[297])^(a[308] & b[298])^(a[307] & b[299])^(a[306] & b[300])^(a[305] & b[301])^(a[304] & b[302])^(a[303] & b[303])^(a[302] & b[304])^(a[301] & b[305])^(a[300] & b[306])^(a[299] & b[307])^(a[298] & b[308])^(a[297] & b[309])^(a[296] & b[310])^(a[295] & b[311])^(a[294] & b[312])^(a[293] & b[313])^(a[292] & b[314])^(a[291] & b[315])^(a[290] & b[316])^(a[289] & b[317])^(a[288] & b[318])^(a[287] & b[319])^(a[286] & b[320])^(a[285] & b[321])^(a[284] & b[322])^(a[283] & b[323])^(a[282] & b[324])^(a[281] & b[325])^(a[280] & b[326])^(a[279] & b[327])^(a[278] & b[328])^(a[277] & b[329])^(a[276] & b[330])^(a[275] & b[331])^(a[274] & b[332])^(a[273] & b[333])^(a[272] & b[334])^(a[271] & b[335])^(a[270] & b[336])^(a[269] & b[337])^(a[268] & b[338])^(a[267] & b[339])^(a[266] & b[340])^(a[265] & b[341])^(a[264] & b[342])^(a[263] & b[343])^(a[262] & b[344])^(a[261] & b[345])^(a[260] & b[346])^(a[259] & b[347])^(a[258] & b[348])^(a[257] & b[349])^(a[256] & b[350])^(a[255] & b[351])^(a[254] & b[352])^(a[253] & b[353])^(a[252] & b[354])^(a[251] & b[355])^(a[250] & b[356])^(a[249] & b[357])^(a[248] & b[358])^(a[247] & b[359])^(a[246] & b[360])^(a[245] & b[361])^(a[244] & b[362])^(a[243] & b[363])^(a[242] & b[364])^(a[241] & b[365])^(a[240] & b[366])^(a[239] & b[367])^(a[238] & b[368])^(a[237] & b[369])^(a[236] & b[370])^(a[235] & b[371])^(a[234] & b[372])^(a[233] & b[373])^(a[232] & b[374])^(a[231] & b[375])^(a[230] & b[376])^(a[229] & b[377])^(a[228] & b[378])^(a[227] & b[379])^(a[226] & b[380])^(a[225] & b[381])^(a[224] & b[382])^(a[223] & b[383])^(a[222] & b[384])^(a[221] & b[385])^(a[220] & b[386])^(a[219] & b[387])^(a[218] & b[388])^(a[217] & b[389])^(a[216] & b[390])^(a[215] & b[391])^(a[214] & b[392])^(a[213] & b[393])^(a[212] & b[394])^(a[211] & b[395])^(a[210] & b[396])^(a[209] & b[397])^(a[208] & b[398])^(a[207] & b[399])^(a[206] & b[400])^(a[205] & b[401])^(a[204] & b[402])^(a[203] & b[403])^(a[202] & b[404])^(a[201] & b[405])^(a[200] & b[406])^(a[199] & b[407])^(a[198] & b[408]);
assign y[607] = (a[408] & b[199])^(a[407] & b[200])^(a[406] & b[201])^(a[405] & b[202])^(a[404] & b[203])^(a[403] & b[204])^(a[402] & b[205])^(a[401] & b[206])^(a[400] & b[207])^(a[399] & b[208])^(a[398] & b[209])^(a[397] & b[210])^(a[396] & b[211])^(a[395] & b[212])^(a[394] & b[213])^(a[393] & b[214])^(a[392] & b[215])^(a[391] & b[216])^(a[390] & b[217])^(a[389] & b[218])^(a[388] & b[219])^(a[387] & b[220])^(a[386] & b[221])^(a[385] & b[222])^(a[384] & b[223])^(a[383] & b[224])^(a[382] & b[225])^(a[381] & b[226])^(a[380] & b[227])^(a[379] & b[228])^(a[378] & b[229])^(a[377] & b[230])^(a[376] & b[231])^(a[375] & b[232])^(a[374] & b[233])^(a[373] & b[234])^(a[372] & b[235])^(a[371] & b[236])^(a[370] & b[237])^(a[369] & b[238])^(a[368] & b[239])^(a[367] & b[240])^(a[366] & b[241])^(a[365] & b[242])^(a[364] & b[243])^(a[363] & b[244])^(a[362] & b[245])^(a[361] & b[246])^(a[360] & b[247])^(a[359] & b[248])^(a[358] & b[249])^(a[357] & b[250])^(a[356] & b[251])^(a[355] & b[252])^(a[354] & b[253])^(a[353] & b[254])^(a[352] & b[255])^(a[351] & b[256])^(a[350] & b[257])^(a[349] & b[258])^(a[348] & b[259])^(a[347] & b[260])^(a[346] & b[261])^(a[345] & b[262])^(a[344] & b[263])^(a[343] & b[264])^(a[342] & b[265])^(a[341] & b[266])^(a[340] & b[267])^(a[339] & b[268])^(a[338] & b[269])^(a[337] & b[270])^(a[336] & b[271])^(a[335] & b[272])^(a[334] & b[273])^(a[333] & b[274])^(a[332] & b[275])^(a[331] & b[276])^(a[330] & b[277])^(a[329] & b[278])^(a[328] & b[279])^(a[327] & b[280])^(a[326] & b[281])^(a[325] & b[282])^(a[324] & b[283])^(a[323] & b[284])^(a[322] & b[285])^(a[321] & b[286])^(a[320] & b[287])^(a[319] & b[288])^(a[318] & b[289])^(a[317] & b[290])^(a[316] & b[291])^(a[315] & b[292])^(a[314] & b[293])^(a[313] & b[294])^(a[312] & b[295])^(a[311] & b[296])^(a[310] & b[297])^(a[309] & b[298])^(a[308] & b[299])^(a[307] & b[300])^(a[306] & b[301])^(a[305] & b[302])^(a[304] & b[303])^(a[303] & b[304])^(a[302] & b[305])^(a[301] & b[306])^(a[300] & b[307])^(a[299] & b[308])^(a[298] & b[309])^(a[297] & b[310])^(a[296] & b[311])^(a[295] & b[312])^(a[294] & b[313])^(a[293] & b[314])^(a[292] & b[315])^(a[291] & b[316])^(a[290] & b[317])^(a[289] & b[318])^(a[288] & b[319])^(a[287] & b[320])^(a[286] & b[321])^(a[285] & b[322])^(a[284] & b[323])^(a[283] & b[324])^(a[282] & b[325])^(a[281] & b[326])^(a[280] & b[327])^(a[279] & b[328])^(a[278] & b[329])^(a[277] & b[330])^(a[276] & b[331])^(a[275] & b[332])^(a[274] & b[333])^(a[273] & b[334])^(a[272] & b[335])^(a[271] & b[336])^(a[270] & b[337])^(a[269] & b[338])^(a[268] & b[339])^(a[267] & b[340])^(a[266] & b[341])^(a[265] & b[342])^(a[264] & b[343])^(a[263] & b[344])^(a[262] & b[345])^(a[261] & b[346])^(a[260] & b[347])^(a[259] & b[348])^(a[258] & b[349])^(a[257] & b[350])^(a[256] & b[351])^(a[255] & b[352])^(a[254] & b[353])^(a[253] & b[354])^(a[252] & b[355])^(a[251] & b[356])^(a[250] & b[357])^(a[249] & b[358])^(a[248] & b[359])^(a[247] & b[360])^(a[246] & b[361])^(a[245] & b[362])^(a[244] & b[363])^(a[243] & b[364])^(a[242] & b[365])^(a[241] & b[366])^(a[240] & b[367])^(a[239] & b[368])^(a[238] & b[369])^(a[237] & b[370])^(a[236] & b[371])^(a[235] & b[372])^(a[234] & b[373])^(a[233] & b[374])^(a[232] & b[375])^(a[231] & b[376])^(a[230] & b[377])^(a[229] & b[378])^(a[228] & b[379])^(a[227] & b[380])^(a[226] & b[381])^(a[225] & b[382])^(a[224] & b[383])^(a[223] & b[384])^(a[222] & b[385])^(a[221] & b[386])^(a[220] & b[387])^(a[219] & b[388])^(a[218] & b[389])^(a[217] & b[390])^(a[216] & b[391])^(a[215] & b[392])^(a[214] & b[393])^(a[213] & b[394])^(a[212] & b[395])^(a[211] & b[396])^(a[210] & b[397])^(a[209] & b[398])^(a[208] & b[399])^(a[207] & b[400])^(a[206] & b[401])^(a[205] & b[402])^(a[204] & b[403])^(a[203] & b[404])^(a[202] & b[405])^(a[201] & b[406])^(a[200] & b[407])^(a[199] & b[408]);
assign y[608] = (a[408] & b[200])^(a[407] & b[201])^(a[406] & b[202])^(a[405] & b[203])^(a[404] & b[204])^(a[403] & b[205])^(a[402] & b[206])^(a[401] & b[207])^(a[400] & b[208])^(a[399] & b[209])^(a[398] & b[210])^(a[397] & b[211])^(a[396] & b[212])^(a[395] & b[213])^(a[394] & b[214])^(a[393] & b[215])^(a[392] & b[216])^(a[391] & b[217])^(a[390] & b[218])^(a[389] & b[219])^(a[388] & b[220])^(a[387] & b[221])^(a[386] & b[222])^(a[385] & b[223])^(a[384] & b[224])^(a[383] & b[225])^(a[382] & b[226])^(a[381] & b[227])^(a[380] & b[228])^(a[379] & b[229])^(a[378] & b[230])^(a[377] & b[231])^(a[376] & b[232])^(a[375] & b[233])^(a[374] & b[234])^(a[373] & b[235])^(a[372] & b[236])^(a[371] & b[237])^(a[370] & b[238])^(a[369] & b[239])^(a[368] & b[240])^(a[367] & b[241])^(a[366] & b[242])^(a[365] & b[243])^(a[364] & b[244])^(a[363] & b[245])^(a[362] & b[246])^(a[361] & b[247])^(a[360] & b[248])^(a[359] & b[249])^(a[358] & b[250])^(a[357] & b[251])^(a[356] & b[252])^(a[355] & b[253])^(a[354] & b[254])^(a[353] & b[255])^(a[352] & b[256])^(a[351] & b[257])^(a[350] & b[258])^(a[349] & b[259])^(a[348] & b[260])^(a[347] & b[261])^(a[346] & b[262])^(a[345] & b[263])^(a[344] & b[264])^(a[343] & b[265])^(a[342] & b[266])^(a[341] & b[267])^(a[340] & b[268])^(a[339] & b[269])^(a[338] & b[270])^(a[337] & b[271])^(a[336] & b[272])^(a[335] & b[273])^(a[334] & b[274])^(a[333] & b[275])^(a[332] & b[276])^(a[331] & b[277])^(a[330] & b[278])^(a[329] & b[279])^(a[328] & b[280])^(a[327] & b[281])^(a[326] & b[282])^(a[325] & b[283])^(a[324] & b[284])^(a[323] & b[285])^(a[322] & b[286])^(a[321] & b[287])^(a[320] & b[288])^(a[319] & b[289])^(a[318] & b[290])^(a[317] & b[291])^(a[316] & b[292])^(a[315] & b[293])^(a[314] & b[294])^(a[313] & b[295])^(a[312] & b[296])^(a[311] & b[297])^(a[310] & b[298])^(a[309] & b[299])^(a[308] & b[300])^(a[307] & b[301])^(a[306] & b[302])^(a[305] & b[303])^(a[304] & b[304])^(a[303] & b[305])^(a[302] & b[306])^(a[301] & b[307])^(a[300] & b[308])^(a[299] & b[309])^(a[298] & b[310])^(a[297] & b[311])^(a[296] & b[312])^(a[295] & b[313])^(a[294] & b[314])^(a[293] & b[315])^(a[292] & b[316])^(a[291] & b[317])^(a[290] & b[318])^(a[289] & b[319])^(a[288] & b[320])^(a[287] & b[321])^(a[286] & b[322])^(a[285] & b[323])^(a[284] & b[324])^(a[283] & b[325])^(a[282] & b[326])^(a[281] & b[327])^(a[280] & b[328])^(a[279] & b[329])^(a[278] & b[330])^(a[277] & b[331])^(a[276] & b[332])^(a[275] & b[333])^(a[274] & b[334])^(a[273] & b[335])^(a[272] & b[336])^(a[271] & b[337])^(a[270] & b[338])^(a[269] & b[339])^(a[268] & b[340])^(a[267] & b[341])^(a[266] & b[342])^(a[265] & b[343])^(a[264] & b[344])^(a[263] & b[345])^(a[262] & b[346])^(a[261] & b[347])^(a[260] & b[348])^(a[259] & b[349])^(a[258] & b[350])^(a[257] & b[351])^(a[256] & b[352])^(a[255] & b[353])^(a[254] & b[354])^(a[253] & b[355])^(a[252] & b[356])^(a[251] & b[357])^(a[250] & b[358])^(a[249] & b[359])^(a[248] & b[360])^(a[247] & b[361])^(a[246] & b[362])^(a[245] & b[363])^(a[244] & b[364])^(a[243] & b[365])^(a[242] & b[366])^(a[241] & b[367])^(a[240] & b[368])^(a[239] & b[369])^(a[238] & b[370])^(a[237] & b[371])^(a[236] & b[372])^(a[235] & b[373])^(a[234] & b[374])^(a[233] & b[375])^(a[232] & b[376])^(a[231] & b[377])^(a[230] & b[378])^(a[229] & b[379])^(a[228] & b[380])^(a[227] & b[381])^(a[226] & b[382])^(a[225] & b[383])^(a[224] & b[384])^(a[223] & b[385])^(a[222] & b[386])^(a[221] & b[387])^(a[220] & b[388])^(a[219] & b[389])^(a[218] & b[390])^(a[217] & b[391])^(a[216] & b[392])^(a[215] & b[393])^(a[214] & b[394])^(a[213] & b[395])^(a[212] & b[396])^(a[211] & b[397])^(a[210] & b[398])^(a[209] & b[399])^(a[208] & b[400])^(a[207] & b[401])^(a[206] & b[402])^(a[205] & b[403])^(a[204] & b[404])^(a[203] & b[405])^(a[202] & b[406])^(a[201] & b[407])^(a[200] & b[408]);
assign y[609] = (a[408] & b[201])^(a[407] & b[202])^(a[406] & b[203])^(a[405] & b[204])^(a[404] & b[205])^(a[403] & b[206])^(a[402] & b[207])^(a[401] & b[208])^(a[400] & b[209])^(a[399] & b[210])^(a[398] & b[211])^(a[397] & b[212])^(a[396] & b[213])^(a[395] & b[214])^(a[394] & b[215])^(a[393] & b[216])^(a[392] & b[217])^(a[391] & b[218])^(a[390] & b[219])^(a[389] & b[220])^(a[388] & b[221])^(a[387] & b[222])^(a[386] & b[223])^(a[385] & b[224])^(a[384] & b[225])^(a[383] & b[226])^(a[382] & b[227])^(a[381] & b[228])^(a[380] & b[229])^(a[379] & b[230])^(a[378] & b[231])^(a[377] & b[232])^(a[376] & b[233])^(a[375] & b[234])^(a[374] & b[235])^(a[373] & b[236])^(a[372] & b[237])^(a[371] & b[238])^(a[370] & b[239])^(a[369] & b[240])^(a[368] & b[241])^(a[367] & b[242])^(a[366] & b[243])^(a[365] & b[244])^(a[364] & b[245])^(a[363] & b[246])^(a[362] & b[247])^(a[361] & b[248])^(a[360] & b[249])^(a[359] & b[250])^(a[358] & b[251])^(a[357] & b[252])^(a[356] & b[253])^(a[355] & b[254])^(a[354] & b[255])^(a[353] & b[256])^(a[352] & b[257])^(a[351] & b[258])^(a[350] & b[259])^(a[349] & b[260])^(a[348] & b[261])^(a[347] & b[262])^(a[346] & b[263])^(a[345] & b[264])^(a[344] & b[265])^(a[343] & b[266])^(a[342] & b[267])^(a[341] & b[268])^(a[340] & b[269])^(a[339] & b[270])^(a[338] & b[271])^(a[337] & b[272])^(a[336] & b[273])^(a[335] & b[274])^(a[334] & b[275])^(a[333] & b[276])^(a[332] & b[277])^(a[331] & b[278])^(a[330] & b[279])^(a[329] & b[280])^(a[328] & b[281])^(a[327] & b[282])^(a[326] & b[283])^(a[325] & b[284])^(a[324] & b[285])^(a[323] & b[286])^(a[322] & b[287])^(a[321] & b[288])^(a[320] & b[289])^(a[319] & b[290])^(a[318] & b[291])^(a[317] & b[292])^(a[316] & b[293])^(a[315] & b[294])^(a[314] & b[295])^(a[313] & b[296])^(a[312] & b[297])^(a[311] & b[298])^(a[310] & b[299])^(a[309] & b[300])^(a[308] & b[301])^(a[307] & b[302])^(a[306] & b[303])^(a[305] & b[304])^(a[304] & b[305])^(a[303] & b[306])^(a[302] & b[307])^(a[301] & b[308])^(a[300] & b[309])^(a[299] & b[310])^(a[298] & b[311])^(a[297] & b[312])^(a[296] & b[313])^(a[295] & b[314])^(a[294] & b[315])^(a[293] & b[316])^(a[292] & b[317])^(a[291] & b[318])^(a[290] & b[319])^(a[289] & b[320])^(a[288] & b[321])^(a[287] & b[322])^(a[286] & b[323])^(a[285] & b[324])^(a[284] & b[325])^(a[283] & b[326])^(a[282] & b[327])^(a[281] & b[328])^(a[280] & b[329])^(a[279] & b[330])^(a[278] & b[331])^(a[277] & b[332])^(a[276] & b[333])^(a[275] & b[334])^(a[274] & b[335])^(a[273] & b[336])^(a[272] & b[337])^(a[271] & b[338])^(a[270] & b[339])^(a[269] & b[340])^(a[268] & b[341])^(a[267] & b[342])^(a[266] & b[343])^(a[265] & b[344])^(a[264] & b[345])^(a[263] & b[346])^(a[262] & b[347])^(a[261] & b[348])^(a[260] & b[349])^(a[259] & b[350])^(a[258] & b[351])^(a[257] & b[352])^(a[256] & b[353])^(a[255] & b[354])^(a[254] & b[355])^(a[253] & b[356])^(a[252] & b[357])^(a[251] & b[358])^(a[250] & b[359])^(a[249] & b[360])^(a[248] & b[361])^(a[247] & b[362])^(a[246] & b[363])^(a[245] & b[364])^(a[244] & b[365])^(a[243] & b[366])^(a[242] & b[367])^(a[241] & b[368])^(a[240] & b[369])^(a[239] & b[370])^(a[238] & b[371])^(a[237] & b[372])^(a[236] & b[373])^(a[235] & b[374])^(a[234] & b[375])^(a[233] & b[376])^(a[232] & b[377])^(a[231] & b[378])^(a[230] & b[379])^(a[229] & b[380])^(a[228] & b[381])^(a[227] & b[382])^(a[226] & b[383])^(a[225] & b[384])^(a[224] & b[385])^(a[223] & b[386])^(a[222] & b[387])^(a[221] & b[388])^(a[220] & b[389])^(a[219] & b[390])^(a[218] & b[391])^(a[217] & b[392])^(a[216] & b[393])^(a[215] & b[394])^(a[214] & b[395])^(a[213] & b[396])^(a[212] & b[397])^(a[211] & b[398])^(a[210] & b[399])^(a[209] & b[400])^(a[208] & b[401])^(a[207] & b[402])^(a[206] & b[403])^(a[205] & b[404])^(a[204] & b[405])^(a[203] & b[406])^(a[202] & b[407])^(a[201] & b[408]);
assign y[610] = (a[408] & b[202])^(a[407] & b[203])^(a[406] & b[204])^(a[405] & b[205])^(a[404] & b[206])^(a[403] & b[207])^(a[402] & b[208])^(a[401] & b[209])^(a[400] & b[210])^(a[399] & b[211])^(a[398] & b[212])^(a[397] & b[213])^(a[396] & b[214])^(a[395] & b[215])^(a[394] & b[216])^(a[393] & b[217])^(a[392] & b[218])^(a[391] & b[219])^(a[390] & b[220])^(a[389] & b[221])^(a[388] & b[222])^(a[387] & b[223])^(a[386] & b[224])^(a[385] & b[225])^(a[384] & b[226])^(a[383] & b[227])^(a[382] & b[228])^(a[381] & b[229])^(a[380] & b[230])^(a[379] & b[231])^(a[378] & b[232])^(a[377] & b[233])^(a[376] & b[234])^(a[375] & b[235])^(a[374] & b[236])^(a[373] & b[237])^(a[372] & b[238])^(a[371] & b[239])^(a[370] & b[240])^(a[369] & b[241])^(a[368] & b[242])^(a[367] & b[243])^(a[366] & b[244])^(a[365] & b[245])^(a[364] & b[246])^(a[363] & b[247])^(a[362] & b[248])^(a[361] & b[249])^(a[360] & b[250])^(a[359] & b[251])^(a[358] & b[252])^(a[357] & b[253])^(a[356] & b[254])^(a[355] & b[255])^(a[354] & b[256])^(a[353] & b[257])^(a[352] & b[258])^(a[351] & b[259])^(a[350] & b[260])^(a[349] & b[261])^(a[348] & b[262])^(a[347] & b[263])^(a[346] & b[264])^(a[345] & b[265])^(a[344] & b[266])^(a[343] & b[267])^(a[342] & b[268])^(a[341] & b[269])^(a[340] & b[270])^(a[339] & b[271])^(a[338] & b[272])^(a[337] & b[273])^(a[336] & b[274])^(a[335] & b[275])^(a[334] & b[276])^(a[333] & b[277])^(a[332] & b[278])^(a[331] & b[279])^(a[330] & b[280])^(a[329] & b[281])^(a[328] & b[282])^(a[327] & b[283])^(a[326] & b[284])^(a[325] & b[285])^(a[324] & b[286])^(a[323] & b[287])^(a[322] & b[288])^(a[321] & b[289])^(a[320] & b[290])^(a[319] & b[291])^(a[318] & b[292])^(a[317] & b[293])^(a[316] & b[294])^(a[315] & b[295])^(a[314] & b[296])^(a[313] & b[297])^(a[312] & b[298])^(a[311] & b[299])^(a[310] & b[300])^(a[309] & b[301])^(a[308] & b[302])^(a[307] & b[303])^(a[306] & b[304])^(a[305] & b[305])^(a[304] & b[306])^(a[303] & b[307])^(a[302] & b[308])^(a[301] & b[309])^(a[300] & b[310])^(a[299] & b[311])^(a[298] & b[312])^(a[297] & b[313])^(a[296] & b[314])^(a[295] & b[315])^(a[294] & b[316])^(a[293] & b[317])^(a[292] & b[318])^(a[291] & b[319])^(a[290] & b[320])^(a[289] & b[321])^(a[288] & b[322])^(a[287] & b[323])^(a[286] & b[324])^(a[285] & b[325])^(a[284] & b[326])^(a[283] & b[327])^(a[282] & b[328])^(a[281] & b[329])^(a[280] & b[330])^(a[279] & b[331])^(a[278] & b[332])^(a[277] & b[333])^(a[276] & b[334])^(a[275] & b[335])^(a[274] & b[336])^(a[273] & b[337])^(a[272] & b[338])^(a[271] & b[339])^(a[270] & b[340])^(a[269] & b[341])^(a[268] & b[342])^(a[267] & b[343])^(a[266] & b[344])^(a[265] & b[345])^(a[264] & b[346])^(a[263] & b[347])^(a[262] & b[348])^(a[261] & b[349])^(a[260] & b[350])^(a[259] & b[351])^(a[258] & b[352])^(a[257] & b[353])^(a[256] & b[354])^(a[255] & b[355])^(a[254] & b[356])^(a[253] & b[357])^(a[252] & b[358])^(a[251] & b[359])^(a[250] & b[360])^(a[249] & b[361])^(a[248] & b[362])^(a[247] & b[363])^(a[246] & b[364])^(a[245] & b[365])^(a[244] & b[366])^(a[243] & b[367])^(a[242] & b[368])^(a[241] & b[369])^(a[240] & b[370])^(a[239] & b[371])^(a[238] & b[372])^(a[237] & b[373])^(a[236] & b[374])^(a[235] & b[375])^(a[234] & b[376])^(a[233] & b[377])^(a[232] & b[378])^(a[231] & b[379])^(a[230] & b[380])^(a[229] & b[381])^(a[228] & b[382])^(a[227] & b[383])^(a[226] & b[384])^(a[225] & b[385])^(a[224] & b[386])^(a[223] & b[387])^(a[222] & b[388])^(a[221] & b[389])^(a[220] & b[390])^(a[219] & b[391])^(a[218] & b[392])^(a[217] & b[393])^(a[216] & b[394])^(a[215] & b[395])^(a[214] & b[396])^(a[213] & b[397])^(a[212] & b[398])^(a[211] & b[399])^(a[210] & b[400])^(a[209] & b[401])^(a[208] & b[402])^(a[207] & b[403])^(a[206] & b[404])^(a[205] & b[405])^(a[204] & b[406])^(a[203] & b[407])^(a[202] & b[408]);
assign y[611] = (a[408] & b[203])^(a[407] & b[204])^(a[406] & b[205])^(a[405] & b[206])^(a[404] & b[207])^(a[403] & b[208])^(a[402] & b[209])^(a[401] & b[210])^(a[400] & b[211])^(a[399] & b[212])^(a[398] & b[213])^(a[397] & b[214])^(a[396] & b[215])^(a[395] & b[216])^(a[394] & b[217])^(a[393] & b[218])^(a[392] & b[219])^(a[391] & b[220])^(a[390] & b[221])^(a[389] & b[222])^(a[388] & b[223])^(a[387] & b[224])^(a[386] & b[225])^(a[385] & b[226])^(a[384] & b[227])^(a[383] & b[228])^(a[382] & b[229])^(a[381] & b[230])^(a[380] & b[231])^(a[379] & b[232])^(a[378] & b[233])^(a[377] & b[234])^(a[376] & b[235])^(a[375] & b[236])^(a[374] & b[237])^(a[373] & b[238])^(a[372] & b[239])^(a[371] & b[240])^(a[370] & b[241])^(a[369] & b[242])^(a[368] & b[243])^(a[367] & b[244])^(a[366] & b[245])^(a[365] & b[246])^(a[364] & b[247])^(a[363] & b[248])^(a[362] & b[249])^(a[361] & b[250])^(a[360] & b[251])^(a[359] & b[252])^(a[358] & b[253])^(a[357] & b[254])^(a[356] & b[255])^(a[355] & b[256])^(a[354] & b[257])^(a[353] & b[258])^(a[352] & b[259])^(a[351] & b[260])^(a[350] & b[261])^(a[349] & b[262])^(a[348] & b[263])^(a[347] & b[264])^(a[346] & b[265])^(a[345] & b[266])^(a[344] & b[267])^(a[343] & b[268])^(a[342] & b[269])^(a[341] & b[270])^(a[340] & b[271])^(a[339] & b[272])^(a[338] & b[273])^(a[337] & b[274])^(a[336] & b[275])^(a[335] & b[276])^(a[334] & b[277])^(a[333] & b[278])^(a[332] & b[279])^(a[331] & b[280])^(a[330] & b[281])^(a[329] & b[282])^(a[328] & b[283])^(a[327] & b[284])^(a[326] & b[285])^(a[325] & b[286])^(a[324] & b[287])^(a[323] & b[288])^(a[322] & b[289])^(a[321] & b[290])^(a[320] & b[291])^(a[319] & b[292])^(a[318] & b[293])^(a[317] & b[294])^(a[316] & b[295])^(a[315] & b[296])^(a[314] & b[297])^(a[313] & b[298])^(a[312] & b[299])^(a[311] & b[300])^(a[310] & b[301])^(a[309] & b[302])^(a[308] & b[303])^(a[307] & b[304])^(a[306] & b[305])^(a[305] & b[306])^(a[304] & b[307])^(a[303] & b[308])^(a[302] & b[309])^(a[301] & b[310])^(a[300] & b[311])^(a[299] & b[312])^(a[298] & b[313])^(a[297] & b[314])^(a[296] & b[315])^(a[295] & b[316])^(a[294] & b[317])^(a[293] & b[318])^(a[292] & b[319])^(a[291] & b[320])^(a[290] & b[321])^(a[289] & b[322])^(a[288] & b[323])^(a[287] & b[324])^(a[286] & b[325])^(a[285] & b[326])^(a[284] & b[327])^(a[283] & b[328])^(a[282] & b[329])^(a[281] & b[330])^(a[280] & b[331])^(a[279] & b[332])^(a[278] & b[333])^(a[277] & b[334])^(a[276] & b[335])^(a[275] & b[336])^(a[274] & b[337])^(a[273] & b[338])^(a[272] & b[339])^(a[271] & b[340])^(a[270] & b[341])^(a[269] & b[342])^(a[268] & b[343])^(a[267] & b[344])^(a[266] & b[345])^(a[265] & b[346])^(a[264] & b[347])^(a[263] & b[348])^(a[262] & b[349])^(a[261] & b[350])^(a[260] & b[351])^(a[259] & b[352])^(a[258] & b[353])^(a[257] & b[354])^(a[256] & b[355])^(a[255] & b[356])^(a[254] & b[357])^(a[253] & b[358])^(a[252] & b[359])^(a[251] & b[360])^(a[250] & b[361])^(a[249] & b[362])^(a[248] & b[363])^(a[247] & b[364])^(a[246] & b[365])^(a[245] & b[366])^(a[244] & b[367])^(a[243] & b[368])^(a[242] & b[369])^(a[241] & b[370])^(a[240] & b[371])^(a[239] & b[372])^(a[238] & b[373])^(a[237] & b[374])^(a[236] & b[375])^(a[235] & b[376])^(a[234] & b[377])^(a[233] & b[378])^(a[232] & b[379])^(a[231] & b[380])^(a[230] & b[381])^(a[229] & b[382])^(a[228] & b[383])^(a[227] & b[384])^(a[226] & b[385])^(a[225] & b[386])^(a[224] & b[387])^(a[223] & b[388])^(a[222] & b[389])^(a[221] & b[390])^(a[220] & b[391])^(a[219] & b[392])^(a[218] & b[393])^(a[217] & b[394])^(a[216] & b[395])^(a[215] & b[396])^(a[214] & b[397])^(a[213] & b[398])^(a[212] & b[399])^(a[211] & b[400])^(a[210] & b[401])^(a[209] & b[402])^(a[208] & b[403])^(a[207] & b[404])^(a[206] & b[405])^(a[205] & b[406])^(a[204] & b[407])^(a[203] & b[408]);
assign y[612] = (a[408] & b[204])^(a[407] & b[205])^(a[406] & b[206])^(a[405] & b[207])^(a[404] & b[208])^(a[403] & b[209])^(a[402] & b[210])^(a[401] & b[211])^(a[400] & b[212])^(a[399] & b[213])^(a[398] & b[214])^(a[397] & b[215])^(a[396] & b[216])^(a[395] & b[217])^(a[394] & b[218])^(a[393] & b[219])^(a[392] & b[220])^(a[391] & b[221])^(a[390] & b[222])^(a[389] & b[223])^(a[388] & b[224])^(a[387] & b[225])^(a[386] & b[226])^(a[385] & b[227])^(a[384] & b[228])^(a[383] & b[229])^(a[382] & b[230])^(a[381] & b[231])^(a[380] & b[232])^(a[379] & b[233])^(a[378] & b[234])^(a[377] & b[235])^(a[376] & b[236])^(a[375] & b[237])^(a[374] & b[238])^(a[373] & b[239])^(a[372] & b[240])^(a[371] & b[241])^(a[370] & b[242])^(a[369] & b[243])^(a[368] & b[244])^(a[367] & b[245])^(a[366] & b[246])^(a[365] & b[247])^(a[364] & b[248])^(a[363] & b[249])^(a[362] & b[250])^(a[361] & b[251])^(a[360] & b[252])^(a[359] & b[253])^(a[358] & b[254])^(a[357] & b[255])^(a[356] & b[256])^(a[355] & b[257])^(a[354] & b[258])^(a[353] & b[259])^(a[352] & b[260])^(a[351] & b[261])^(a[350] & b[262])^(a[349] & b[263])^(a[348] & b[264])^(a[347] & b[265])^(a[346] & b[266])^(a[345] & b[267])^(a[344] & b[268])^(a[343] & b[269])^(a[342] & b[270])^(a[341] & b[271])^(a[340] & b[272])^(a[339] & b[273])^(a[338] & b[274])^(a[337] & b[275])^(a[336] & b[276])^(a[335] & b[277])^(a[334] & b[278])^(a[333] & b[279])^(a[332] & b[280])^(a[331] & b[281])^(a[330] & b[282])^(a[329] & b[283])^(a[328] & b[284])^(a[327] & b[285])^(a[326] & b[286])^(a[325] & b[287])^(a[324] & b[288])^(a[323] & b[289])^(a[322] & b[290])^(a[321] & b[291])^(a[320] & b[292])^(a[319] & b[293])^(a[318] & b[294])^(a[317] & b[295])^(a[316] & b[296])^(a[315] & b[297])^(a[314] & b[298])^(a[313] & b[299])^(a[312] & b[300])^(a[311] & b[301])^(a[310] & b[302])^(a[309] & b[303])^(a[308] & b[304])^(a[307] & b[305])^(a[306] & b[306])^(a[305] & b[307])^(a[304] & b[308])^(a[303] & b[309])^(a[302] & b[310])^(a[301] & b[311])^(a[300] & b[312])^(a[299] & b[313])^(a[298] & b[314])^(a[297] & b[315])^(a[296] & b[316])^(a[295] & b[317])^(a[294] & b[318])^(a[293] & b[319])^(a[292] & b[320])^(a[291] & b[321])^(a[290] & b[322])^(a[289] & b[323])^(a[288] & b[324])^(a[287] & b[325])^(a[286] & b[326])^(a[285] & b[327])^(a[284] & b[328])^(a[283] & b[329])^(a[282] & b[330])^(a[281] & b[331])^(a[280] & b[332])^(a[279] & b[333])^(a[278] & b[334])^(a[277] & b[335])^(a[276] & b[336])^(a[275] & b[337])^(a[274] & b[338])^(a[273] & b[339])^(a[272] & b[340])^(a[271] & b[341])^(a[270] & b[342])^(a[269] & b[343])^(a[268] & b[344])^(a[267] & b[345])^(a[266] & b[346])^(a[265] & b[347])^(a[264] & b[348])^(a[263] & b[349])^(a[262] & b[350])^(a[261] & b[351])^(a[260] & b[352])^(a[259] & b[353])^(a[258] & b[354])^(a[257] & b[355])^(a[256] & b[356])^(a[255] & b[357])^(a[254] & b[358])^(a[253] & b[359])^(a[252] & b[360])^(a[251] & b[361])^(a[250] & b[362])^(a[249] & b[363])^(a[248] & b[364])^(a[247] & b[365])^(a[246] & b[366])^(a[245] & b[367])^(a[244] & b[368])^(a[243] & b[369])^(a[242] & b[370])^(a[241] & b[371])^(a[240] & b[372])^(a[239] & b[373])^(a[238] & b[374])^(a[237] & b[375])^(a[236] & b[376])^(a[235] & b[377])^(a[234] & b[378])^(a[233] & b[379])^(a[232] & b[380])^(a[231] & b[381])^(a[230] & b[382])^(a[229] & b[383])^(a[228] & b[384])^(a[227] & b[385])^(a[226] & b[386])^(a[225] & b[387])^(a[224] & b[388])^(a[223] & b[389])^(a[222] & b[390])^(a[221] & b[391])^(a[220] & b[392])^(a[219] & b[393])^(a[218] & b[394])^(a[217] & b[395])^(a[216] & b[396])^(a[215] & b[397])^(a[214] & b[398])^(a[213] & b[399])^(a[212] & b[400])^(a[211] & b[401])^(a[210] & b[402])^(a[209] & b[403])^(a[208] & b[404])^(a[207] & b[405])^(a[206] & b[406])^(a[205] & b[407])^(a[204] & b[408]);
assign y[613] = (a[408] & b[205])^(a[407] & b[206])^(a[406] & b[207])^(a[405] & b[208])^(a[404] & b[209])^(a[403] & b[210])^(a[402] & b[211])^(a[401] & b[212])^(a[400] & b[213])^(a[399] & b[214])^(a[398] & b[215])^(a[397] & b[216])^(a[396] & b[217])^(a[395] & b[218])^(a[394] & b[219])^(a[393] & b[220])^(a[392] & b[221])^(a[391] & b[222])^(a[390] & b[223])^(a[389] & b[224])^(a[388] & b[225])^(a[387] & b[226])^(a[386] & b[227])^(a[385] & b[228])^(a[384] & b[229])^(a[383] & b[230])^(a[382] & b[231])^(a[381] & b[232])^(a[380] & b[233])^(a[379] & b[234])^(a[378] & b[235])^(a[377] & b[236])^(a[376] & b[237])^(a[375] & b[238])^(a[374] & b[239])^(a[373] & b[240])^(a[372] & b[241])^(a[371] & b[242])^(a[370] & b[243])^(a[369] & b[244])^(a[368] & b[245])^(a[367] & b[246])^(a[366] & b[247])^(a[365] & b[248])^(a[364] & b[249])^(a[363] & b[250])^(a[362] & b[251])^(a[361] & b[252])^(a[360] & b[253])^(a[359] & b[254])^(a[358] & b[255])^(a[357] & b[256])^(a[356] & b[257])^(a[355] & b[258])^(a[354] & b[259])^(a[353] & b[260])^(a[352] & b[261])^(a[351] & b[262])^(a[350] & b[263])^(a[349] & b[264])^(a[348] & b[265])^(a[347] & b[266])^(a[346] & b[267])^(a[345] & b[268])^(a[344] & b[269])^(a[343] & b[270])^(a[342] & b[271])^(a[341] & b[272])^(a[340] & b[273])^(a[339] & b[274])^(a[338] & b[275])^(a[337] & b[276])^(a[336] & b[277])^(a[335] & b[278])^(a[334] & b[279])^(a[333] & b[280])^(a[332] & b[281])^(a[331] & b[282])^(a[330] & b[283])^(a[329] & b[284])^(a[328] & b[285])^(a[327] & b[286])^(a[326] & b[287])^(a[325] & b[288])^(a[324] & b[289])^(a[323] & b[290])^(a[322] & b[291])^(a[321] & b[292])^(a[320] & b[293])^(a[319] & b[294])^(a[318] & b[295])^(a[317] & b[296])^(a[316] & b[297])^(a[315] & b[298])^(a[314] & b[299])^(a[313] & b[300])^(a[312] & b[301])^(a[311] & b[302])^(a[310] & b[303])^(a[309] & b[304])^(a[308] & b[305])^(a[307] & b[306])^(a[306] & b[307])^(a[305] & b[308])^(a[304] & b[309])^(a[303] & b[310])^(a[302] & b[311])^(a[301] & b[312])^(a[300] & b[313])^(a[299] & b[314])^(a[298] & b[315])^(a[297] & b[316])^(a[296] & b[317])^(a[295] & b[318])^(a[294] & b[319])^(a[293] & b[320])^(a[292] & b[321])^(a[291] & b[322])^(a[290] & b[323])^(a[289] & b[324])^(a[288] & b[325])^(a[287] & b[326])^(a[286] & b[327])^(a[285] & b[328])^(a[284] & b[329])^(a[283] & b[330])^(a[282] & b[331])^(a[281] & b[332])^(a[280] & b[333])^(a[279] & b[334])^(a[278] & b[335])^(a[277] & b[336])^(a[276] & b[337])^(a[275] & b[338])^(a[274] & b[339])^(a[273] & b[340])^(a[272] & b[341])^(a[271] & b[342])^(a[270] & b[343])^(a[269] & b[344])^(a[268] & b[345])^(a[267] & b[346])^(a[266] & b[347])^(a[265] & b[348])^(a[264] & b[349])^(a[263] & b[350])^(a[262] & b[351])^(a[261] & b[352])^(a[260] & b[353])^(a[259] & b[354])^(a[258] & b[355])^(a[257] & b[356])^(a[256] & b[357])^(a[255] & b[358])^(a[254] & b[359])^(a[253] & b[360])^(a[252] & b[361])^(a[251] & b[362])^(a[250] & b[363])^(a[249] & b[364])^(a[248] & b[365])^(a[247] & b[366])^(a[246] & b[367])^(a[245] & b[368])^(a[244] & b[369])^(a[243] & b[370])^(a[242] & b[371])^(a[241] & b[372])^(a[240] & b[373])^(a[239] & b[374])^(a[238] & b[375])^(a[237] & b[376])^(a[236] & b[377])^(a[235] & b[378])^(a[234] & b[379])^(a[233] & b[380])^(a[232] & b[381])^(a[231] & b[382])^(a[230] & b[383])^(a[229] & b[384])^(a[228] & b[385])^(a[227] & b[386])^(a[226] & b[387])^(a[225] & b[388])^(a[224] & b[389])^(a[223] & b[390])^(a[222] & b[391])^(a[221] & b[392])^(a[220] & b[393])^(a[219] & b[394])^(a[218] & b[395])^(a[217] & b[396])^(a[216] & b[397])^(a[215] & b[398])^(a[214] & b[399])^(a[213] & b[400])^(a[212] & b[401])^(a[211] & b[402])^(a[210] & b[403])^(a[209] & b[404])^(a[208] & b[405])^(a[207] & b[406])^(a[206] & b[407])^(a[205] & b[408]);
assign y[614] = (a[408] & b[206])^(a[407] & b[207])^(a[406] & b[208])^(a[405] & b[209])^(a[404] & b[210])^(a[403] & b[211])^(a[402] & b[212])^(a[401] & b[213])^(a[400] & b[214])^(a[399] & b[215])^(a[398] & b[216])^(a[397] & b[217])^(a[396] & b[218])^(a[395] & b[219])^(a[394] & b[220])^(a[393] & b[221])^(a[392] & b[222])^(a[391] & b[223])^(a[390] & b[224])^(a[389] & b[225])^(a[388] & b[226])^(a[387] & b[227])^(a[386] & b[228])^(a[385] & b[229])^(a[384] & b[230])^(a[383] & b[231])^(a[382] & b[232])^(a[381] & b[233])^(a[380] & b[234])^(a[379] & b[235])^(a[378] & b[236])^(a[377] & b[237])^(a[376] & b[238])^(a[375] & b[239])^(a[374] & b[240])^(a[373] & b[241])^(a[372] & b[242])^(a[371] & b[243])^(a[370] & b[244])^(a[369] & b[245])^(a[368] & b[246])^(a[367] & b[247])^(a[366] & b[248])^(a[365] & b[249])^(a[364] & b[250])^(a[363] & b[251])^(a[362] & b[252])^(a[361] & b[253])^(a[360] & b[254])^(a[359] & b[255])^(a[358] & b[256])^(a[357] & b[257])^(a[356] & b[258])^(a[355] & b[259])^(a[354] & b[260])^(a[353] & b[261])^(a[352] & b[262])^(a[351] & b[263])^(a[350] & b[264])^(a[349] & b[265])^(a[348] & b[266])^(a[347] & b[267])^(a[346] & b[268])^(a[345] & b[269])^(a[344] & b[270])^(a[343] & b[271])^(a[342] & b[272])^(a[341] & b[273])^(a[340] & b[274])^(a[339] & b[275])^(a[338] & b[276])^(a[337] & b[277])^(a[336] & b[278])^(a[335] & b[279])^(a[334] & b[280])^(a[333] & b[281])^(a[332] & b[282])^(a[331] & b[283])^(a[330] & b[284])^(a[329] & b[285])^(a[328] & b[286])^(a[327] & b[287])^(a[326] & b[288])^(a[325] & b[289])^(a[324] & b[290])^(a[323] & b[291])^(a[322] & b[292])^(a[321] & b[293])^(a[320] & b[294])^(a[319] & b[295])^(a[318] & b[296])^(a[317] & b[297])^(a[316] & b[298])^(a[315] & b[299])^(a[314] & b[300])^(a[313] & b[301])^(a[312] & b[302])^(a[311] & b[303])^(a[310] & b[304])^(a[309] & b[305])^(a[308] & b[306])^(a[307] & b[307])^(a[306] & b[308])^(a[305] & b[309])^(a[304] & b[310])^(a[303] & b[311])^(a[302] & b[312])^(a[301] & b[313])^(a[300] & b[314])^(a[299] & b[315])^(a[298] & b[316])^(a[297] & b[317])^(a[296] & b[318])^(a[295] & b[319])^(a[294] & b[320])^(a[293] & b[321])^(a[292] & b[322])^(a[291] & b[323])^(a[290] & b[324])^(a[289] & b[325])^(a[288] & b[326])^(a[287] & b[327])^(a[286] & b[328])^(a[285] & b[329])^(a[284] & b[330])^(a[283] & b[331])^(a[282] & b[332])^(a[281] & b[333])^(a[280] & b[334])^(a[279] & b[335])^(a[278] & b[336])^(a[277] & b[337])^(a[276] & b[338])^(a[275] & b[339])^(a[274] & b[340])^(a[273] & b[341])^(a[272] & b[342])^(a[271] & b[343])^(a[270] & b[344])^(a[269] & b[345])^(a[268] & b[346])^(a[267] & b[347])^(a[266] & b[348])^(a[265] & b[349])^(a[264] & b[350])^(a[263] & b[351])^(a[262] & b[352])^(a[261] & b[353])^(a[260] & b[354])^(a[259] & b[355])^(a[258] & b[356])^(a[257] & b[357])^(a[256] & b[358])^(a[255] & b[359])^(a[254] & b[360])^(a[253] & b[361])^(a[252] & b[362])^(a[251] & b[363])^(a[250] & b[364])^(a[249] & b[365])^(a[248] & b[366])^(a[247] & b[367])^(a[246] & b[368])^(a[245] & b[369])^(a[244] & b[370])^(a[243] & b[371])^(a[242] & b[372])^(a[241] & b[373])^(a[240] & b[374])^(a[239] & b[375])^(a[238] & b[376])^(a[237] & b[377])^(a[236] & b[378])^(a[235] & b[379])^(a[234] & b[380])^(a[233] & b[381])^(a[232] & b[382])^(a[231] & b[383])^(a[230] & b[384])^(a[229] & b[385])^(a[228] & b[386])^(a[227] & b[387])^(a[226] & b[388])^(a[225] & b[389])^(a[224] & b[390])^(a[223] & b[391])^(a[222] & b[392])^(a[221] & b[393])^(a[220] & b[394])^(a[219] & b[395])^(a[218] & b[396])^(a[217] & b[397])^(a[216] & b[398])^(a[215] & b[399])^(a[214] & b[400])^(a[213] & b[401])^(a[212] & b[402])^(a[211] & b[403])^(a[210] & b[404])^(a[209] & b[405])^(a[208] & b[406])^(a[207] & b[407])^(a[206] & b[408]);
assign y[615] = (a[408] & b[207])^(a[407] & b[208])^(a[406] & b[209])^(a[405] & b[210])^(a[404] & b[211])^(a[403] & b[212])^(a[402] & b[213])^(a[401] & b[214])^(a[400] & b[215])^(a[399] & b[216])^(a[398] & b[217])^(a[397] & b[218])^(a[396] & b[219])^(a[395] & b[220])^(a[394] & b[221])^(a[393] & b[222])^(a[392] & b[223])^(a[391] & b[224])^(a[390] & b[225])^(a[389] & b[226])^(a[388] & b[227])^(a[387] & b[228])^(a[386] & b[229])^(a[385] & b[230])^(a[384] & b[231])^(a[383] & b[232])^(a[382] & b[233])^(a[381] & b[234])^(a[380] & b[235])^(a[379] & b[236])^(a[378] & b[237])^(a[377] & b[238])^(a[376] & b[239])^(a[375] & b[240])^(a[374] & b[241])^(a[373] & b[242])^(a[372] & b[243])^(a[371] & b[244])^(a[370] & b[245])^(a[369] & b[246])^(a[368] & b[247])^(a[367] & b[248])^(a[366] & b[249])^(a[365] & b[250])^(a[364] & b[251])^(a[363] & b[252])^(a[362] & b[253])^(a[361] & b[254])^(a[360] & b[255])^(a[359] & b[256])^(a[358] & b[257])^(a[357] & b[258])^(a[356] & b[259])^(a[355] & b[260])^(a[354] & b[261])^(a[353] & b[262])^(a[352] & b[263])^(a[351] & b[264])^(a[350] & b[265])^(a[349] & b[266])^(a[348] & b[267])^(a[347] & b[268])^(a[346] & b[269])^(a[345] & b[270])^(a[344] & b[271])^(a[343] & b[272])^(a[342] & b[273])^(a[341] & b[274])^(a[340] & b[275])^(a[339] & b[276])^(a[338] & b[277])^(a[337] & b[278])^(a[336] & b[279])^(a[335] & b[280])^(a[334] & b[281])^(a[333] & b[282])^(a[332] & b[283])^(a[331] & b[284])^(a[330] & b[285])^(a[329] & b[286])^(a[328] & b[287])^(a[327] & b[288])^(a[326] & b[289])^(a[325] & b[290])^(a[324] & b[291])^(a[323] & b[292])^(a[322] & b[293])^(a[321] & b[294])^(a[320] & b[295])^(a[319] & b[296])^(a[318] & b[297])^(a[317] & b[298])^(a[316] & b[299])^(a[315] & b[300])^(a[314] & b[301])^(a[313] & b[302])^(a[312] & b[303])^(a[311] & b[304])^(a[310] & b[305])^(a[309] & b[306])^(a[308] & b[307])^(a[307] & b[308])^(a[306] & b[309])^(a[305] & b[310])^(a[304] & b[311])^(a[303] & b[312])^(a[302] & b[313])^(a[301] & b[314])^(a[300] & b[315])^(a[299] & b[316])^(a[298] & b[317])^(a[297] & b[318])^(a[296] & b[319])^(a[295] & b[320])^(a[294] & b[321])^(a[293] & b[322])^(a[292] & b[323])^(a[291] & b[324])^(a[290] & b[325])^(a[289] & b[326])^(a[288] & b[327])^(a[287] & b[328])^(a[286] & b[329])^(a[285] & b[330])^(a[284] & b[331])^(a[283] & b[332])^(a[282] & b[333])^(a[281] & b[334])^(a[280] & b[335])^(a[279] & b[336])^(a[278] & b[337])^(a[277] & b[338])^(a[276] & b[339])^(a[275] & b[340])^(a[274] & b[341])^(a[273] & b[342])^(a[272] & b[343])^(a[271] & b[344])^(a[270] & b[345])^(a[269] & b[346])^(a[268] & b[347])^(a[267] & b[348])^(a[266] & b[349])^(a[265] & b[350])^(a[264] & b[351])^(a[263] & b[352])^(a[262] & b[353])^(a[261] & b[354])^(a[260] & b[355])^(a[259] & b[356])^(a[258] & b[357])^(a[257] & b[358])^(a[256] & b[359])^(a[255] & b[360])^(a[254] & b[361])^(a[253] & b[362])^(a[252] & b[363])^(a[251] & b[364])^(a[250] & b[365])^(a[249] & b[366])^(a[248] & b[367])^(a[247] & b[368])^(a[246] & b[369])^(a[245] & b[370])^(a[244] & b[371])^(a[243] & b[372])^(a[242] & b[373])^(a[241] & b[374])^(a[240] & b[375])^(a[239] & b[376])^(a[238] & b[377])^(a[237] & b[378])^(a[236] & b[379])^(a[235] & b[380])^(a[234] & b[381])^(a[233] & b[382])^(a[232] & b[383])^(a[231] & b[384])^(a[230] & b[385])^(a[229] & b[386])^(a[228] & b[387])^(a[227] & b[388])^(a[226] & b[389])^(a[225] & b[390])^(a[224] & b[391])^(a[223] & b[392])^(a[222] & b[393])^(a[221] & b[394])^(a[220] & b[395])^(a[219] & b[396])^(a[218] & b[397])^(a[217] & b[398])^(a[216] & b[399])^(a[215] & b[400])^(a[214] & b[401])^(a[213] & b[402])^(a[212] & b[403])^(a[211] & b[404])^(a[210] & b[405])^(a[209] & b[406])^(a[208] & b[407])^(a[207] & b[408]);
assign y[616] = (a[408] & b[208])^(a[407] & b[209])^(a[406] & b[210])^(a[405] & b[211])^(a[404] & b[212])^(a[403] & b[213])^(a[402] & b[214])^(a[401] & b[215])^(a[400] & b[216])^(a[399] & b[217])^(a[398] & b[218])^(a[397] & b[219])^(a[396] & b[220])^(a[395] & b[221])^(a[394] & b[222])^(a[393] & b[223])^(a[392] & b[224])^(a[391] & b[225])^(a[390] & b[226])^(a[389] & b[227])^(a[388] & b[228])^(a[387] & b[229])^(a[386] & b[230])^(a[385] & b[231])^(a[384] & b[232])^(a[383] & b[233])^(a[382] & b[234])^(a[381] & b[235])^(a[380] & b[236])^(a[379] & b[237])^(a[378] & b[238])^(a[377] & b[239])^(a[376] & b[240])^(a[375] & b[241])^(a[374] & b[242])^(a[373] & b[243])^(a[372] & b[244])^(a[371] & b[245])^(a[370] & b[246])^(a[369] & b[247])^(a[368] & b[248])^(a[367] & b[249])^(a[366] & b[250])^(a[365] & b[251])^(a[364] & b[252])^(a[363] & b[253])^(a[362] & b[254])^(a[361] & b[255])^(a[360] & b[256])^(a[359] & b[257])^(a[358] & b[258])^(a[357] & b[259])^(a[356] & b[260])^(a[355] & b[261])^(a[354] & b[262])^(a[353] & b[263])^(a[352] & b[264])^(a[351] & b[265])^(a[350] & b[266])^(a[349] & b[267])^(a[348] & b[268])^(a[347] & b[269])^(a[346] & b[270])^(a[345] & b[271])^(a[344] & b[272])^(a[343] & b[273])^(a[342] & b[274])^(a[341] & b[275])^(a[340] & b[276])^(a[339] & b[277])^(a[338] & b[278])^(a[337] & b[279])^(a[336] & b[280])^(a[335] & b[281])^(a[334] & b[282])^(a[333] & b[283])^(a[332] & b[284])^(a[331] & b[285])^(a[330] & b[286])^(a[329] & b[287])^(a[328] & b[288])^(a[327] & b[289])^(a[326] & b[290])^(a[325] & b[291])^(a[324] & b[292])^(a[323] & b[293])^(a[322] & b[294])^(a[321] & b[295])^(a[320] & b[296])^(a[319] & b[297])^(a[318] & b[298])^(a[317] & b[299])^(a[316] & b[300])^(a[315] & b[301])^(a[314] & b[302])^(a[313] & b[303])^(a[312] & b[304])^(a[311] & b[305])^(a[310] & b[306])^(a[309] & b[307])^(a[308] & b[308])^(a[307] & b[309])^(a[306] & b[310])^(a[305] & b[311])^(a[304] & b[312])^(a[303] & b[313])^(a[302] & b[314])^(a[301] & b[315])^(a[300] & b[316])^(a[299] & b[317])^(a[298] & b[318])^(a[297] & b[319])^(a[296] & b[320])^(a[295] & b[321])^(a[294] & b[322])^(a[293] & b[323])^(a[292] & b[324])^(a[291] & b[325])^(a[290] & b[326])^(a[289] & b[327])^(a[288] & b[328])^(a[287] & b[329])^(a[286] & b[330])^(a[285] & b[331])^(a[284] & b[332])^(a[283] & b[333])^(a[282] & b[334])^(a[281] & b[335])^(a[280] & b[336])^(a[279] & b[337])^(a[278] & b[338])^(a[277] & b[339])^(a[276] & b[340])^(a[275] & b[341])^(a[274] & b[342])^(a[273] & b[343])^(a[272] & b[344])^(a[271] & b[345])^(a[270] & b[346])^(a[269] & b[347])^(a[268] & b[348])^(a[267] & b[349])^(a[266] & b[350])^(a[265] & b[351])^(a[264] & b[352])^(a[263] & b[353])^(a[262] & b[354])^(a[261] & b[355])^(a[260] & b[356])^(a[259] & b[357])^(a[258] & b[358])^(a[257] & b[359])^(a[256] & b[360])^(a[255] & b[361])^(a[254] & b[362])^(a[253] & b[363])^(a[252] & b[364])^(a[251] & b[365])^(a[250] & b[366])^(a[249] & b[367])^(a[248] & b[368])^(a[247] & b[369])^(a[246] & b[370])^(a[245] & b[371])^(a[244] & b[372])^(a[243] & b[373])^(a[242] & b[374])^(a[241] & b[375])^(a[240] & b[376])^(a[239] & b[377])^(a[238] & b[378])^(a[237] & b[379])^(a[236] & b[380])^(a[235] & b[381])^(a[234] & b[382])^(a[233] & b[383])^(a[232] & b[384])^(a[231] & b[385])^(a[230] & b[386])^(a[229] & b[387])^(a[228] & b[388])^(a[227] & b[389])^(a[226] & b[390])^(a[225] & b[391])^(a[224] & b[392])^(a[223] & b[393])^(a[222] & b[394])^(a[221] & b[395])^(a[220] & b[396])^(a[219] & b[397])^(a[218] & b[398])^(a[217] & b[399])^(a[216] & b[400])^(a[215] & b[401])^(a[214] & b[402])^(a[213] & b[403])^(a[212] & b[404])^(a[211] & b[405])^(a[210] & b[406])^(a[209] & b[407])^(a[208] & b[408]);
assign y[617] = (a[408] & b[209])^(a[407] & b[210])^(a[406] & b[211])^(a[405] & b[212])^(a[404] & b[213])^(a[403] & b[214])^(a[402] & b[215])^(a[401] & b[216])^(a[400] & b[217])^(a[399] & b[218])^(a[398] & b[219])^(a[397] & b[220])^(a[396] & b[221])^(a[395] & b[222])^(a[394] & b[223])^(a[393] & b[224])^(a[392] & b[225])^(a[391] & b[226])^(a[390] & b[227])^(a[389] & b[228])^(a[388] & b[229])^(a[387] & b[230])^(a[386] & b[231])^(a[385] & b[232])^(a[384] & b[233])^(a[383] & b[234])^(a[382] & b[235])^(a[381] & b[236])^(a[380] & b[237])^(a[379] & b[238])^(a[378] & b[239])^(a[377] & b[240])^(a[376] & b[241])^(a[375] & b[242])^(a[374] & b[243])^(a[373] & b[244])^(a[372] & b[245])^(a[371] & b[246])^(a[370] & b[247])^(a[369] & b[248])^(a[368] & b[249])^(a[367] & b[250])^(a[366] & b[251])^(a[365] & b[252])^(a[364] & b[253])^(a[363] & b[254])^(a[362] & b[255])^(a[361] & b[256])^(a[360] & b[257])^(a[359] & b[258])^(a[358] & b[259])^(a[357] & b[260])^(a[356] & b[261])^(a[355] & b[262])^(a[354] & b[263])^(a[353] & b[264])^(a[352] & b[265])^(a[351] & b[266])^(a[350] & b[267])^(a[349] & b[268])^(a[348] & b[269])^(a[347] & b[270])^(a[346] & b[271])^(a[345] & b[272])^(a[344] & b[273])^(a[343] & b[274])^(a[342] & b[275])^(a[341] & b[276])^(a[340] & b[277])^(a[339] & b[278])^(a[338] & b[279])^(a[337] & b[280])^(a[336] & b[281])^(a[335] & b[282])^(a[334] & b[283])^(a[333] & b[284])^(a[332] & b[285])^(a[331] & b[286])^(a[330] & b[287])^(a[329] & b[288])^(a[328] & b[289])^(a[327] & b[290])^(a[326] & b[291])^(a[325] & b[292])^(a[324] & b[293])^(a[323] & b[294])^(a[322] & b[295])^(a[321] & b[296])^(a[320] & b[297])^(a[319] & b[298])^(a[318] & b[299])^(a[317] & b[300])^(a[316] & b[301])^(a[315] & b[302])^(a[314] & b[303])^(a[313] & b[304])^(a[312] & b[305])^(a[311] & b[306])^(a[310] & b[307])^(a[309] & b[308])^(a[308] & b[309])^(a[307] & b[310])^(a[306] & b[311])^(a[305] & b[312])^(a[304] & b[313])^(a[303] & b[314])^(a[302] & b[315])^(a[301] & b[316])^(a[300] & b[317])^(a[299] & b[318])^(a[298] & b[319])^(a[297] & b[320])^(a[296] & b[321])^(a[295] & b[322])^(a[294] & b[323])^(a[293] & b[324])^(a[292] & b[325])^(a[291] & b[326])^(a[290] & b[327])^(a[289] & b[328])^(a[288] & b[329])^(a[287] & b[330])^(a[286] & b[331])^(a[285] & b[332])^(a[284] & b[333])^(a[283] & b[334])^(a[282] & b[335])^(a[281] & b[336])^(a[280] & b[337])^(a[279] & b[338])^(a[278] & b[339])^(a[277] & b[340])^(a[276] & b[341])^(a[275] & b[342])^(a[274] & b[343])^(a[273] & b[344])^(a[272] & b[345])^(a[271] & b[346])^(a[270] & b[347])^(a[269] & b[348])^(a[268] & b[349])^(a[267] & b[350])^(a[266] & b[351])^(a[265] & b[352])^(a[264] & b[353])^(a[263] & b[354])^(a[262] & b[355])^(a[261] & b[356])^(a[260] & b[357])^(a[259] & b[358])^(a[258] & b[359])^(a[257] & b[360])^(a[256] & b[361])^(a[255] & b[362])^(a[254] & b[363])^(a[253] & b[364])^(a[252] & b[365])^(a[251] & b[366])^(a[250] & b[367])^(a[249] & b[368])^(a[248] & b[369])^(a[247] & b[370])^(a[246] & b[371])^(a[245] & b[372])^(a[244] & b[373])^(a[243] & b[374])^(a[242] & b[375])^(a[241] & b[376])^(a[240] & b[377])^(a[239] & b[378])^(a[238] & b[379])^(a[237] & b[380])^(a[236] & b[381])^(a[235] & b[382])^(a[234] & b[383])^(a[233] & b[384])^(a[232] & b[385])^(a[231] & b[386])^(a[230] & b[387])^(a[229] & b[388])^(a[228] & b[389])^(a[227] & b[390])^(a[226] & b[391])^(a[225] & b[392])^(a[224] & b[393])^(a[223] & b[394])^(a[222] & b[395])^(a[221] & b[396])^(a[220] & b[397])^(a[219] & b[398])^(a[218] & b[399])^(a[217] & b[400])^(a[216] & b[401])^(a[215] & b[402])^(a[214] & b[403])^(a[213] & b[404])^(a[212] & b[405])^(a[211] & b[406])^(a[210] & b[407])^(a[209] & b[408]);
assign y[618] = (a[408] & b[210])^(a[407] & b[211])^(a[406] & b[212])^(a[405] & b[213])^(a[404] & b[214])^(a[403] & b[215])^(a[402] & b[216])^(a[401] & b[217])^(a[400] & b[218])^(a[399] & b[219])^(a[398] & b[220])^(a[397] & b[221])^(a[396] & b[222])^(a[395] & b[223])^(a[394] & b[224])^(a[393] & b[225])^(a[392] & b[226])^(a[391] & b[227])^(a[390] & b[228])^(a[389] & b[229])^(a[388] & b[230])^(a[387] & b[231])^(a[386] & b[232])^(a[385] & b[233])^(a[384] & b[234])^(a[383] & b[235])^(a[382] & b[236])^(a[381] & b[237])^(a[380] & b[238])^(a[379] & b[239])^(a[378] & b[240])^(a[377] & b[241])^(a[376] & b[242])^(a[375] & b[243])^(a[374] & b[244])^(a[373] & b[245])^(a[372] & b[246])^(a[371] & b[247])^(a[370] & b[248])^(a[369] & b[249])^(a[368] & b[250])^(a[367] & b[251])^(a[366] & b[252])^(a[365] & b[253])^(a[364] & b[254])^(a[363] & b[255])^(a[362] & b[256])^(a[361] & b[257])^(a[360] & b[258])^(a[359] & b[259])^(a[358] & b[260])^(a[357] & b[261])^(a[356] & b[262])^(a[355] & b[263])^(a[354] & b[264])^(a[353] & b[265])^(a[352] & b[266])^(a[351] & b[267])^(a[350] & b[268])^(a[349] & b[269])^(a[348] & b[270])^(a[347] & b[271])^(a[346] & b[272])^(a[345] & b[273])^(a[344] & b[274])^(a[343] & b[275])^(a[342] & b[276])^(a[341] & b[277])^(a[340] & b[278])^(a[339] & b[279])^(a[338] & b[280])^(a[337] & b[281])^(a[336] & b[282])^(a[335] & b[283])^(a[334] & b[284])^(a[333] & b[285])^(a[332] & b[286])^(a[331] & b[287])^(a[330] & b[288])^(a[329] & b[289])^(a[328] & b[290])^(a[327] & b[291])^(a[326] & b[292])^(a[325] & b[293])^(a[324] & b[294])^(a[323] & b[295])^(a[322] & b[296])^(a[321] & b[297])^(a[320] & b[298])^(a[319] & b[299])^(a[318] & b[300])^(a[317] & b[301])^(a[316] & b[302])^(a[315] & b[303])^(a[314] & b[304])^(a[313] & b[305])^(a[312] & b[306])^(a[311] & b[307])^(a[310] & b[308])^(a[309] & b[309])^(a[308] & b[310])^(a[307] & b[311])^(a[306] & b[312])^(a[305] & b[313])^(a[304] & b[314])^(a[303] & b[315])^(a[302] & b[316])^(a[301] & b[317])^(a[300] & b[318])^(a[299] & b[319])^(a[298] & b[320])^(a[297] & b[321])^(a[296] & b[322])^(a[295] & b[323])^(a[294] & b[324])^(a[293] & b[325])^(a[292] & b[326])^(a[291] & b[327])^(a[290] & b[328])^(a[289] & b[329])^(a[288] & b[330])^(a[287] & b[331])^(a[286] & b[332])^(a[285] & b[333])^(a[284] & b[334])^(a[283] & b[335])^(a[282] & b[336])^(a[281] & b[337])^(a[280] & b[338])^(a[279] & b[339])^(a[278] & b[340])^(a[277] & b[341])^(a[276] & b[342])^(a[275] & b[343])^(a[274] & b[344])^(a[273] & b[345])^(a[272] & b[346])^(a[271] & b[347])^(a[270] & b[348])^(a[269] & b[349])^(a[268] & b[350])^(a[267] & b[351])^(a[266] & b[352])^(a[265] & b[353])^(a[264] & b[354])^(a[263] & b[355])^(a[262] & b[356])^(a[261] & b[357])^(a[260] & b[358])^(a[259] & b[359])^(a[258] & b[360])^(a[257] & b[361])^(a[256] & b[362])^(a[255] & b[363])^(a[254] & b[364])^(a[253] & b[365])^(a[252] & b[366])^(a[251] & b[367])^(a[250] & b[368])^(a[249] & b[369])^(a[248] & b[370])^(a[247] & b[371])^(a[246] & b[372])^(a[245] & b[373])^(a[244] & b[374])^(a[243] & b[375])^(a[242] & b[376])^(a[241] & b[377])^(a[240] & b[378])^(a[239] & b[379])^(a[238] & b[380])^(a[237] & b[381])^(a[236] & b[382])^(a[235] & b[383])^(a[234] & b[384])^(a[233] & b[385])^(a[232] & b[386])^(a[231] & b[387])^(a[230] & b[388])^(a[229] & b[389])^(a[228] & b[390])^(a[227] & b[391])^(a[226] & b[392])^(a[225] & b[393])^(a[224] & b[394])^(a[223] & b[395])^(a[222] & b[396])^(a[221] & b[397])^(a[220] & b[398])^(a[219] & b[399])^(a[218] & b[400])^(a[217] & b[401])^(a[216] & b[402])^(a[215] & b[403])^(a[214] & b[404])^(a[213] & b[405])^(a[212] & b[406])^(a[211] & b[407])^(a[210] & b[408]);
assign y[619] = (a[408] & b[211])^(a[407] & b[212])^(a[406] & b[213])^(a[405] & b[214])^(a[404] & b[215])^(a[403] & b[216])^(a[402] & b[217])^(a[401] & b[218])^(a[400] & b[219])^(a[399] & b[220])^(a[398] & b[221])^(a[397] & b[222])^(a[396] & b[223])^(a[395] & b[224])^(a[394] & b[225])^(a[393] & b[226])^(a[392] & b[227])^(a[391] & b[228])^(a[390] & b[229])^(a[389] & b[230])^(a[388] & b[231])^(a[387] & b[232])^(a[386] & b[233])^(a[385] & b[234])^(a[384] & b[235])^(a[383] & b[236])^(a[382] & b[237])^(a[381] & b[238])^(a[380] & b[239])^(a[379] & b[240])^(a[378] & b[241])^(a[377] & b[242])^(a[376] & b[243])^(a[375] & b[244])^(a[374] & b[245])^(a[373] & b[246])^(a[372] & b[247])^(a[371] & b[248])^(a[370] & b[249])^(a[369] & b[250])^(a[368] & b[251])^(a[367] & b[252])^(a[366] & b[253])^(a[365] & b[254])^(a[364] & b[255])^(a[363] & b[256])^(a[362] & b[257])^(a[361] & b[258])^(a[360] & b[259])^(a[359] & b[260])^(a[358] & b[261])^(a[357] & b[262])^(a[356] & b[263])^(a[355] & b[264])^(a[354] & b[265])^(a[353] & b[266])^(a[352] & b[267])^(a[351] & b[268])^(a[350] & b[269])^(a[349] & b[270])^(a[348] & b[271])^(a[347] & b[272])^(a[346] & b[273])^(a[345] & b[274])^(a[344] & b[275])^(a[343] & b[276])^(a[342] & b[277])^(a[341] & b[278])^(a[340] & b[279])^(a[339] & b[280])^(a[338] & b[281])^(a[337] & b[282])^(a[336] & b[283])^(a[335] & b[284])^(a[334] & b[285])^(a[333] & b[286])^(a[332] & b[287])^(a[331] & b[288])^(a[330] & b[289])^(a[329] & b[290])^(a[328] & b[291])^(a[327] & b[292])^(a[326] & b[293])^(a[325] & b[294])^(a[324] & b[295])^(a[323] & b[296])^(a[322] & b[297])^(a[321] & b[298])^(a[320] & b[299])^(a[319] & b[300])^(a[318] & b[301])^(a[317] & b[302])^(a[316] & b[303])^(a[315] & b[304])^(a[314] & b[305])^(a[313] & b[306])^(a[312] & b[307])^(a[311] & b[308])^(a[310] & b[309])^(a[309] & b[310])^(a[308] & b[311])^(a[307] & b[312])^(a[306] & b[313])^(a[305] & b[314])^(a[304] & b[315])^(a[303] & b[316])^(a[302] & b[317])^(a[301] & b[318])^(a[300] & b[319])^(a[299] & b[320])^(a[298] & b[321])^(a[297] & b[322])^(a[296] & b[323])^(a[295] & b[324])^(a[294] & b[325])^(a[293] & b[326])^(a[292] & b[327])^(a[291] & b[328])^(a[290] & b[329])^(a[289] & b[330])^(a[288] & b[331])^(a[287] & b[332])^(a[286] & b[333])^(a[285] & b[334])^(a[284] & b[335])^(a[283] & b[336])^(a[282] & b[337])^(a[281] & b[338])^(a[280] & b[339])^(a[279] & b[340])^(a[278] & b[341])^(a[277] & b[342])^(a[276] & b[343])^(a[275] & b[344])^(a[274] & b[345])^(a[273] & b[346])^(a[272] & b[347])^(a[271] & b[348])^(a[270] & b[349])^(a[269] & b[350])^(a[268] & b[351])^(a[267] & b[352])^(a[266] & b[353])^(a[265] & b[354])^(a[264] & b[355])^(a[263] & b[356])^(a[262] & b[357])^(a[261] & b[358])^(a[260] & b[359])^(a[259] & b[360])^(a[258] & b[361])^(a[257] & b[362])^(a[256] & b[363])^(a[255] & b[364])^(a[254] & b[365])^(a[253] & b[366])^(a[252] & b[367])^(a[251] & b[368])^(a[250] & b[369])^(a[249] & b[370])^(a[248] & b[371])^(a[247] & b[372])^(a[246] & b[373])^(a[245] & b[374])^(a[244] & b[375])^(a[243] & b[376])^(a[242] & b[377])^(a[241] & b[378])^(a[240] & b[379])^(a[239] & b[380])^(a[238] & b[381])^(a[237] & b[382])^(a[236] & b[383])^(a[235] & b[384])^(a[234] & b[385])^(a[233] & b[386])^(a[232] & b[387])^(a[231] & b[388])^(a[230] & b[389])^(a[229] & b[390])^(a[228] & b[391])^(a[227] & b[392])^(a[226] & b[393])^(a[225] & b[394])^(a[224] & b[395])^(a[223] & b[396])^(a[222] & b[397])^(a[221] & b[398])^(a[220] & b[399])^(a[219] & b[400])^(a[218] & b[401])^(a[217] & b[402])^(a[216] & b[403])^(a[215] & b[404])^(a[214] & b[405])^(a[213] & b[406])^(a[212] & b[407])^(a[211] & b[408]);
assign y[620] = (a[408] & b[212])^(a[407] & b[213])^(a[406] & b[214])^(a[405] & b[215])^(a[404] & b[216])^(a[403] & b[217])^(a[402] & b[218])^(a[401] & b[219])^(a[400] & b[220])^(a[399] & b[221])^(a[398] & b[222])^(a[397] & b[223])^(a[396] & b[224])^(a[395] & b[225])^(a[394] & b[226])^(a[393] & b[227])^(a[392] & b[228])^(a[391] & b[229])^(a[390] & b[230])^(a[389] & b[231])^(a[388] & b[232])^(a[387] & b[233])^(a[386] & b[234])^(a[385] & b[235])^(a[384] & b[236])^(a[383] & b[237])^(a[382] & b[238])^(a[381] & b[239])^(a[380] & b[240])^(a[379] & b[241])^(a[378] & b[242])^(a[377] & b[243])^(a[376] & b[244])^(a[375] & b[245])^(a[374] & b[246])^(a[373] & b[247])^(a[372] & b[248])^(a[371] & b[249])^(a[370] & b[250])^(a[369] & b[251])^(a[368] & b[252])^(a[367] & b[253])^(a[366] & b[254])^(a[365] & b[255])^(a[364] & b[256])^(a[363] & b[257])^(a[362] & b[258])^(a[361] & b[259])^(a[360] & b[260])^(a[359] & b[261])^(a[358] & b[262])^(a[357] & b[263])^(a[356] & b[264])^(a[355] & b[265])^(a[354] & b[266])^(a[353] & b[267])^(a[352] & b[268])^(a[351] & b[269])^(a[350] & b[270])^(a[349] & b[271])^(a[348] & b[272])^(a[347] & b[273])^(a[346] & b[274])^(a[345] & b[275])^(a[344] & b[276])^(a[343] & b[277])^(a[342] & b[278])^(a[341] & b[279])^(a[340] & b[280])^(a[339] & b[281])^(a[338] & b[282])^(a[337] & b[283])^(a[336] & b[284])^(a[335] & b[285])^(a[334] & b[286])^(a[333] & b[287])^(a[332] & b[288])^(a[331] & b[289])^(a[330] & b[290])^(a[329] & b[291])^(a[328] & b[292])^(a[327] & b[293])^(a[326] & b[294])^(a[325] & b[295])^(a[324] & b[296])^(a[323] & b[297])^(a[322] & b[298])^(a[321] & b[299])^(a[320] & b[300])^(a[319] & b[301])^(a[318] & b[302])^(a[317] & b[303])^(a[316] & b[304])^(a[315] & b[305])^(a[314] & b[306])^(a[313] & b[307])^(a[312] & b[308])^(a[311] & b[309])^(a[310] & b[310])^(a[309] & b[311])^(a[308] & b[312])^(a[307] & b[313])^(a[306] & b[314])^(a[305] & b[315])^(a[304] & b[316])^(a[303] & b[317])^(a[302] & b[318])^(a[301] & b[319])^(a[300] & b[320])^(a[299] & b[321])^(a[298] & b[322])^(a[297] & b[323])^(a[296] & b[324])^(a[295] & b[325])^(a[294] & b[326])^(a[293] & b[327])^(a[292] & b[328])^(a[291] & b[329])^(a[290] & b[330])^(a[289] & b[331])^(a[288] & b[332])^(a[287] & b[333])^(a[286] & b[334])^(a[285] & b[335])^(a[284] & b[336])^(a[283] & b[337])^(a[282] & b[338])^(a[281] & b[339])^(a[280] & b[340])^(a[279] & b[341])^(a[278] & b[342])^(a[277] & b[343])^(a[276] & b[344])^(a[275] & b[345])^(a[274] & b[346])^(a[273] & b[347])^(a[272] & b[348])^(a[271] & b[349])^(a[270] & b[350])^(a[269] & b[351])^(a[268] & b[352])^(a[267] & b[353])^(a[266] & b[354])^(a[265] & b[355])^(a[264] & b[356])^(a[263] & b[357])^(a[262] & b[358])^(a[261] & b[359])^(a[260] & b[360])^(a[259] & b[361])^(a[258] & b[362])^(a[257] & b[363])^(a[256] & b[364])^(a[255] & b[365])^(a[254] & b[366])^(a[253] & b[367])^(a[252] & b[368])^(a[251] & b[369])^(a[250] & b[370])^(a[249] & b[371])^(a[248] & b[372])^(a[247] & b[373])^(a[246] & b[374])^(a[245] & b[375])^(a[244] & b[376])^(a[243] & b[377])^(a[242] & b[378])^(a[241] & b[379])^(a[240] & b[380])^(a[239] & b[381])^(a[238] & b[382])^(a[237] & b[383])^(a[236] & b[384])^(a[235] & b[385])^(a[234] & b[386])^(a[233] & b[387])^(a[232] & b[388])^(a[231] & b[389])^(a[230] & b[390])^(a[229] & b[391])^(a[228] & b[392])^(a[227] & b[393])^(a[226] & b[394])^(a[225] & b[395])^(a[224] & b[396])^(a[223] & b[397])^(a[222] & b[398])^(a[221] & b[399])^(a[220] & b[400])^(a[219] & b[401])^(a[218] & b[402])^(a[217] & b[403])^(a[216] & b[404])^(a[215] & b[405])^(a[214] & b[406])^(a[213] & b[407])^(a[212] & b[408]);
assign y[621] = (a[408] & b[213])^(a[407] & b[214])^(a[406] & b[215])^(a[405] & b[216])^(a[404] & b[217])^(a[403] & b[218])^(a[402] & b[219])^(a[401] & b[220])^(a[400] & b[221])^(a[399] & b[222])^(a[398] & b[223])^(a[397] & b[224])^(a[396] & b[225])^(a[395] & b[226])^(a[394] & b[227])^(a[393] & b[228])^(a[392] & b[229])^(a[391] & b[230])^(a[390] & b[231])^(a[389] & b[232])^(a[388] & b[233])^(a[387] & b[234])^(a[386] & b[235])^(a[385] & b[236])^(a[384] & b[237])^(a[383] & b[238])^(a[382] & b[239])^(a[381] & b[240])^(a[380] & b[241])^(a[379] & b[242])^(a[378] & b[243])^(a[377] & b[244])^(a[376] & b[245])^(a[375] & b[246])^(a[374] & b[247])^(a[373] & b[248])^(a[372] & b[249])^(a[371] & b[250])^(a[370] & b[251])^(a[369] & b[252])^(a[368] & b[253])^(a[367] & b[254])^(a[366] & b[255])^(a[365] & b[256])^(a[364] & b[257])^(a[363] & b[258])^(a[362] & b[259])^(a[361] & b[260])^(a[360] & b[261])^(a[359] & b[262])^(a[358] & b[263])^(a[357] & b[264])^(a[356] & b[265])^(a[355] & b[266])^(a[354] & b[267])^(a[353] & b[268])^(a[352] & b[269])^(a[351] & b[270])^(a[350] & b[271])^(a[349] & b[272])^(a[348] & b[273])^(a[347] & b[274])^(a[346] & b[275])^(a[345] & b[276])^(a[344] & b[277])^(a[343] & b[278])^(a[342] & b[279])^(a[341] & b[280])^(a[340] & b[281])^(a[339] & b[282])^(a[338] & b[283])^(a[337] & b[284])^(a[336] & b[285])^(a[335] & b[286])^(a[334] & b[287])^(a[333] & b[288])^(a[332] & b[289])^(a[331] & b[290])^(a[330] & b[291])^(a[329] & b[292])^(a[328] & b[293])^(a[327] & b[294])^(a[326] & b[295])^(a[325] & b[296])^(a[324] & b[297])^(a[323] & b[298])^(a[322] & b[299])^(a[321] & b[300])^(a[320] & b[301])^(a[319] & b[302])^(a[318] & b[303])^(a[317] & b[304])^(a[316] & b[305])^(a[315] & b[306])^(a[314] & b[307])^(a[313] & b[308])^(a[312] & b[309])^(a[311] & b[310])^(a[310] & b[311])^(a[309] & b[312])^(a[308] & b[313])^(a[307] & b[314])^(a[306] & b[315])^(a[305] & b[316])^(a[304] & b[317])^(a[303] & b[318])^(a[302] & b[319])^(a[301] & b[320])^(a[300] & b[321])^(a[299] & b[322])^(a[298] & b[323])^(a[297] & b[324])^(a[296] & b[325])^(a[295] & b[326])^(a[294] & b[327])^(a[293] & b[328])^(a[292] & b[329])^(a[291] & b[330])^(a[290] & b[331])^(a[289] & b[332])^(a[288] & b[333])^(a[287] & b[334])^(a[286] & b[335])^(a[285] & b[336])^(a[284] & b[337])^(a[283] & b[338])^(a[282] & b[339])^(a[281] & b[340])^(a[280] & b[341])^(a[279] & b[342])^(a[278] & b[343])^(a[277] & b[344])^(a[276] & b[345])^(a[275] & b[346])^(a[274] & b[347])^(a[273] & b[348])^(a[272] & b[349])^(a[271] & b[350])^(a[270] & b[351])^(a[269] & b[352])^(a[268] & b[353])^(a[267] & b[354])^(a[266] & b[355])^(a[265] & b[356])^(a[264] & b[357])^(a[263] & b[358])^(a[262] & b[359])^(a[261] & b[360])^(a[260] & b[361])^(a[259] & b[362])^(a[258] & b[363])^(a[257] & b[364])^(a[256] & b[365])^(a[255] & b[366])^(a[254] & b[367])^(a[253] & b[368])^(a[252] & b[369])^(a[251] & b[370])^(a[250] & b[371])^(a[249] & b[372])^(a[248] & b[373])^(a[247] & b[374])^(a[246] & b[375])^(a[245] & b[376])^(a[244] & b[377])^(a[243] & b[378])^(a[242] & b[379])^(a[241] & b[380])^(a[240] & b[381])^(a[239] & b[382])^(a[238] & b[383])^(a[237] & b[384])^(a[236] & b[385])^(a[235] & b[386])^(a[234] & b[387])^(a[233] & b[388])^(a[232] & b[389])^(a[231] & b[390])^(a[230] & b[391])^(a[229] & b[392])^(a[228] & b[393])^(a[227] & b[394])^(a[226] & b[395])^(a[225] & b[396])^(a[224] & b[397])^(a[223] & b[398])^(a[222] & b[399])^(a[221] & b[400])^(a[220] & b[401])^(a[219] & b[402])^(a[218] & b[403])^(a[217] & b[404])^(a[216] & b[405])^(a[215] & b[406])^(a[214] & b[407])^(a[213] & b[408]);
assign y[622] = (a[408] & b[214])^(a[407] & b[215])^(a[406] & b[216])^(a[405] & b[217])^(a[404] & b[218])^(a[403] & b[219])^(a[402] & b[220])^(a[401] & b[221])^(a[400] & b[222])^(a[399] & b[223])^(a[398] & b[224])^(a[397] & b[225])^(a[396] & b[226])^(a[395] & b[227])^(a[394] & b[228])^(a[393] & b[229])^(a[392] & b[230])^(a[391] & b[231])^(a[390] & b[232])^(a[389] & b[233])^(a[388] & b[234])^(a[387] & b[235])^(a[386] & b[236])^(a[385] & b[237])^(a[384] & b[238])^(a[383] & b[239])^(a[382] & b[240])^(a[381] & b[241])^(a[380] & b[242])^(a[379] & b[243])^(a[378] & b[244])^(a[377] & b[245])^(a[376] & b[246])^(a[375] & b[247])^(a[374] & b[248])^(a[373] & b[249])^(a[372] & b[250])^(a[371] & b[251])^(a[370] & b[252])^(a[369] & b[253])^(a[368] & b[254])^(a[367] & b[255])^(a[366] & b[256])^(a[365] & b[257])^(a[364] & b[258])^(a[363] & b[259])^(a[362] & b[260])^(a[361] & b[261])^(a[360] & b[262])^(a[359] & b[263])^(a[358] & b[264])^(a[357] & b[265])^(a[356] & b[266])^(a[355] & b[267])^(a[354] & b[268])^(a[353] & b[269])^(a[352] & b[270])^(a[351] & b[271])^(a[350] & b[272])^(a[349] & b[273])^(a[348] & b[274])^(a[347] & b[275])^(a[346] & b[276])^(a[345] & b[277])^(a[344] & b[278])^(a[343] & b[279])^(a[342] & b[280])^(a[341] & b[281])^(a[340] & b[282])^(a[339] & b[283])^(a[338] & b[284])^(a[337] & b[285])^(a[336] & b[286])^(a[335] & b[287])^(a[334] & b[288])^(a[333] & b[289])^(a[332] & b[290])^(a[331] & b[291])^(a[330] & b[292])^(a[329] & b[293])^(a[328] & b[294])^(a[327] & b[295])^(a[326] & b[296])^(a[325] & b[297])^(a[324] & b[298])^(a[323] & b[299])^(a[322] & b[300])^(a[321] & b[301])^(a[320] & b[302])^(a[319] & b[303])^(a[318] & b[304])^(a[317] & b[305])^(a[316] & b[306])^(a[315] & b[307])^(a[314] & b[308])^(a[313] & b[309])^(a[312] & b[310])^(a[311] & b[311])^(a[310] & b[312])^(a[309] & b[313])^(a[308] & b[314])^(a[307] & b[315])^(a[306] & b[316])^(a[305] & b[317])^(a[304] & b[318])^(a[303] & b[319])^(a[302] & b[320])^(a[301] & b[321])^(a[300] & b[322])^(a[299] & b[323])^(a[298] & b[324])^(a[297] & b[325])^(a[296] & b[326])^(a[295] & b[327])^(a[294] & b[328])^(a[293] & b[329])^(a[292] & b[330])^(a[291] & b[331])^(a[290] & b[332])^(a[289] & b[333])^(a[288] & b[334])^(a[287] & b[335])^(a[286] & b[336])^(a[285] & b[337])^(a[284] & b[338])^(a[283] & b[339])^(a[282] & b[340])^(a[281] & b[341])^(a[280] & b[342])^(a[279] & b[343])^(a[278] & b[344])^(a[277] & b[345])^(a[276] & b[346])^(a[275] & b[347])^(a[274] & b[348])^(a[273] & b[349])^(a[272] & b[350])^(a[271] & b[351])^(a[270] & b[352])^(a[269] & b[353])^(a[268] & b[354])^(a[267] & b[355])^(a[266] & b[356])^(a[265] & b[357])^(a[264] & b[358])^(a[263] & b[359])^(a[262] & b[360])^(a[261] & b[361])^(a[260] & b[362])^(a[259] & b[363])^(a[258] & b[364])^(a[257] & b[365])^(a[256] & b[366])^(a[255] & b[367])^(a[254] & b[368])^(a[253] & b[369])^(a[252] & b[370])^(a[251] & b[371])^(a[250] & b[372])^(a[249] & b[373])^(a[248] & b[374])^(a[247] & b[375])^(a[246] & b[376])^(a[245] & b[377])^(a[244] & b[378])^(a[243] & b[379])^(a[242] & b[380])^(a[241] & b[381])^(a[240] & b[382])^(a[239] & b[383])^(a[238] & b[384])^(a[237] & b[385])^(a[236] & b[386])^(a[235] & b[387])^(a[234] & b[388])^(a[233] & b[389])^(a[232] & b[390])^(a[231] & b[391])^(a[230] & b[392])^(a[229] & b[393])^(a[228] & b[394])^(a[227] & b[395])^(a[226] & b[396])^(a[225] & b[397])^(a[224] & b[398])^(a[223] & b[399])^(a[222] & b[400])^(a[221] & b[401])^(a[220] & b[402])^(a[219] & b[403])^(a[218] & b[404])^(a[217] & b[405])^(a[216] & b[406])^(a[215] & b[407])^(a[214] & b[408]);
assign y[623] = (a[408] & b[215])^(a[407] & b[216])^(a[406] & b[217])^(a[405] & b[218])^(a[404] & b[219])^(a[403] & b[220])^(a[402] & b[221])^(a[401] & b[222])^(a[400] & b[223])^(a[399] & b[224])^(a[398] & b[225])^(a[397] & b[226])^(a[396] & b[227])^(a[395] & b[228])^(a[394] & b[229])^(a[393] & b[230])^(a[392] & b[231])^(a[391] & b[232])^(a[390] & b[233])^(a[389] & b[234])^(a[388] & b[235])^(a[387] & b[236])^(a[386] & b[237])^(a[385] & b[238])^(a[384] & b[239])^(a[383] & b[240])^(a[382] & b[241])^(a[381] & b[242])^(a[380] & b[243])^(a[379] & b[244])^(a[378] & b[245])^(a[377] & b[246])^(a[376] & b[247])^(a[375] & b[248])^(a[374] & b[249])^(a[373] & b[250])^(a[372] & b[251])^(a[371] & b[252])^(a[370] & b[253])^(a[369] & b[254])^(a[368] & b[255])^(a[367] & b[256])^(a[366] & b[257])^(a[365] & b[258])^(a[364] & b[259])^(a[363] & b[260])^(a[362] & b[261])^(a[361] & b[262])^(a[360] & b[263])^(a[359] & b[264])^(a[358] & b[265])^(a[357] & b[266])^(a[356] & b[267])^(a[355] & b[268])^(a[354] & b[269])^(a[353] & b[270])^(a[352] & b[271])^(a[351] & b[272])^(a[350] & b[273])^(a[349] & b[274])^(a[348] & b[275])^(a[347] & b[276])^(a[346] & b[277])^(a[345] & b[278])^(a[344] & b[279])^(a[343] & b[280])^(a[342] & b[281])^(a[341] & b[282])^(a[340] & b[283])^(a[339] & b[284])^(a[338] & b[285])^(a[337] & b[286])^(a[336] & b[287])^(a[335] & b[288])^(a[334] & b[289])^(a[333] & b[290])^(a[332] & b[291])^(a[331] & b[292])^(a[330] & b[293])^(a[329] & b[294])^(a[328] & b[295])^(a[327] & b[296])^(a[326] & b[297])^(a[325] & b[298])^(a[324] & b[299])^(a[323] & b[300])^(a[322] & b[301])^(a[321] & b[302])^(a[320] & b[303])^(a[319] & b[304])^(a[318] & b[305])^(a[317] & b[306])^(a[316] & b[307])^(a[315] & b[308])^(a[314] & b[309])^(a[313] & b[310])^(a[312] & b[311])^(a[311] & b[312])^(a[310] & b[313])^(a[309] & b[314])^(a[308] & b[315])^(a[307] & b[316])^(a[306] & b[317])^(a[305] & b[318])^(a[304] & b[319])^(a[303] & b[320])^(a[302] & b[321])^(a[301] & b[322])^(a[300] & b[323])^(a[299] & b[324])^(a[298] & b[325])^(a[297] & b[326])^(a[296] & b[327])^(a[295] & b[328])^(a[294] & b[329])^(a[293] & b[330])^(a[292] & b[331])^(a[291] & b[332])^(a[290] & b[333])^(a[289] & b[334])^(a[288] & b[335])^(a[287] & b[336])^(a[286] & b[337])^(a[285] & b[338])^(a[284] & b[339])^(a[283] & b[340])^(a[282] & b[341])^(a[281] & b[342])^(a[280] & b[343])^(a[279] & b[344])^(a[278] & b[345])^(a[277] & b[346])^(a[276] & b[347])^(a[275] & b[348])^(a[274] & b[349])^(a[273] & b[350])^(a[272] & b[351])^(a[271] & b[352])^(a[270] & b[353])^(a[269] & b[354])^(a[268] & b[355])^(a[267] & b[356])^(a[266] & b[357])^(a[265] & b[358])^(a[264] & b[359])^(a[263] & b[360])^(a[262] & b[361])^(a[261] & b[362])^(a[260] & b[363])^(a[259] & b[364])^(a[258] & b[365])^(a[257] & b[366])^(a[256] & b[367])^(a[255] & b[368])^(a[254] & b[369])^(a[253] & b[370])^(a[252] & b[371])^(a[251] & b[372])^(a[250] & b[373])^(a[249] & b[374])^(a[248] & b[375])^(a[247] & b[376])^(a[246] & b[377])^(a[245] & b[378])^(a[244] & b[379])^(a[243] & b[380])^(a[242] & b[381])^(a[241] & b[382])^(a[240] & b[383])^(a[239] & b[384])^(a[238] & b[385])^(a[237] & b[386])^(a[236] & b[387])^(a[235] & b[388])^(a[234] & b[389])^(a[233] & b[390])^(a[232] & b[391])^(a[231] & b[392])^(a[230] & b[393])^(a[229] & b[394])^(a[228] & b[395])^(a[227] & b[396])^(a[226] & b[397])^(a[225] & b[398])^(a[224] & b[399])^(a[223] & b[400])^(a[222] & b[401])^(a[221] & b[402])^(a[220] & b[403])^(a[219] & b[404])^(a[218] & b[405])^(a[217] & b[406])^(a[216] & b[407])^(a[215] & b[408]);
assign y[624] = (a[408] & b[216])^(a[407] & b[217])^(a[406] & b[218])^(a[405] & b[219])^(a[404] & b[220])^(a[403] & b[221])^(a[402] & b[222])^(a[401] & b[223])^(a[400] & b[224])^(a[399] & b[225])^(a[398] & b[226])^(a[397] & b[227])^(a[396] & b[228])^(a[395] & b[229])^(a[394] & b[230])^(a[393] & b[231])^(a[392] & b[232])^(a[391] & b[233])^(a[390] & b[234])^(a[389] & b[235])^(a[388] & b[236])^(a[387] & b[237])^(a[386] & b[238])^(a[385] & b[239])^(a[384] & b[240])^(a[383] & b[241])^(a[382] & b[242])^(a[381] & b[243])^(a[380] & b[244])^(a[379] & b[245])^(a[378] & b[246])^(a[377] & b[247])^(a[376] & b[248])^(a[375] & b[249])^(a[374] & b[250])^(a[373] & b[251])^(a[372] & b[252])^(a[371] & b[253])^(a[370] & b[254])^(a[369] & b[255])^(a[368] & b[256])^(a[367] & b[257])^(a[366] & b[258])^(a[365] & b[259])^(a[364] & b[260])^(a[363] & b[261])^(a[362] & b[262])^(a[361] & b[263])^(a[360] & b[264])^(a[359] & b[265])^(a[358] & b[266])^(a[357] & b[267])^(a[356] & b[268])^(a[355] & b[269])^(a[354] & b[270])^(a[353] & b[271])^(a[352] & b[272])^(a[351] & b[273])^(a[350] & b[274])^(a[349] & b[275])^(a[348] & b[276])^(a[347] & b[277])^(a[346] & b[278])^(a[345] & b[279])^(a[344] & b[280])^(a[343] & b[281])^(a[342] & b[282])^(a[341] & b[283])^(a[340] & b[284])^(a[339] & b[285])^(a[338] & b[286])^(a[337] & b[287])^(a[336] & b[288])^(a[335] & b[289])^(a[334] & b[290])^(a[333] & b[291])^(a[332] & b[292])^(a[331] & b[293])^(a[330] & b[294])^(a[329] & b[295])^(a[328] & b[296])^(a[327] & b[297])^(a[326] & b[298])^(a[325] & b[299])^(a[324] & b[300])^(a[323] & b[301])^(a[322] & b[302])^(a[321] & b[303])^(a[320] & b[304])^(a[319] & b[305])^(a[318] & b[306])^(a[317] & b[307])^(a[316] & b[308])^(a[315] & b[309])^(a[314] & b[310])^(a[313] & b[311])^(a[312] & b[312])^(a[311] & b[313])^(a[310] & b[314])^(a[309] & b[315])^(a[308] & b[316])^(a[307] & b[317])^(a[306] & b[318])^(a[305] & b[319])^(a[304] & b[320])^(a[303] & b[321])^(a[302] & b[322])^(a[301] & b[323])^(a[300] & b[324])^(a[299] & b[325])^(a[298] & b[326])^(a[297] & b[327])^(a[296] & b[328])^(a[295] & b[329])^(a[294] & b[330])^(a[293] & b[331])^(a[292] & b[332])^(a[291] & b[333])^(a[290] & b[334])^(a[289] & b[335])^(a[288] & b[336])^(a[287] & b[337])^(a[286] & b[338])^(a[285] & b[339])^(a[284] & b[340])^(a[283] & b[341])^(a[282] & b[342])^(a[281] & b[343])^(a[280] & b[344])^(a[279] & b[345])^(a[278] & b[346])^(a[277] & b[347])^(a[276] & b[348])^(a[275] & b[349])^(a[274] & b[350])^(a[273] & b[351])^(a[272] & b[352])^(a[271] & b[353])^(a[270] & b[354])^(a[269] & b[355])^(a[268] & b[356])^(a[267] & b[357])^(a[266] & b[358])^(a[265] & b[359])^(a[264] & b[360])^(a[263] & b[361])^(a[262] & b[362])^(a[261] & b[363])^(a[260] & b[364])^(a[259] & b[365])^(a[258] & b[366])^(a[257] & b[367])^(a[256] & b[368])^(a[255] & b[369])^(a[254] & b[370])^(a[253] & b[371])^(a[252] & b[372])^(a[251] & b[373])^(a[250] & b[374])^(a[249] & b[375])^(a[248] & b[376])^(a[247] & b[377])^(a[246] & b[378])^(a[245] & b[379])^(a[244] & b[380])^(a[243] & b[381])^(a[242] & b[382])^(a[241] & b[383])^(a[240] & b[384])^(a[239] & b[385])^(a[238] & b[386])^(a[237] & b[387])^(a[236] & b[388])^(a[235] & b[389])^(a[234] & b[390])^(a[233] & b[391])^(a[232] & b[392])^(a[231] & b[393])^(a[230] & b[394])^(a[229] & b[395])^(a[228] & b[396])^(a[227] & b[397])^(a[226] & b[398])^(a[225] & b[399])^(a[224] & b[400])^(a[223] & b[401])^(a[222] & b[402])^(a[221] & b[403])^(a[220] & b[404])^(a[219] & b[405])^(a[218] & b[406])^(a[217] & b[407])^(a[216] & b[408]);
assign y[625] = (a[408] & b[217])^(a[407] & b[218])^(a[406] & b[219])^(a[405] & b[220])^(a[404] & b[221])^(a[403] & b[222])^(a[402] & b[223])^(a[401] & b[224])^(a[400] & b[225])^(a[399] & b[226])^(a[398] & b[227])^(a[397] & b[228])^(a[396] & b[229])^(a[395] & b[230])^(a[394] & b[231])^(a[393] & b[232])^(a[392] & b[233])^(a[391] & b[234])^(a[390] & b[235])^(a[389] & b[236])^(a[388] & b[237])^(a[387] & b[238])^(a[386] & b[239])^(a[385] & b[240])^(a[384] & b[241])^(a[383] & b[242])^(a[382] & b[243])^(a[381] & b[244])^(a[380] & b[245])^(a[379] & b[246])^(a[378] & b[247])^(a[377] & b[248])^(a[376] & b[249])^(a[375] & b[250])^(a[374] & b[251])^(a[373] & b[252])^(a[372] & b[253])^(a[371] & b[254])^(a[370] & b[255])^(a[369] & b[256])^(a[368] & b[257])^(a[367] & b[258])^(a[366] & b[259])^(a[365] & b[260])^(a[364] & b[261])^(a[363] & b[262])^(a[362] & b[263])^(a[361] & b[264])^(a[360] & b[265])^(a[359] & b[266])^(a[358] & b[267])^(a[357] & b[268])^(a[356] & b[269])^(a[355] & b[270])^(a[354] & b[271])^(a[353] & b[272])^(a[352] & b[273])^(a[351] & b[274])^(a[350] & b[275])^(a[349] & b[276])^(a[348] & b[277])^(a[347] & b[278])^(a[346] & b[279])^(a[345] & b[280])^(a[344] & b[281])^(a[343] & b[282])^(a[342] & b[283])^(a[341] & b[284])^(a[340] & b[285])^(a[339] & b[286])^(a[338] & b[287])^(a[337] & b[288])^(a[336] & b[289])^(a[335] & b[290])^(a[334] & b[291])^(a[333] & b[292])^(a[332] & b[293])^(a[331] & b[294])^(a[330] & b[295])^(a[329] & b[296])^(a[328] & b[297])^(a[327] & b[298])^(a[326] & b[299])^(a[325] & b[300])^(a[324] & b[301])^(a[323] & b[302])^(a[322] & b[303])^(a[321] & b[304])^(a[320] & b[305])^(a[319] & b[306])^(a[318] & b[307])^(a[317] & b[308])^(a[316] & b[309])^(a[315] & b[310])^(a[314] & b[311])^(a[313] & b[312])^(a[312] & b[313])^(a[311] & b[314])^(a[310] & b[315])^(a[309] & b[316])^(a[308] & b[317])^(a[307] & b[318])^(a[306] & b[319])^(a[305] & b[320])^(a[304] & b[321])^(a[303] & b[322])^(a[302] & b[323])^(a[301] & b[324])^(a[300] & b[325])^(a[299] & b[326])^(a[298] & b[327])^(a[297] & b[328])^(a[296] & b[329])^(a[295] & b[330])^(a[294] & b[331])^(a[293] & b[332])^(a[292] & b[333])^(a[291] & b[334])^(a[290] & b[335])^(a[289] & b[336])^(a[288] & b[337])^(a[287] & b[338])^(a[286] & b[339])^(a[285] & b[340])^(a[284] & b[341])^(a[283] & b[342])^(a[282] & b[343])^(a[281] & b[344])^(a[280] & b[345])^(a[279] & b[346])^(a[278] & b[347])^(a[277] & b[348])^(a[276] & b[349])^(a[275] & b[350])^(a[274] & b[351])^(a[273] & b[352])^(a[272] & b[353])^(a[271] & b[354])^(a[270] & b[355])^(a[269] & b[356])^(a[268] & b[357])^(a[267] & b[358])^(a[266] & b[359])^(a[265] & b[360])^(a[264] & b[361])^(a[263] & b[362])^(a[262] & b[363])^(a[261] & b[364])^(a[260] & b[365])^(a[259] & b[366])^(a[258] & b[367])^(a[257] & b[368])^(a[256] & b[369])^(a[255] & b[370])^(a[254] & b[371])^(a[253] & b[372])^(a[252] & b[373])^(a[251] & b[374])^(a[250] & b[375])^(a[249] & b[376])^(a[248] & b[377])^(a[247] & b[378])^(a[246] & b[379])^(a[245] & b[380])^(a[244] & b[381])^(a[243] & b[382])^(a[242] & b[383])^(a[241] & b[384])^(a[240] & b[385])^(a[239] & b[386])^(a[238] & b[387])^(a[237] & b[388])^(a[236] & b[389])^(a[235] & b[390])^(a[234] & b[391])^(a[233] & b[392])^(a[232] & b[393])^(a[231] & b[394])^(a[230] & b[395])^(a[229] & b[396])^(a[228] & b[397])^(a[227] & b[398])^(a[226] & b[399])^(a[225] & b[400])^(a[224] & b[401])^(a[223] & b[402])^(a[222] & b[403])^(a[221] & b[404])^(a[220] & b[405])^(a[219] & b[406])^(a[218] & b[407])^(a[217] & b[408]);
assign y[626] = (a[408] & b[218])^(a[407] & b[219])^(a[406] & b[220])^(a[405] & b[221])^(a[404] & b[222])^(a[403] & b[223])^(a[402] & b[224])^(a[401] & b[225])^(a[400] & b[226])^(a[399] & b[227])^(a[398] & b[228])^(a[397] & b[229])^(a[396] & b[230])^(a[395] & b[231])^(a[394] & b[232])^(a[393] & b[233])^(a[392] & b[234])^(a[391] & b[235])^(a[390] & b[236])^(a[389] & b[237])^(a[388] & b[238])^(a[387] & b[239])^(a[386] & b[240])^(a[385] & b[241])^(a[384] & b[242])^(a[383] & b[243])^(a[382] & b[244])^(a[381] & b[245])^(a[380] & b[246])^(a[379] & b[247])^(a[378] & b[248])^(a[377] & b[249])^(a[376] & b[250])^(a[375] & b[251])^(a[374] & b[252])^(a[373] & b[253])^(a[372] & b[254])^(a[371] & b[255])^(a[370] & b[256])^(a[369] & b[257])^(a[368] & b[258])^(a[367] & b[259])^(a[366] & b[260])^(a[365] & b[261])^(a[364] & b[262])^(a[363] & b[263])^(a[362] & b[264])^(a[361] & b[265])^(a[360] & b[266])^(a[359] & b[267])^(a[358] & b[268])^(a[357] & b[269])^(a[356] & b[270])^(a[355] & b[271])^(a[354] & b[272])^(a[353] & b[273])^(a[352] & b[274])^(a[351] & b[275])^(a[350] & b[276])^(a[349] & b[277])^(a[348] & b[278])^(a[347] & b[279])^(a[346] & b[280])^(a[345] & b[281])^(a[344] & b[282])^(a[343] & b[283])^(a[342] & b[284])^(a[341] & b[285])^(a[340] & b[286])^(a[339] & b[287])^(a[338] & b[288])^(a[337] & b[289])^(a[336] & b[290])^(a[335] & b[291])^(a[334] & b[292])^(a[333] & b[293])^(a[332] & b[294])^(a[331] & b[295])^(a[330] & b[296])^(a[329] & b[297])^(a[328] & b[298])^(a[327] & b[299])^(a[326] & b[300])^(a[325] & b[301])^(a[324] & b[302])^(a[323] & b[303])^(a[322] & b[304])^(a[321] & b[305])^(a[320] & b[306])^(a[319] & b[307])^(a[318] & b[308])^(a[317] & b[309])^(a[316] & b[310])^(a[315] & b[311])^(a[314] & b[312])^(a[313] & b[313])^(a[312] & b[314])^(a[311] & b[315])^(a[310] & b[316])^(a[309] & b[317])^(a[308] & b[318])^(a[307] & b[319])^(a[306] & b[320])^(a[305] & b[321])^(a[304] & b[322])^(a[303] & b[323])^(a[302] & b[324])^(a[301] & b[325])^(a[300] & b[326])^(a[299] & b[327])^(a[298] & b[328])^(a[297] & b[329])^(a[296] & b[330])^(a[295] & b[331])^(a[294] & b[332])^(a[293] & b[333])^(a[292] & b[334])^(a[291] & b[335])^(a[290] & b[336])^(a[289] & b[337])^(a[288] & b[338])^(a[287] & b[339])^(a[286] & b[340])^(a[285] & b[341])^(a[284] & b[342])^(a[283] & b[343])^(a[282] & b[344])^(a[281] & b[345])^(a[280] & b[346])^(a[279] & b[347])^(a[278] & b[348])^(a[277] & b[349])^(a[276] & b[350])^(a[275] & b[351])^(a[274] & b[352])^(a[273] & b[353])^(a[272] & b[354])^(a[271] & b[355])^(a[270] & b[356])^(a[269] & b[357])^(a[268] & b[358])^(a[267] & b[359])^(a[266] & b[360])^(a[265] & b[361])^(a[264] & b[362])^(a[263] & b[363])^(a[262] & b[364])^(a[261] & b[365])^(a[260] & b[366])^(a[259] & b[367])^(a[258] & b[368])^(a[257] & b[369])^(a[256] & b[370])^(a[255] & b[371])^(a[254] & b[372])^(a[253] & b[373])^(a[252] & b[374])^(a[251] & b[375])^(a[250] & b[376])^(a[249] & b[377])^(a[248] & b[378])^(a[247] & b[379])^(a[246] & b[380])^(a[245] & b[381])^(a[244] & b[382])^(a[243] & b[383])^(a[242] & b[384])^(a[241] & b[385])^(a[240] & b[386])^(a[239] & b[387])^(a[238] & b[388])^(a[237] & b[389])^(a[236] & b[390])^(a[235] & b[391])^(a[234] & b[392])^(a[233] & b[393])^(a[232] & b[394])^(a[231] & b[395])^(a[230] & b[396])^(a[229] & b[397])^(a[228] & b[398])^(a[227] & b[399])^(a[226] & b[400])^(a[225] & b[401])^(a[224] & b[402])^(a[223] & b[403])^(a[222] & b[404])^(a[221] & b[405])^(a[220] & b[406])^(a[219] & b[407])^(a[218] & b[408]);
assign y[627] = (a[408] & b[219])^(a[407] & b[220])^(a[406] & b[221])^(a[405] & b[222])^(a[404] & b[223])^(a[403] & b[224])^(a[402] & b[225])^(a[401] & b[226])^(a[400] & b[227])^(a[399] & b[228])^(a[398] & b[229])^(a[397] & b[230])^(a[396] & b[231])^(a[395] & b[232])^(a[394] & b[233])^(a[393] & b[234])^(a[392] & b[235])^(a[391] & b[236])^(a[390] & b[237])^(a[389] & b[238])^(a[388] & b[239])^(a[387] & b[240])^(a[386] & b[241])^(a[385] & b[242])^(a[384] & b[243])^(a[383] & b[244])^(a[382] & b[245])^(a[381] & b[246])^(a[380] & b[247])^(a[379] & b[248])^(a[378] & b[249])^(a[377] & b[250])^(a[376] & b[251])^(a[375] & b[252])^(a[374] & b[253])^(a[373] & b[254])^(a[372] & b[255])^(a[371] & b[256])^(a[370] & b[257])^(a[369] & b[258])^(a[368] & b[259])^(a[367] & b[260])^(a[366] & b[261])^(a[365] & b[262])^(a[364] & b[263])^(a[363] & b[264])^(a[362] & b[265])^(a[361] & b[266])^(a[360] & b[267])^(a[359] & b[268])^(a[358] & b[269])^(a[357] & b[270])^(a[356] & b[271])^(a[355] & b[272])^(a[354] & b[273])^(a[353] & b[274])^(a[352] & b[275])^(a[351] & b[276])^(a[350] & b[277])^(a[349] & b[278])^(a[348] & b[279])^(a[347] & b[280])^(a[346] & b[281])^(a[345] & b[282])^(a[344] & b[283])^(a[343] & b[284])^(a[342] & b[285])^(a[341] & b[286])^(a[340] & b[287])^(a[339] & b[288])^(a[338] & b[289])^(a[337] & b[290])^(a[336] & b[291])^(a[335] & b[292])^(a[334] & b[293])^(a[333] & b[294])^(a[332] & b[295])^(a[331] & b[296])^(a[330] & b[297])^(a[329] & b[298])^(a[328] & b[299])^(a[327] & b[300])^(a[326] & b[301])^(a[325] & b[302])^(a[324] & b[303])^(a[323] & b[304])^(a[322] & b[305])^(a[321] & b[306])^(a[320] & b[307])^(a[319] & b[308])^(a[318] & b[309])^(a[317] & b[310])^(a[316] & b[311])^(a[315] & b[312])^(a[314] & b[313])^(a[313] & b[314])^(a[312] & b[315])^(a[311] & b[316])^(a[310] & b[317])^(a[309] & b[318])^(a[308] & b[319])^(a[307] & b[320])^(a[306] & b[321])^(a[305] & b[322])^(a[304] & b[323])^(a[303] & b[324])^(a[302] & b[325])^(a[301] & b[326])^(a[300] & b[327])^(a[299] & b[328])^(a[298] & b[329])^(a[297] & b[330])^(a[296] & b[331])^(a[295] & b[332])^(a[294] & b[333])^(a[293] & b[334])^(a[292] & b[335])^(a[291] & b[336])^(a[290] & b[337])^(a[289] & b[338])^(a[288] & b[339])^(a[287] & b[340])^(a[286] & b[341])^(a[285] & b[342])^(a[284] & b[343])^(a[283] & b[344])^(a[282] & b[345])^(a[281] & b[346])^(a[280] & b[347])^(a[279] & b[348])^(a[278] & b[349])^(a[277] & b[350])^(a[276] & b[351])^(a[275] & b[352])^(a[274] & b[353])^(a[273] & b[354])^(a[272] & b[355])^(a[271] & b[356])^(a[270] & b[357])^(a[269] & b[358])^(a[268] & b[359])^(a[267] & b[360])^(a[266] & b[361])^(a[265] & b[362])^(a[264] & b[363])^(a[263] & b[364])^(a[262] & b[365])^(a[261] & b[366])^(a[260] & b[367])^(a[259] & b[368])^(a[258] & b[369])^(a[257] & b[370])^(a[256] & b[371])^(a[255] & b[372])^(a[254] & b[373])^(a[253] & b[374])^(a[252] & b[375])^(a[251] & b[376])^(a[250] & b[377])^(a[249] & b[378])^(a[248] & b[379])^(a[247] & b[380])^(a[246] & b[381])^(a[245] & b[382])^(a[244] & b[383])^(a[243] & b[384])^(a[242] & b[385])^(a[241] & b[386])^(a[240] & b[387])^(a[239] & b[388])^(a[238] & b[389])^(a[237] & b[390])^(a[236] & b[391])^(a[235] & b[392])^(a[234] & b[393])^(a[233] & b[394])^(a[232] & b[395])^(a[231] & b[396])^(a[230] & b[397])^(a[229] & b[398])^(a[228] & b[399])^(a[227] & b[400])^(a[226] & b[401])^(a[225] & b[402])^(a[224] & b[403])^(a[223] & b[404])^(a[222] & b[405])^(a[221] & b[406])^(a[220] & b[407])^(a[219] & b[408]);
assign y[628] = (a[408] & b[220])^(a[407] & b[221])^(a[406] & b[222])^(a[405] & b[223])^(a[404] & b[224])^(a[403] & b[225])^(a[402] & b[226])^(a[401] & b[227])^(a[400] & b[228])^(a[399] & b[229])^(a[398] & b[230])^(a[397] & b[231])^(a[396] & b[232])^(a[395] & b[233])^(a[394] & b[234])^(a[393] & b[235])^(a[392] & b[236])^(a[391] & b[237])^(a[390] & b[238])^(a[389] & b[239])^(a[388] & b[240])^(a[387] & b[241])^(a[386] & b[242])^(a[385] & b[243])^(a[384] & b[244])^(a[383] & b[245])^(a[382] & b[246])^(a[381] & b[247])^(a[380] & b[248])^(a[379] & b[249])^(a[378] & b[250])^(a[377] & b[251])^(a[376] & b[252])^(a[375] & b[253])^(a[374] & b[254])^(a[373] & b[255])^(a[372] & b[256])^(a[371] & b[257])^(a[370] & b[258])^(a[369] & b[259])^(a[368] & b[260])^(a[367] & b[261])^(a[366] & b[262])^(a[365] & b[263])^(a[364] & b[264])^(a[363] & b[265])^(a[362] & b[266])^(a[361] & b[267])^(a[360] & b[268])^(a[359] & b[269])^(a[358] & b[270])^(a[357] & b[271])^(a[356] & b[272])^(a[355] & b[273])^(a[354] & b[274])^(a[353] & b[275])^(a[352] & b[276])^(a[351] & b[277])^(a[350] & b[278])^(a[349] & b[279])^(a[348] & b[280])^(a[347] & b[281])^(a[346] & b[282])^(a[345] & b[283])^(a[344] & b[284])^(a[343] & b[285])^(a[342] & b[286])^(a[341] & b[287])^(a[340] & b[288])^(a[339] & b[289])^(a[338] & b[290])^(a[337] & b[291])^(a[336] & b[292])^(a[335] & b[293])^(a[334] & b[294])^(a[333] & b[295])^(a[332] & b[296])^(a[331] & b[297])^(a[330] & b[298])^(a[329] & b[299])^(a[328] & b[300])^(a[327] & b[301])^(a[326] & b[302])^(a[325] & b[303])^(a[324] & b[304])^(a[323] & b[305])^(a[322] & b[306])^(a[321] & b[307])^(a[320] & b[308])^(a[319] & b[309])^(a[318] & b[310])^(a[317] & b[311])^(a[316] & b[312])^(a[315] & b[313])^(a[314] & b[314])^(a[313] & b[315])^(a[312] & b[316])^(a[311] & b[317])^(a[310] & b[318])^(a[309] & b[319])^(a[308] & b[320])^(a[307] & b[321])^(a[306] & b[322])^(a[305] & b[323])^(a[304] & b[324])^(a[303] & b[325])^(a[302] & b[326])^(a[301] & b[327])^(a[300] & b[328])^(a[299] & b[329])^(a[298] & b[330])^(a[297] & b[331])^(a[296] & b[332])^(a[295] & b[333])^(a[294] & b[334])^(a[293] & b[335])^(a[292] & b[336])^(a[291] & b[337])^(a[290] & b[338])^(a[289] & b[339])^(a[288] & b[340])^(a[287] & b[341])^(a[286] & b[342])^(a[285] & b[343])^(a[284] & b[344])^(a[283] & b[345])^(a[282] & b[346])^(a[281] & b[347])^(a[280] & b[348])^(a[279] & b[349])^(a[278] & b[350])^(a[277] & b[351])^(a[276] & b[352])^(a[275] & b[353])^(a[274] & b[354])^(a[273] & b[355])^(a[272] & b[356])^(a[271] & b[357])^(a[270] & b[358])^(a[269] & b[359])^(a[268] & b[360])^(a[267] & b[361])^(a[266] & b[362])^(a[265] & b[363])^(a[264] & b[364])^(a[263] & b[365])^(a[262] & b[366])^(a[261] & b[367])^(a[260] & b[368])^(a[259] & b[369])^(a[258] & b[370])^(a[257] & b[371])^(a[256] & b[372])^(a[255] & b[373])^(a[254] & b[374])^(a[253] & b[375])^(a[252] & b[376])^(a[251] & b[377])^(a[250] & b[378])^(a[249] & b[379])^(a[248] & b[380])^(a[247] & b[381])^(a[246] & b[382])^(a[245] & b[383])^(a[244] & b[384])^(a[243] & b[385])^(a[242] & b[386])^(a[241] & b[387])^(a[240] & b[388])^(a[239] & b[389])^(a[238] & b[390])^(a[237] & b[391])^(a[236] & b[392])^(a[235] & b[393])^(a[234] & b[394])^(a[233] & b[395])^(a[232] & b[396])^(a[231] & b[397])^(a[230] & b[398])^(a[229] & b[399])^(a[228] & b[400])^(a[227] & b[401])^(a[226] & b[402])^(a[225] & b[403])^(a[224] & b[404])^(a[223] & b[405])^(a[222] & b[406])^(a[221] & b[407])^(a[220] & b[408]);
assign y[629] = (a[408] & b[221])^(a[407] & b[222])^(a[406] & b[223])^(a[405] & b[224])^(a[404] & b[225])^(a[403] & b[226])^(a[402] & b[227])^(a[401] & b[228])^(a[400] & b[229])^(a[399] & b[230])^(a[398] & b[231])^(a[397] & b[232])^(a[396] & b[233])^(a[395] & b[234])^(a[394] & b[235])^(a[393] & b[236])^(a[392] & b[237])^(a[391] & b[238])^(a[390] & b[239])^(a[389] & b[240])^(a[388] & b[241])^(a[387] & b[242])^(a[386] & b[243])^(a[385] & b[244])^(a[384] & b[245])^(a[383] & b[246])^(a[382] & b[247])^(a[381] & b[248])^(a[380] & b[249])^(a[379] & b[250])^(a[378] & b[251])^(a[377] & b[252])^(a[376] & b[253])^(a[375] & b[254])^(a[374] & b[255])^(a[373] & b[256])^(a[372] & b[257])^(a[371] & b[258])^(a[370] & b[259])^(a[369] & b[260])^(a[368] & b[261])^(a[367] & b[262])^(a[366] & b[263])^(a[365] & b[264])^(a[364] & b[265])^(a[363] & b[266])^(a[362] & b[267])^(a[361] & b[268])^(a[360] & b[269])^(a[359] & b[270])^(a[358] & b[271])^(a[357] & b[272])^(a[356] & b[273])^(a[355] & b[274])^(a[354] & b[275])^(a[353] & b[276])^(a[352] & b[277])^(a[351] & b[278])^(a[350] & b[279])^(a[349] & b[280])^(a[348] & b[281])^(a[347] & b[282])^(a[346] & b[283])^(a[345] & b[284])^(a[344] & b[285])^(a[343] & b[286])^(a[342] & b[287])^(a[341] & b[288])^(a[340] & b[289])^(a[339] & b[290])^(a[338] & b[291])^(a[337] & b[292])^(a[336] & b[293])^(a[335] & b[294])^(a[334] & b[295])^(a[333] & b[296])^(a[332] & b[297])^(a[331] & b[298])^(a[330] & b[299])^(a[329] & b[300])^(a[328] & b[301])^(a[327] & b[302])^(a[326] & b[303])^(a[325] & b[304])^(a[324] & b[305])^(a[323] & b[306])^(a[322] & b[307])^(a[321] & b[308])^(a[320] & b[309])^(a[319] & b[310])^(a[318] & b[311])^(a[317] & b[312])^(a[316] & b[313])^(a[315] & b[314])^(a[314] & b[315])^(a[313] & b[316])^(a[312] & b[317])^(a[311] & b[318])^(a[310] & b[319])^(a[309] & b[320])^(a[308] & b[321])^(a[307] & b[322])^(a[306] & b[323])^(a[305] & b[324])^(a[304] & b[325])^(a[303] & b[326])^(a[302] & b[327])^(a[301] & b[328])^(a[300] & b[329])^(a[299] & b[330])^(a[298] & b[331])^(a[297] & b[332])^(a[296] & b[333])^(a[295] & b[334])^(a[294] & b[335])^(a[293] & b[336])^(a[292] & b[337])^(a[291] & b[338])^(a[290] & b[339])^(a[289] & b[340])^(a[288] & b[341])^(a[287] & b[342])^(a[286] & b[343])^(a[285] & b[344])^(a[284] & b[345])^(a[283] & b[346])^(a[282] & b[347])^(a[281] & b[348])^(a[280] & b[349])^(a[279] & b[350])^(a[278] & b[351])^(a[277] & b[352])^(a[276] & b[353])^(a[275] & b[354])^(a[274] & b[355])^(a[273] & b[356])^(a[272] & b[357])^(a[271] & b[358])^(a[270] & b[359])^(a[269] & b[360])^(a[268] & b[361])^(a[267] & b[362])^(a[266] & b[363])^(a[265] & b[364])^(a[264] & b[365])^(a[263] & b[366])^(a[262] & b[367])^(a[261] & b[368])^(a[260] & b[369])^(a[259] & b[370])^(a[258] & b[371])^(a[257] & b[372])^(a[256] & b[373])^(a[255] & b[374])^(a[254] & b[375])^(a[253] & b[376])^(a[252] & b[377])^(a[251] & b[378])^(a[250] & b[379])^(a[249] & b[380])^(a[248] & b[381])^(a[247] & b[382])^(a[246] & b[383])^(a[245] & b[384])^(a[244] & b[385])^(a[243] & b[386])^(a[242] & b[387])^(a[241] & b[388])^(a[240] & b[389])^(a[239] & b[390])^(a[238] & b[391])^(a[237] & b[392])^(a[236] & b[393])^(a[235] & b[394])^(a[234] & b[395])^(a[233] & b[396])^(a[232] & b[397])^(a[231] & b[398])^(a[230] & b[399])^(a[229] & b[400])^(a[228] & b[401])^(a[227] & b[402])^(a[226] & b[403])^(a[225] & b[404])^(a[224] & b[405])^(a[223] & b[406])^(a[222] & b[407])^(a[221] & b[408]);
assign y[630] = (a[408] & b[222])^(a[407] & b[223])^(a[406] & b[224])^(a[405] & b[225])^(a[404] & b[226])^(a[403] & b[227])^(a[402] & b[228])^(a[401] & b[229])^(a[400] & b[230])^(a[399] & b[231])^(a[398] & b[232])^(a[397] & b[233])^(a[396] & b[234])^(a[395] & b[235])^(a[394] & b[236])^(a[393] & b[237])^(a[392] & b[238])^(a[391] & b[239])^(a[390] & b[240])^(a[389] & b[241])^(a[388] & b[242])^(a[387] & b[243])^(a[386] & b[244])^(a[385] & b[245])^(a[384] & b[246])^(a[383] & b[247])^(a[382] & b[248])^(a[381] & b[249])^(a[380] & b[250])^(a[379] & b[251])^(a[378] & b[252])^(a[377] & b[253])^(a[376] & b[254])^(a[375] & b[255])^(a[374] & b[256])^(a[373] & b[257])^(a[372] & b[258])^(a[371] & b[259])^(a[370] & b[260])^(a[369] & b[261])^(a[368] & b[262])^(a[367] & b[263])^(a[366] & b[264])^(a[365] & b[265])^(a[364] & b[266])^(a[363] & b[267])^(a[362] & b[268])^(a[361] & b[269])^(a[360] & b[270])^(a[359] & b[271])^(a[358] & b[272])^(a[357] & b[273])^(a[356] & b[274])^(a[355] & b[275])^(a[354] & b[276])^(a[353] & b[277])^(a[352] & b[278])^(a[351] & b[279])^(a[350] & b[280])^(a[349] & b[281])^(a[348] & b[282])^(a[347] & b[283])^(a[346] & b[284])^(a[345] & b[285])^(a[344] & b[286])^(a[343] & b[287])^(a[342] & b[288])^(a[341] & b[289])^(a[340] & b[290])^(a[339] & b[291])^(a[338] & b[292])^(a[337] & b[293])^(a[336] & b[294])^(a[335] & b[295])^(a[334] & b[296])^(a[333] & b[297])^(a[332] & b[298])^(a[331] & b[299])^(a[330] & b[300])^(a[329] & b[301])^(a[328] & b[302])^(a[327] & b[303])^(a[326] & b[304])^(a[325] & b[305])^(a[324] & b[306])^(a[323] & b[307])^(a[322] & b[308])^(a[321] & b[309])^(a[320] & b[310])^(a[319] & b[311])^(a[318] & b[312])^(a[317] & b[313])^(a[316] & b[314])^(a[315] & b[315])^(a[314] & b[316])^(a[313] & b[317])^(a[312] & b[318])^(a[311] & b[319])^(a[310] & b[320])^(a[309] & b[321])^(a[308] & b[322])^(a[307] & b[323])^(a[306] & b[324])^(a[305] & b[325])^(a[304] & b[326])^(a[303] & b[327])^(a[302] & b[328])^(a[301] & b[329])^(a[300] & b[330])^(a[299] & b[331])^(a[298] & b[332])^(a[297] & b[333])^(a[296] & b[334])^(a[295] & b[335])^(a[294] & b[336])^(a[293] & b[337])^(a[292] & b[338])^(a[291] & b[339])^(a[290] & b[340])^(a[289] & b[341])^(a[288] & b[342])^(a[287] & b[343])^(a[286] & b[344])^(a[285] & b[345])^(a[284] & b[346])^(a[283] & b[347])^(a[282] & b[348])^(a[281] & b[349])^(a[280] & b[350])^(a[279] & b[351])^(a[278] & b[352])^(a[277] & b[353])^(a[276] & b[354])^(a[275] & b[355])^(a[274] & b[356])^(a[273] & b[357])^(a[272] & b[358])^(a[271] & b[359])^(a[270] & b[360])^(a[269] & b[361])^(a[268] & b[362])^(a[267] & b[363])^(a[266] & b[364])^(a[265] & b[365])^(a[264] & b[366])^(a[263] & b[367])^(a[262] & b[368])^(a[261] & b[369])^(a[260] & b[370])^(a[259] & b[371])^(a[258] & b[372])^(a[257] & b[373])^(a[256] & b[374])^(a[255] & b[375])^(a[254] & b[376])^(a[253] & b[377])^(a[252] & b[378])^(a[251] & b[379])^(a[250] & b[380])^(a[249] & b[381])^(a[248] & b[382])^(a[247] & b[383])^(a[246] & b[384])^(a[245] & b[385])^(a[244] & b[386])^(a[243] & b[387])^(a[242] & b[388])^(a[241] & b[389])^(a[240] & b[390])^(a[239] & b[391])^(a[238] & b[392])^(a[237] & b[393])^(a[236] & b[394])^(a[235] & b[395])^(a[234] & b[396])^(a[233] & b[397])^(a[232] & b[398])^(a[231] & b[399])^(a[230] & b[400])^(a[229] & b[401])^(a[228] & b[402])^(a[227] & b[403])^(a[226] & b[404])^(a[225] & b[405])^(a[224] & b[406])^(a[223] & b[407])^(a[222] & b[408]);
assign y[631] = (a[408] & b[223])^(a[407] & b[224])^(a[406] & b[225])^(a[405] & b[226])^(a[404] & b[227])^(a[403] & b[228])^(a[402] & b[229])^(a[401] & b[230])^(a[400] & b[231])^(a[399] & b[232])^(a[398] & b[233])^(a[397] & b[234])^(a[396] & b[235])^(a[395] & b[236])^(a[394] & b[237])^(a[393] & b[238])^(a[392] & b[239])^(a[391] & b[240])^(a[390] & b[241])^(a[389] & b[242])^(a[388] & b[243])^(a[387] & b[244])^(a[386] & b[245])^(a[385] & b[246])^(a[384] & b[247])^(a[383] & b[248])^(a[382] & b[249])^(a[381] & b[250])^(a[380] & b[251])^(a[379] & b[252])^(a[378] & b[253])^(a[377] & b[254])^(a[376] & b[255])^(a[375] & b[256])^(a[374] & b[257])^(a[373] & b[258])^(a[372] & b[259])^(a[371] & b[260])^(a[370] & b[261])^(a[369] & b[262])^(a[368] & b[263])^(a[367] & b[264])^(a[366] & b[265])^(a[365] & b[266])^(a[364] & b[267])^(a[363] & b[268])^(a[362] & b[269])^(a[361] & b[270])^(a[360] & b[271])^(a[359] & b[272])^(a[358] & b[273])^(a[357] & b[274])^(a[356] & b[275])^(a[355] & b[276])^(a[354] & b[277])^(a[353] & b[278])^(a[352] & b[279])^(a[351] & b[280])^(a[350] & b[281])^(a[349] & b[282])^(a[348] & b[283])^(a[347] & b[284])^(a[346] & b[285])^(a[345] & b[286])^(a[344] & b[287])^(a[343] & b[288])^(a[342] & b[289])^(a[341] & b[290])^(a[340] & b[291])^(a[339] & b[292])^(a[338] & b[293])^(a[337] & b[294])^(a[336] & b[295])^(a[335] & b[296])^(a[334] & b[297])^(a[333] & b[298])^(a[332] & b[299])^(a[331] & b[300])^(a[330] & b[301])^(a[329] & b[302])^(a[328] & b[303])^(a[327] & b[304])^(a[326] & b[305])^(a[325] & b[306])^(a[324] & b[307])^(a[323] & b[308])^(a[322] & b[309])^(a[321] & b[310])^(a[320] & b[311])^(a[319] & b[312])^(a[318] & b[313])^(a[317] & b[314])^(a[316] & b[315])^(a[315] & b[316])^(a[314] & b[317])^(a[313] & b[318])^(a[312] & b[319])^(a[311] & b[320])^(a[310] & b[321])^(a[309] & b[322])^(a[308] & b[323])^(a[307] & b[324])^(a[306] & b[325])^(a[305] & b[326])^(a[304] & b[327])^(a[303] & b[328])^(a[302] & b[329])^(a[301] & b[330])^(a[300] & b[331])^(a[299] & b[332])^(a[298] & b[333])^(a[297] & b[334])^(a[296] & b[335])^(a[295] & b[336])^(a[294] & b[337])^(a[293] & b[338])^(a[292] & b[339])^(a[291] & b[340])^(a[290] & b[341])^(a[289] & b[342])^(a[288] & b[343])^(a[287] & b[344])^(a[286] & b[345])^(a[285] & b[346])^(a[284] & b[347])^(a[283] & b[348])^(a[282] & b[349])^(a[281] & b[350])^(a[280] & b[351])^(a[279] & b[352])^(a[278] & b[353])^(a[277] & b[354])^(a[276] & b[355])^(a[275] & b[356])^(a[274] & b[357])^(a[273] & b[358])^(a[272] & b[359])^(a[271] & b[360])^(a[270] & b[361])^(a[269] & b[362])^(a[268] & b[363])^(a[267] & b[364])^(a[266] & b[365])^(a[265] & b[366])^(a[264] & b[367])^(a[263] & b[368])^(a[262] & b[369])^(a[261] & b[370])^(a[260] & b[371])^(a[259] & b[372])^(a[258] & b[373])^(a[257] & b[374])^(a[256] & b[375])^(a[255] & b[376])^(a[254] & b[377])^(a[253] & b[378])^(a[252] & b[379])^(a[251] & b[380])^(a[250] & b[381])^(a[249] & b[382])^(a[248] & b[383])^(a[247] & b[384])^(a[246] & b[385])^(a[245] & b[386])^(a[244] & b[387])^(a[243] & b[388])^(a[242] & b[389])^(a[241] & b[390])^(a[240] & b[391])^(a[239] & b[392])^(a[238] & b[393])^(a[237] & b[394])^(a[236] & b[395])^(a[235] & b[396])^(a[234] & b[397])^(a[233] & b[398])^(a[232] & b[399])^(a[231] & b[400])^(a[230] & b[401])^(a[229] & b[402])^(a[228] & b[403])^(a[227] & b[404])^(a[226] & b[405])^(a[225] & b[406])^(a[224] & b[407])^(a[223] & b[408]);
assign y[632] = (a[408] & b[224])^(a[407] & b[225])^(a[406] & b[226])^(a[405] & b[227])^(a[404] & b[228])^(a[403] & b[229])^(a[402] & b[230])^(a[401] & b[231])^(a[400] & b[232])^(a[399] & b[233])^(a[398] & b[234])^(a[397] & b[235])^(a[396] & b[236])^(a[395] & b[237])^(a[394] & b[238])^(a[393] & b[239])^(a[392] & b[240])^(a[391] & b[241])^(a[390] & b[242])^(a[389] & b[243])^(a[388] & b[244])^(a[387] & b[245])^(a[386] & b[246])^(a[385] & b[247])^(a[384] & b[248])^(a[383] & b[249])^(a[382] & b[250])^(a[381] & b[251])^(a[380] & b[252])^(a[379] & b[253])^(a[378] & b[254])^(a[377] & b[255])^(a[376] & b[256])^(a[375] & b[257])^(a[374] & b[258])^(a[373] & b[259])^(a[372] & b[260])^(a[371] & b[261])^(a[370] & b[262])^(a[369] & b[263])^(a[368] & b[264])^(a[367] & b[265])^(a[366] & b[266])^(a[365] & b[267])^(a[364] & b[268])^(a[363] & b[269])^(a[362] & b[270])^(a[361] & b[271])^(a[360] & b[272])^(a[359] & b[273])^(a[358] & b[274])^(a[357] & b[275])^(a[356] & b[276])^(a[355] & b[277])^(a[354] & b[278])^(a[353] & b[279])^(a[352] & b[280])^(a[351] & b[281])^(a[350] & b[282])^(a[349] & b[283])^(a[348] & b[284])^(a[347] & b[285])^(a[346] & b[286])^(a[345] & b[287])^(a[344] & b[288])^(a[343] & b[289])^(a[342] & b[290])^(a[341] & b[291])^(a[340] & b[292])^(a[339] & b[293])^(a[338] & b[294])^(a[337] & b[295])^(a[336] & b[296])^(a[335] & b[297])^(a[334] & b[298])^(a[333] & b[299])^(a[332] & b[300])^(a[331] & b[301])^(a[330] & b[302])^(a[329] & b[303])^(a[328] & b[304])^(a[327] & b[305])^(a[326] & b[306])^(a[325] & b[307])^(a[324] & b[308])^(a[323] & b[309])^(a[322] & b[310])^(a[321] & b[311])^(a[320] & b[312])^(a[319] & b[313])^(a[318] & b[314])^(a[317] & b[315])^(a[316] & b[316])^(a[315] & b[317])^(a[314] & b[318])^(a[313] & b[319])^(a[312] & b[320])^(a[311] & b[321])^(a[310] & b[322])^(a[309] & b[323])^(a[308] & b[324])^(a[307] & b[325])^(a[306] & b[326])^(a[305] & b[327])^(a[304] & b[328])^(a[303] & b[329])^(a[302] & b[330])^(a[301] & b[331])^(a[300] & b[332])^(a[299] & b[333])^(a[298] & b[334])^(a[297] & b[335])^(a[296] & b[336])^(a[295] & b[337])^(a[294] & b[338])^(a[293] & b[339])^(a[292] & b[340])^(a[291] & b[341])^(a[290] & b[342])^(a[289] & b[343])^(a[288] & b[344])^(a[287] & b[345])^(a[286] & b[346])^(a[285] & b[347])^(a[284] & b[348])^(a[283] & b[349])^(a[282] & b[350])^(a[281] & b[351])^(a[280] & b[352])^(a[279] & b[353])^(a[278] & b[354])^(a[277] & b[355])^(a[276] & b[356])^(a[275] & b[357])^(a[274] & b[358])^(a[273] & b[359])^(a[272] & b[360])^(a[271] & b[361])^(a[270] & b[362])^(a[269] & b[363])^(a[268] & b[364])^(a[267] & b[365])^(a[266] & b[366])^(a[265] & b[367])^(a[264] & b[368])^(a[263] & b[369])^(a[262] & b[370])^(a[261] & b[371])^(a[260] & b[372])^(a[259] & b[373])^(a[258] & b[374])^(a[257] & b[375])^(a[256] & b[376])^(a[255] & b[377])^(a[254] & b[378])^(a[253] & b[379])^(a[252] & b[380])^(a[251] & b[381])^(a[250] & b[382])^(a[249] & b[383])^(a[248] & b[384])^(a[247] & b[385])^(a[246] & b[386])^(a[245] & b[387])^(a[244] & b[388])^(a[243] & b[389])^(a[242] & b[390])^(a[241] & b[391])^(a[240] & b[392])^(a[239] & b[393])^(a[238] & b[394])^(a[237] & b[395])^(a[236] & b[396])^(a[235] & b[397])^(a[234] & b[398])^(a[233] & b[399])^(a[232] & b[400])^(a[231] & b[401])^(a[230] & b[402])^(a[229] & b[403])^(a[228] & b[404])^(a[227] & b[405])^(a[226] & b[406])^(a[225] & b[407])^(a[224] & b[408]);
assign y[633] = (a[408] & b[225])^(a[407] & b[226])^(a[406] & b[227])^(a[405] & b[228])^(a[404] & b[229])^(a[403] & b[230])^(a[402] & b[231])^(a[401] & b[232])^(a[400] & b[233])^(a[399] & b[234])^(a[398] & b[235])^(a[397] & b[236])^(a[396] & b[237])^(a[395] & b[238])^(a[394] & b[239])^(a[393] & b[240])^(a[392] & b[241])^(a[391] & b[242])^(a[390] & b[243])^(a[389] & b[244])^(a[388] & b[245])^(a[387] & b[246])^(a[386] & b[247])^(a[385] & b[248])^(a[384] & b[249])^(a[383] & b[250])^(a[382] & b[251])^(a[381] & b[252])^(a[380] & b[253])^(a[379] & b[254])^(a[378] & b[255])^(a[377] & b[256])^(a[376] & b[257])^(a[375] & b[258])^(a[374] & b[259])^(a[373] & b[260])^(a[372] & b[261])^(a[371] & b[262])^(a[370] & b[263])^(a[369] & b[264])^(a[368] & b[265])^(a[367] & b[266])^(a[366] & b[267])^(a[365] & b[268])^(a[364] & b[269])^(a[363] & b[270])^(a[362] & b[271])^(a[361] & b[272])^(a[360] & b[273])^(a[359] & b[274])^(a[358] & b[275])^(a[357] & b[276])^(a[356] & b[277])^(a[355] & b[278])^(a[354] & b[279])^(a[353] & b[280])^(a[352] & b[281])^(a[351] & b[282])^(a[350] & b[283])^(a[349] & b[284])^(a[348] & b[285])^(a[347] & b[286])^(a[346] & b[287])^(a[345] & b[288])^(a[344] & b[289])^(a[343] & b[290])^(a[342] & b[291])^(a[341] & b[292])^(a[340] & b[293])^(a[339] & b[294])^(a[338] & b[295])^(a[337] & b[296])^(a[336] & b[297])^(a[335] & b[298])^(a[334] & b[299])^(a[333] & b[300])^(a[332] & b[301])^(a[331] & b[302])^(a[330] & b[303])^(a[329] & b[304])^(a[328] & b[305])^(a[327] & b[306])^(a[326] & b[307])^(a[325] & b[308])^(a[324] & b[309])^(a[323] & b[310])^(a[322] & b[311])^(a[321] & b[312])^(a[320] & b[313])^(a[319] & b[314])^(a[318] & b[315])^(a[317] & b[316])^(a[316] & b[317])^(a[315] & b[318])^(a[314] & b[319])^(a[313] & b[320])^(a[312] & b[321])^(a[311] & b[322])^(a[310] & b[323])^(a[309] & b[324])^(a[308] & b[325])^(a[307] & b[326])^(a[306] & b[327])^(a[305] & b[328])^(a[304] & b[329])^(a[303] & b[330])^(a[302] & b[331])^(a[301] & b[332])^(a[300] & b[333])^(a[299] & b[334])^(a[298] & b[335])^(a[297] & b[336])^(a[296] & b[337])^(a[295] & b[338])^(a[294] & b[339])^(a[293] & b[340])^(a[292] & b[341])^(a[291] & b[342])^(a[290] & b[343])^(a[289] & b[344])^(a[288] & b[345])^(a[287] & b[346])^(a[286] & b[347])^(a[285] & b[348])^(a[284] & b[349])^(a[283] & b[350])^(a[282] & b[351])^(a[281] & b[352])^(a[280] & b[353])^(a[279] & b[354])^(a[278] & b[355])^(a[277] & b[356])^(a[276] & b[357])^(a[275] & b[358])^(a[274] & b[359])^(a[273] & b[360])^(a[272] & b[361])^(a[271] & b[362])^(a[270] & b[363])^(a[269] & b[364])^(a[268] & b[365])^(a[267] & b[366])^(a[266] & b[367])^(a[265] & b[368])^(a[264] & b[369])^(a[263] & b[370])^(a[262] & b[371])^(a[261] & b[372])^(a[260] & b[373])^(a[259] & b[374])^(a[258] & b[375])^(a[257] & b[376])^(a[256] & b[377])^(a[255] & b[378])^(a[254] & b[379])^(a[253] & b[380])^(a[252] & b[381])^(a[251] & b[382])^(a[250] & b[383])^(a[249] & b[384])^(a[248] & b[385])^(a[247] & b[386])^(a[246] & b[387])^(a[245] & b[388])^(a[244] & b[389])^(a[243] & b[390])^(a[242] & b[391])^(a[241] & b[392])^(a[240] & b[393])^(a[239] & b[394])^(a[238] & b[395])^(a[237] & b[396])^(a[236] & b[397])^(a[235] & b[398])^(a[234] & b[399])^(a[233] & b[400])^(a[232] & b[401])^(a[231] & b[402])^(a[230] & b[403])^(a[229] & b[404])^(a[228] & b[405])^(a[227] & b[406])^(a[226] & b[407])^(a[225] & b[408]);
assign y[634] = (a[408] & b[226])^(a[407] & b[227])^(a[406] & b[228])^(a[405] & b[229])^(a[404] & b[230])^(a[403] & b[231])^(a[402] & b[232])^(a[401] & b[233])^(a[400] & b[234])^(a[399] & b[235])^(a[398] & b[236])^(a[397] & b[237])^(a[396] & b[238])^(a[395] & b[239])^(a[394] & b[240])^(a[393] & b[241])^(a[392] & b[242])^(a[391] & b[243])^(a[390] & b[244])^(a[389] & b[245])^(a[388] & b[246])^(a[387] & b[247])^(a[386] & b[248])^(a[385] & b[249])^(a[384] & b[250])^(a[383] & b[251])^(a[382] & b[252])^(a[381] & b[253])^(a[380] & b[254])^(a[379] & b[255])^(a[378] & b[256])^(a[377] & b[257])^(a[376] & b[258])^(a[375] & b[259])^(a[374] & b[260])^(a[373] & b[261])^(a[372] & b[262])^(a[371] & b[263])^(a[370] & b[264])^(a[369] & b[265])^(a[368] & b[266])^(a[367] & b[267])^(a[366] & b[268])^(a[365] & b[269])^(a[364] & b[270])^(a[363] & b[271])^(a[362] & b[272])^(a[361] & b[273])^(a[360] & b[274])^(a[359] & b[275])^(a[358] & b[276])^(a[357] & b[277])^(a[356] & b[278])^(a[355] & b[279])^(a[354] & b[280])^(a[353] & b[281])^(a[352] & b[282])^(a[351] & b[283])^(a[350] & b[284])^(a[349] & b[285])^(a[348] & b[286])^(a[347] & b[287])^(a[346] & b[288])^(a[345] & b[289])^(a[344] & b[290])^(a[343] & b[291])^(a[342] & b[292])^(a[341] & b[293])^(a[340] & b[294])^(a[339] & b[295])^(a[338] & b[296])^(a[337] & b[297])^(a[336] & b[298])^(a[335] & b[299])^(a[334] & b[300])^(a[333] & b[301])^(a[332] & b[302])^(a[331] & b[303])^(a[330] & b[304])^(a[329] & b[305])^(a[328] & b[306])^(a[327] & b[307])^(a[326] & b[308])^(a[325] & b[309])^(a[324] & b[310])^(a[323] & b[311])^(a[322] & b[312])^(a[321] & b[313])^(a[320] & b[314])^(a[319] & b[315])^(a[318] & b[316])^(a[317] & b[317])^(a[316] & b[318])^(a[315] & b[319])^(a[314] & b[320])^(a[313] & b[321])^(a[312] & b[322])^(a[311] & b[323])^(a[310] & b[324])^(a[309] & b[325])^(a[308] & b[326])^(a[307] & b[327])^(a[306] & b[328])^(a[305] & b[329])^(a[304] & b[330])^(a[303] & b[331])^(a[302] & b[332])^(a[301] & b[333])^(a[300] & b[334])^(a[299] & b[335])^(a[298] & b[336])^(a[297] & b[337])^(a[296] & b[338])^(a[295] & b[339])^(a[294] & b[340])^(a[293] & b[341])^(a[292] & b[342])^(a[291] & b[343])^(a[290] & b[344])^(a[289] & b[345])^(a[288] & b[346])^(a[287] & b[347])^(a[286] & b[348])^(a[285] & b[349])^(a[284] & b[350])^(a[283] & b[351])^(a[282] & b[352])^(a[281] & b[353])^(a[280] & b[354])^(a[279] & b[355])^(a[278] & b[356])^(a[277] & b[357])^(a[276] & b[358])^(a[275] & b[359])^(a[274] & b[360])^(a[273] & b[361])^(a[272] & b[362])^(a[271] & b[363])^(a[270] & b[364])^(a[269] & b[365])^(a[268] & b[366])^(a[267] & b[367])^(a[266] & b[368])^(a[265] & b[369])^(a[264] & b[370])^(a[263] & b[371])^(a[262] & b[372])^(a[261] & b[373])^(a[260] & b[374])^(a[259] & b[375])^(a[258] & b[376])^(a[257] & b[377])^(a[256] & b[378])^(a[255] & b[379])^(a[254] & b[380])^(a[253] & b[381])^(a[252] & b[382])^(a[251] & b[383])^(a[250] & b[384])^(a[249] & b[385])^(a[248] & b[386])^(a[247] & b[387])^(a[246] & b[388])^(a[245] & b[389])^(a[244] & b[390])^(a[243] & b[391])^(a[242] & b[392])^(a[241] & b[393])^(a[240] & b[394])^(a[239] & b[395])^(a[238] & b[396])^(a[237] & b[397])^(a[236] & b[398])^(a[235] & b[399])^(a[234] & b[400])^(a[233] & b[401])^(a[232] & b[402])^(a[231] & b[403])^(a[230] & b[404])^(a[229] & b[405])^(a[228] & b[406])^(a[227] & b[407])^(a[226] & b[408]);
assign y[635] = (a[408] & b[227])^(a[407] & b[228])^(a[406] & b[229])^(a[405] & b[230])^(a[404] & b[231])^(a[403] & b[232])^(a[402] & b[233])^(a[401] & b[234])^(a[400] & b[235])^(a[399] & b[236])^(a[398] & b[237])^(a[397] & b[238])^(a[396] & b[239])^(a[395] & b[240])^(a[394] & b[241])^(a[393] & b[242])^(a[392] & b[243])^(a[391] & b[244])^(a[390] & b[245])^(a[389] & b[246])^(a[388] & b[247])^(a[387] & b[248])^(a[386] & b[249])^(a[385] & b[250])^(a[384] & b[251])^(a[383] & b[252])^(a[382] & b[253])^(a[381] & b[254])^(a[380] & b[255])^(a[379] & b[256])^(a[378] & b[257])^(a[377] & b[258])^(a[376] & b[259])^(a[375] & b[260])^(a[374] & b[261])^(a[373] & b[262])^(a[372] & b[263])^(a[371] & b[264])^(a[370] & b[265])^(a[369] & b[266])^(a[368] & b[267])^(a[367] & b[268])^(a[366] & b[269])^(a[365] & b[270])^(a[364] & b[271])^(a[363] & b[272])^(a[362] & b[273])^(a[361] & b[274])^(a[360] & b[275])^(a[359] & b[276])^(a[358] & b[277])^(a[357] & b[278])^(a[356] & b[279])^(a[355] & b[280])^(a[354] & b[281])^(a[353] & b[282])^(a[352] & b[283])^(a[351] & b[284])^(a[350] & b[285])^(a[349] & b[286])^(a[348] & b[287])^(a[347] & b[288])^(a[346] & b[289])^(a[345] & b[290])^(a[344] & b[291])^(a[343] & b[292])^(a[342] & b[293])^(a[341] & b[294])^(a[340] & b[295])^(a[339] & b[296])^(a[338] & b[297])^(a[337] & b[298])^(a[336] & b[299])^(a[335] & b[300])^(a[334] & b[301])^(a[333] & b[302])^(a[332] & b[303])^(a[331] & b[304])^(a[330] & b[305])^(a[329] & b[306])^(a[328] & b[307])^(a[327] & b[308])^(a[326] & b[309])^(a[325] & b[310])^(a[324] & b[311])^(a[323] & b[312])^(a[322] & b[313])^(a[321] & b[314])^(a[320] & b[315])^(a[319] & b[316])^(a[318] & b[317])^(a[317] & b[318])^(a[316] & b[319])^(a[315] & b[320])^(a[314] & b[321])^(a[313] & b[322])^(a[312] & b[323])^(a[311] & b[324])^(a[310] & b[325])^(a[309] & b[326])^(a[308] & b[327])^(a[307] & b[328])^(a[306] & b[329])^(a[305] & b[330])^(a[304] & b[331])^(a[303] & b[332])^(a[302] & b[333])^(a[301] & b[334])^(a[300] & b[335])^(a[299] & b[336])^(a[298] & b[337])^(a[297] & b[338])^(a[296] & b[339])^(a[295] & b[340])^(a[294] & b[341])^(a[293] & b[342])^(a[292] & b[343])^(a[291] & b[344])^(a[290] & b[345])^(a[289] & b[346])^(a[288] & b[347])^(a[287] & b[348])^(a[286] & b[349])^(a[285] & b[350])^(a[284] & b[351])^(a[283] & b[352])^(a[282] & b[353])^(a[281] & b[354])^(a[280] & b[355])^(a[279] & b[356])^(a[278] & b[357])^(a[277] & b[358])^(a[276] & b[359])^(a[275] & b[360])^(a[274] & b[361])^(a[273] & b[362])^(a[272] & b[363])^(a[271] & b[364])^(a[270] & b[365])^(a[269] & b[366])^(a[268] & b[367])^(a[267] & b[368])^(a[266] & b[369])^(a[265] & b[370])^(a[264] & b[371])^(a[263] & b[372])^(a[262] & b[373])^(a[261] & b[374])^(a[260] & b[375])^(a[259] & b[376])^(a[258] & b[377])^(a[257] & b[378])^(a[256] & b[379])^(a[255] & b[380])^(a[254] & b[381])^(a[253] & b[382])^(a[252] & b[383])^(a[251] & b[384])^(a[250] & b[385])^(a[249] & b[386])^(a[248] & b[387])^(a[247] & b[388])^(a[246] & b[389])^(a[245] & b[390])^(a[244] & b[391])^(a[243] & b[392])^(a[242] & b[393])^(a[241] & b[394])^(a[240] & b[395])^(a[239] & b[396])^(a[238] & b[397])^(a[237] & b[398])^(a[236] & b[399])^(a[235] & b[400])^(a[234] & b[401])^(a[233] & b[402])^(a[232] & b[403])^(a[231] & b[404])^(a[230] & b[405])^(a[229] & b[406])^(a[228] & b[407])^(a[227] & b[408]);
assign y[636] = (a[408] & b[228])^(a[407] & b[229])^(a[406] & b[230])^(a[405] & b[231])^(a[404] & b[232])^(a[403] & b[233])^(a[402] & b[234])^(a[401] & b[235])^(a[400] & b[236])^(a[399] & b[237])^(a[398] & b[238])^(a[397] & b[239])^(a[396] & b[240])^(a[395] & b[241])^(a[394] & b[242])^(a[393] & b[243])^(a[392] & b[244])^(a[391] & b[245])^(a[390] & b[246])^(a[389] & b[247])^(a[388] & b[248])^(a[387] & b[249])^(a[386] & b[250])^(a[385] & b[251])^(a[384] & b[252])^(a[383] & b[253])^(a[382] & b[254])^(a[381] & b[255])^(a[380] & b[256])^(a[379] & b[257])^(a[378] & b[258])^(a[377] & b[259])^(a[376] & b[260])^(a[375] & b[261])^(a[374] & b[262])^(a[373] & b[263])^(a[372] & b[264])^(a[371] & b[265])^(a[370] & b[266])^(a[369] & b[267])^(a[368] & b[268])^(a[367] & b[269])^(a[366] & b[270])^(a[365] & b[271])^(a[364] & b[272])^(a[363] & b[273])^(a[362] & b[274])^(a[361] & b[275])^(a[360] & b[276])^(a[359] & b[277])^(a[358] & b[278])^(a[357] & b[279])^(a[356] & b[280])^(a[355] & b[281])^(a[354] & b[282])^(a[353] & b[283])^(a[352] & b[284])^(a[351] & b[285])^(a[350] & b[286])^(a[349] & b[287])^(a[348] & b[288])^(a[347] & b[289])^(a[346] & b[290])^(a[345] & b[291])^(a[344] & b[292])^(a[343] & b[293])^(a[342] & b[294])^(a[341] & b[295])^(a[340] & b[296])^(a[339] & b[297])^(a[338] & b[298])^(a[337] & b[299])^(a[336] & b[300])^(a[335] & b[301])^(a[334] & b[302])^(a[333] & b[303])^(a[332] & b[304])^(a[331] & b[305])^(a[330] & b[306])^(a[329] & b[307])^(a[328] & b[308])^(a[327] & b[309])^(a[326] & b[310])^(a[325] & b[311])^(a[324] & b[312])^(a[323] & b[313])^(a[322] & b[314])^(a[321] & b[315])^(a[320] & b[316])^(a[319] & b[317])^(a[318] & b[318])^(a[317] & b[319])^(a[316] & b[320])^(a[315] & b[321])^(a[314] & b[322])^(a[313] & b[323])^(a[312] & b[324])^(a[311] & b[325])^(a[310] & b[326])^(a[309] & b[327])^(a[308] & b[328])^(a[307] & b[329])^(a[306] & b[330])^(a[305] & b[331])^(a[304] & b[332])^(a[303] & b[333])^(a[302] & b[334])^(a[301] & b[335])^(a[300] & b[336])^(a[299] & b[337])^(a[298] & b[338])^(a[297] & b[339])^(a[296] & b[340])^(a[295] & b[341])^(a[294] & b[342])^(a[293] & b[343])^(a[292] & b[344])^(a[291] & b[345])^(a[290] & b[346])^(a[289] & b[347])^(a[288] & b[348])^(a[287] & b[349])^(a[286] & b[350])^(a[285] & b[351])^(a[284] & b[352])^(a[283] & b[353])^(a[282] & b[354])^(a[281] & b[355])^(a[280] & b[356])^(a[279] & b[357])^(a[278] & b[358])^(a[277] & b[359])^(a[276] & b[360])^(a[275] & b[361])^(a[274] & b[362])^(a[273] & b[363])^(a[272] & b[364])^(a[271] & b[365])^(a[270] & b[366])^(a[269] & b[367])^(a[268] & b[368])^(a[267] & b[369])^(a[266] & b[370])^(a[265] & b[371])^(a[264] & b[372])^(a[263] & b[373])^(a[262] & b[374])^(a[261] & b[375])^(a[260] & b[376])^(a[259] & b[377])^(a[258] & b[378])^(a[257] & b[379])^(a[256] & b[380])^(a[255] & b[381])^(a[254] & b[382])^(a[253] & b[383])^(a[252] & b[384])^(a[251] & b[385])^(a[250] & b[386])^(a[249] & b[387])^(a[248] & b[388])^(a[247] & b[389])^(a[246] & b[390])^(a[245] & b[391])^(a[244] & b[392])^(a[243] & b[393])^(a[242] & b[394])^(a[241] & b[395])^(a[240] & b[396])^(a[239] & b[397])^(a[238] & b[398])^(a[237] & b[399])^(a[236] & b[400])^(a[235] & b[401])^(a[234] & b[402])^(a[233] & b[403])^(a[232] & b[404])^(a[231] & b[405])^(a[230] & b[406])^(a[229] & b[407])^(a[228] & b[408]);
assign y[637] = (a[408] & b[229])^(a[407] & b[230])^(a[406] & b[231])^(a[405] & b[232])^(a[404] & b[233])^(a[403] & b[234])^(a[402] & b[235])^(a[401] & b[236])^(a[400] & b[237])^(a[399] & b[238])^(a[398] & b[239])^(a[397] & b[240])^(a[396] & b[241])^(a[395] & b[242])^(a[394] & b[243])^(a[393] & b[244])^(a[392] & b[245])^(a[391] & b[246])^(a[390] & b[247])^(a[389] & b[248])^(a[388] & b[249])^(a[387] & b[250])^(a[386] & b[251])^(a[385] & b[252])^(a[384] & b[253])^(a[383] & b[254])^(a[382] & b[255])^(a[381] & b[256])^(a[380] & b[257])^(a[379] & b[258])^(a[378] & b[259])^(a[377] & b[260])^(a[376] & b[261])^(a[375] & b[262])^(a[374] & b[263])^(a[373] & b[264])^(a[372] & b[265])^(a[371] & b[266])^(a[370] & b[267])^(a[369] & b[268])^(a[368] & b[269])^(a[367] & b[270])^(a[366] & b[271])^(a[365] & b[272])^(a[364] & b[273])^(a[363] & b[274])^(a[362] & b[275])^(a[361] & b[276])^(a[360] & b[277])^(a[359] & b[278])^(a[358] & b[279])^(a[357] & b[280])^(a[356] & b[281])^(a[355] & b[282])^(a[354] & b[283])^(a[353] & b[284])^(a[352] & b[285])^(a[351] & b[286])^(a[350] & b[287])^(a[349] & b[288])^(a[348] & b[289])^(a[347] & b[290])^(a[346] & b[291])^(a[345] & b[292])^(a[344] & b[293])^(a[343] & b[294])^(a[342] & b[295])^(a[341] & b[296])^(a[340] & b[297])^(a[339] & b[298])^(a[338] & b[299])^(a[337] & b[300])^(a[336] & b[301])^(a[335] & b[302])^(a[334] & b[303])^(a[333] & b[304])^(a[332] & b[305])^(a[331] & b[306])^(a[330] & b[307])^(a[329] & b[308])^(a[328] & b[309])^(a[327] & b[310])^(a[326] & b[311])^(a[325] & b[312])^(a[324] & b[313])^(a[323] & b[314])^(a[322] & b[315])^(a[321] & b[316])^(a[320] & b[317])^(a[319] & b[318])^(a[318] & b[319])^(a[317] & b[320])^(a[316] & b[321])^(a[315] & b[322])^(a[314] & b[323])^(a[313] & b[324])^(a[312] & b[325])^(a[311] & b[326])^(a[310] & b[327])^(a[309] & b[328])^(a[308] & b[329])^(a[307] & b[330])^(a[306] & b[331])^(a[305] & b[332])^(a[304] & b[333])^(a[303] & b[334])^(a[302] & b[335])^(a[301] & b[336])^(a[300] & b[337])^(a[299] & b[338])^(a[298] & b[339])^(a[297] & b[340])^(a[296] & b[341])^(a[295] & b[342])^(a[294] & b[343])^(a[293] & b[344])^(a[292] & b[345])^(a[291] & b[346])^(a[290] & b[347])^(a[289] & b[348])^(a[288] & b[349])^(a[287] & b[350])^(a[286] & b[351])^(a[285] & b[352])^(a[284] & b[353])^(a[283] & b[354])^(a[282] & b[355])^(a[281] & b[356])^(a[280] & b[357])^(a[279] & b[358])^(a[278] & b[359])^(a[277] & b[360])^(a[276] & b[361])^(a[275] & b[362])^(a[274] & b[363])^(a[273] & b[364])^(a[272] & b[365])^(a[271] & b[366])^(a[270] & b[367])^(a[269] & b[368])^(a[268] & b[369])^(a[267] & b[370])^(a[266] & b[371])^(a[265] & b[372])^(a[264] & b[373])^(a[263] & b[374])^(a[262] & b[375])^(a[261] & b[376])^(a[260] & b[377])^(a[259] & b[378])^(a[258] & b[379])^(a[257] & b[380])^(a[256] & b[381])^(a[255] & b[382])^(a[254] & b[383])^(a[253] & b[384])^(a[252] & b[385])^(a[251] & b[386])^(a[250] & b[387])^(a[249] & b[388])^(a[248] & b[389])^(a[247] & b[390])^(a[246] & b[391])^(a[245] & b[392])^(a[244] & b[393])^(a[243] & b[394])^(a[242] & b[395])^(a[241] & b[396])^(a[240] & b[397])^(a[239] & b[398])^(a[238] & b[399])^(a[237] & b[400])^(a[236] & b[401])^(a[235] & b[402])^(a[234] & b[403])^(a[233] & b[404])^(a[232] & b[405])^(a[231] & b[406])^(a[230] & b[407])^(a[229] & b[408]);
assign y[638] = (a[408] & b[230])^(a[407] & b[231])^(a[406] & b[232])^(a[405] & b[233])^(a[404] & b[234])^(a[403] & b[235])^(a[402] & b[236])^(a[401] & b[237])^(a[400] & b[238])^(a[399] & b[239])^(a[398] & b[240])^(a[397] & b[241])^(a[396] & b[242])^(a[395] & b[243])^(a[394] & b[244])^(a[393] & b[245])^(a[392] & b[246])^(a[391] & b[247])^(a[390] & b[248])^(a[389] & b[249])^(a[388] & b[250])^(a[387] & b[251])^(a[386] & b[252])^(a[385] & b[253])^(a[384] & b[254])^(a[383] & b[255])^(a[382] & b[256])^(a[381] & b[257])^(a[380] & b[258])^(a[379] & b[259])^(a[378] & b[260])^(a[377] & b[261])^(a[376] & b[262])^(a[375] & b[263])^(a[374] & b[264])^(a[373] & b[265])^(a[372] & b[266])^(a[371] & b[267])^(a[370] & b[268])^(a[369] & b[269])^(a[368] & b[270])^(a[367] & b[271])^(a[366] & b[272])^(a[365] & b[273])^(a[364] & b[274])^(a[363] & b[275])^(a[362] & b[276])^(a[361] & b[277])^(a[360] & b[278])^(a[359] & b[279])^(a[358] & b[280])^(a[357] & b[281])^(a[356] & b[282])^(a[355] & b[283])^(a[354] & b[284])^(a[353] & b[285])^(a[352] & b[286])^(a[351] & b[287])^(a[350] & b[288])^(a[349] & b[289])^(a[348] & b[290])^(a[347] & b[291])^(a[346] & b[292])^(a[345] & b[293])^(a[344] & b[294])^(a[343] & b[295])^(a[342] & b[296])^(a[341] & b[297])^(a[340] & b[298])^(a[339] & b[299])^(a[338] & b[300])^(a[337] & b[301])^(a[336] & b[302])^(a[335] & b[303])^(a[334] & b[304])^(a[333] & b[305])^(a[332] & b[306])^(a[331] & b[307])^(a[330] & b[308])^(a[329] & b[309])^(a[328] & b[310])^(a[327] & b[311])^(a[326] & b[312])^(a[325] & b[313])^(a[324] & b[314])^(a[323] & b[315])^(a[322] & b[316])^(a[321] & b[317])^(a[320] & b[318])^(a[319] & b[319])^(a[318] & b[320])^(a[317] & b[321])^(a[316] & b[322])^(a[315] & b[323])^(a[314] & b[324])^(a[313] & b[325])^(a[312] & b[326])^(a[311] & b[327])^(a[310] & b[328])^(a[309] & b[329])^(a[308] & b[330])^(a[307] & b[331])^(a[306] & b[332])^(a[305] & b[333])^(a[304] & b[334])^(a[303] & b[335])^(a[302] & b[336])^(a[301] & b[337])^(a[300] & b[338])^(a[299] & b[339])^(a[298] & b[340])^(a[297] & b[341])^(a[296] & b[342])^(a[295] & b[343])^(a[294] & b[344])^(a[293] & b[345])^(a[292] & b[346])^(a[291] & b[347])^(a[290] & b[348])^(a[289] & b[349])^(a[288] & b[350])^(a[287] & b[351])^(a[286] & b[352])^(a[285] & b[353])^(a[284] & b[354])^(a[283] & b[355])^(a[282] & b[356])^(a[281] & b[357])^(a[280] & b[358])^(a[279] & b[359])^(a[278] & b[360])^(a[277] & b[361])^(a[276] & b[362])^(a[275] & b[363])^(a[274] & b[364])^(a[273] & b[365])^(a[272] & b[366])^(a[271] & b[367])^(a[270] & b[368])^(a[269] & b[369])^(a[268] & b[370])^(a[267] & b[371])^(a[266] & b[372])^(a[265] & b[373])^(a[264] & b[374])^(a[263] & b[375])^(a[262] & b[376])^(a[261] & b[377])^(a[260] & b[378])^(a[259] & b[379])^(a[258] & b[380])^(a[257] & b[381])^(a[256] & b[382])^(a[255] & b[383])^(a[254] & b[384])^(a[253] & b[385])^(a[252] & b[386])^(a[251] & b[387])^(a[250] & b[388])^(a[249] & b[389])^(a[248] & b[390])^(a[247] & b[391])^(a[246] & b[392])^(a[245] & b[393])^(a[244] & b[394])^(a[243] & b[395])^(a[242] & b[396])^(a[241] & b[397])^(a[240] & b[398])^(a[239] & b[399])^(a[238] & b[400])^(a[237] & b[401])^(a[236] & b[402])^(a[235] & b[403])^(a[234] & b[404])^(a[233] & b[405])^(a[232] & b[406])^(a[231] & b[407])^(a[230] & b[408]);
assign y[639] = (a[408] & b[231])^(a[407] & b[232])^(a[406] & b[233])^(a[405] & b[234])^(a[404] & b[235])^(a[403] & b[236])^(a[402] & b[237])^(a[401] & b[238])^(a[400] & b[239])^(a[399] & b[240])^(a[398] & b[241])^(a[397] & b[242])^(a[396] & b[243])^(a[395] & b[244])^(a[394] & b[245])^(a[393] & b[246])^(a[392] & b[247])^(a[391] & b[248])^(a[390] & b[249])^(a[389] & b[250])^(a[388] & b[251])^(a[387] & b[252])^(a[386] & b[253])^(a[385] & b[254])^(a[384] & b[255])^(a[383] & b[256])^(a[382] & b[257])^(a[381] & b[258])^(a[380] & b[259])^(a[379] & b[260])^(a[378] & b[261])^(a[377] & b[262])^(a[376] & b[263])^(a[375] & b[264])^(a[374] & b[265])^(a[373] & b[266])^(a[372] & b[267])^(a[371] & b[268])^(a[370] & b[269])^(a[369] & b[270])^(a[368] & b[271])^(a[367] & b[272])^(a[366] & b[273])^(a[365] & b[274])^(a[364] & b[275])^(a[363] & b[276])^(a[362] & b[277])^(a[361] & b[278])^(a[360] & b[279])^(a[359] & b[280])^(a[358] & b[281])^(a[357] & b[282])^(a[356] & b[283])^(a[355] & b[284])^(a[354] & b[285])^(a[353] & b[286])^(a[352] & b[287])^(a[351] & b[288])^(a[350] & b[289])^(a[349] & b[290])^(a[348] & b[291])^(a[347] & b[292])^(a[346] & b[293])^(a[345] & b[294])^(a[344] & b[295])^(a[343] & b[296])^(a[342] & b[297])^(a[341] & b[298])^(a[340] & b[299])^(a[339] & b[300])^(a[338] & b[301])^(a[337] & b[302])^(a[336] & b[303])^(a[335] & b[304])^(a[334] & b[305])^(a[333] & b[306])^(a[332] & b[307])^(a[331] & b[308])^(a[330] & b[309])^(a[329] & b[310])^(a[328] & b[311])^(a[327] & b[312])^(a[326] & b[313])^(a[325] & b[314])^(a[324] & b[315])^(a[323] & b[316])^(a[322] & b[317])^(a[321] & b[318])^(a[320] & b[319])^(a[319] & b[320])^(a[318] & b[321])^(a[317] & b[322])^(a[316] & b[323])^(a[315] & b[324])^(a[314] & b[325])^(a[313] & b[326])^(a[312] & b[327])^(a[311] & b[328])^(a[310] & b[329])^(a[309] & b[330])^(a[308] & b[331])^(a[307] & b[332])^(a[306] & b[333])^(a[305] & b[334])^(a[304] & b[335])^(a[303] & b[336])^(a[302] & b[337])^(a[301] & b[338])^(a[300] & b[339])^(a[299] & b[340])^(a[298] & b[341])^(a[297] & b[342])^(a[296] & b[343])^(a[295] & b[344])^(a[294] & b[345])^(a[293] & b[346])^(a[292] & b[347])^(a[291] & b[348])^(a[290] & b[349])^(a[289] & b[350])^(a[288] & b[351])^(a[287] & b[352])^(a[286] & b[353])^(a[285] & b[354])^(a[284] & b[355])^(a[283] & b[356])^(a[282] & b[357])^(a[281] & b[358])^(a[280] & b[359])^(a[279] & b[360])^(a[278] & b[361])^(a[277] & b[362])^(a[276] & b[363])^(a[275] & b[364])^(a[274] & b[365])^(a[273] & b[366])^(a[272] & b[367])^(a[271] & b[368])^(a[270] & b[369])^(a[269] & b[370])^(a[268] & b[371])^(a[267] & b[372])^(a[266] & b[373])^(a[265] & b[374])^(a[264] & b[375])^(a[263] & b[376])^(a[262] & b[377])^(a[261] & b[378])^(a[260] & b[379])^(a[259] & b[380])^(a[258] & b[381])^(a[257] & b[382])^(a[256] & b[383])^(a[255] & b[384])^(a[254] & b[385])^(a[253] & b[386])^(a[252] & b[387])^(a[251] & b[388])^(a[250] & b[389])^(a[249] & b[390])^(a[248] & b[391])^(a[247] & b[392])^(a[246] & b[393])^(a[245] & b[394])^(a[244] & b[395])^(a[243] & b[396])^(a[242] & b[397])^(a[241] & b[398])^(a[240] & b[399])^(a[239] & b[400])^(a[238] & b[401])^(a[237] & b[402])^(a[236] & b[403])^(a[235] & b[404])^(a[234] & b[405])^(a[233] & b[406])^(a[232] & b[407])^(a[231] & b[408]);
assign y[640] = (a[408] & b[232])^(a[407] & b[233])^(a[406] & b[234])^(a[405] & b[235])^(a[404] & b[236])^(a[403] & b[237])^(a[402] & b[238])^(a[401] & b[239])^(a[400] & b[240])^(a[399] & b[241])^(a[398] & b[242])^(a[397] & b[243])^(a[396] & b[244])^(a[395] & b[245])^(a[394] & b[246])^(a[393] & b[247])^(a[392] & b[248])^(a[391] & b[249])^(a[390] & b[250])^(a[389] & b[251])^(a[388] & b[252])^(a[387] & b[253])^(a[386] & b[254])^(a[385] & b[255])^(a[384] & b[256])^(a[383] & b[257])^(a[382] & b[258])^(a[381] & b[259])^(a[380] & b[260])^(a[379] & b[261])^(a[378] & b[262])^(a[377] & b[263])^(a[376] & b[264])^(a[375] & b[265])^(a[374] & b[266])^(a[373] & b[267])^(a[372] & b[268])^(a[371] & b[269])^(a[370] & b[270])^(a[369] & b[271])^(a[368] & b[272])^(a[367] & b[273])^(a[366] & b[274])^(a[365] & b[275])^(a[364] & b[276])^(a[363] & b[277])^(a[362] & b[278])^(a[361] & b[279])^(a[360] & b[280])^(a[359] & b[281])^(a[358] & b[282])^(a[357] & b[283])^(a[356] & b[284])^(a[355] & b[285])^(a[354] & b[286])^(a[353] & b[287])^(a[352] & b[288])^(a[351] & b[289])^(a[350] & b[290])^(a[349] & b[291])^(a[348] & b[292])^(a[347] & b[293])^(a[346] & b[294])^(a[345] & b[295])^(a[344] & b[296])^(a[343] & b[297])^(a[342] & b[298])^(a[341] & b[299])^(a[340] & b[300])^(a[339] & b[301])^(a[338] & b[302])^(a[337] & b[303])^(a[336] & b[304])^(a[335] & b[305])^(a[334] & b[306])^(a[333] & b[307])^(a[332] & b[308])^(a[331] & b[309])^(a[330] & b[310])^(a[329] & b[311])^(a[328] & b[312])^(a[327] & b[313])^(a[326] & b[314])^(a[325] & b[315])^(a[324] & b[316])^(a[323] & b[317])^(a[322] & b[318])^(a[321] & b[319])^(a[320] & b[320])^(a[319] & b[321])^(a[318] & b[322])^(a[317] & b[323])^(a[316] & b[324])^(a[315] & b[325])^(a[314] & b[326])^(a[313] & b[327])^(a[312] & b[328])^(a[311] & b[329])^(a[310] & b[330])^(a[309] & b[331])^(a[308] & b[332])^(a[307] & b[333])^(a[306] & b[334])^(a[305] & b[335])^(a[304] & b[336])^(a[303] & b[337])^(a[302] & b[338])^(a[301] & b[339])^(a[300] & b[340])^(a[299] & b[341])^(a[298] & b[342])^(a[297] & b[343])^(a[296] & b[344])^(a[295] & b[345])^(a[294] & b[346])^(a[293] & b[347])^(a[292] & b[348])^(a[291] & b[349])^(a[290] & b[350])^(a[289] & b[351])^(a[288] & b[352])^(a[287] & b[353])^(a[286] & b[354])^(a[285] & b[355])^(a[284] & b[356])^(a[283] & b[357])^(a[282] & b[358])^(a[281] & b[359])^(a[280] & b[360])^(a[279] & b[361])^(a[278] & b[362])^(a[277] & b[363])^(a[276] & b[364])^(a[275] & b[365])^(a[274] & b[366])^(a[273] & b[367])^(a[272] & b[368])^(a[271] & b[369])^(a[270] & b[370])^(a[269] & b[371])^(a[268] & b[372])^(a[267] & b[373])^(a[266] & b[374])^(a[265] & b[375])^(a[264] & b[376])^(a[263] & b[377])^(a[262] & b[378])^(a[261] & b[379])^(a[260] & b[380])^(a[259] & b[381])^(a[258] & b[382])^(a[257] & b[383])^(a[256] & b[384])^(a[255] & b[385])^(a[254] & b[386])^(a[253] & b[387])^(a[252] & b[388])^(a[251] & b[389])^(a[250] & b[390])^(a[249] & b[391])^(a[248] & b[392])^(a[247] & b[393])^(a[246] & b[394])^(a[245] & b[395])^(a[244] & b[396])^(a[243] & b[397])^(a[242] & b[398])^(a[241] & b[399])^(a[240] & b[400])^(a[239] & b[401])^(a[238] & b[402])^(a[237] & b[403])^(a[236] & b[404])^(a[235] & b[405])^(a[234] & b[406])^(a[233] & b[407])^(a[232] & b[408]);
assign y[641] = (a[408] & b[233])^(a[407] & b[234])^(a[406] & b[235])^(a[405] & b[236])^(a[404] & b[237])^(a[403] & b[238])^(a[402] & b[239])^(a[401] & b[240])^(a[400] & b[241])^(a[399] & b[242])^(a[398] & b[243])^(a[397] & b[244])^(a[396] & b[245])^(a[395] & b[246])^(a[394] & b[247])^(a[393] & b[248])^(a[392] & b[249])^(a[391] & b[250])^(a[390] & b[251])^(a[389] & b[252])^(a[388] & b[253])^(a[387] & b[254])^(a[386] & b[255])^(a[385] & b[256])^(a[384] & b[257])^(a[383] & b[258])^(a[382] & b[259])^(a[381] & b[260])^(a[380] & b[261])^(a[379] & b[262])^(a[378] & b[263])^(a[377] & b[264])^(a[376] & b[265])^(a[375] & b[266])^(a[374] & b[267])^(a[373] & b[268])^(a[372] & b[269])^(a[371] & b[270])^(a[370] & b[271])^(a[369] & b[272])^(a[368] & b[273])^(a[367] & b[274])^(a[366] & b[275])^(a[365] & b[276])^(a[364] & b[277])^(a[363] & b[278])^(a[362] & b[279])^(a[361] & b[280])^(a[360] & b[281])^(a[359] & b[282])^(a[358] & b[283])^(a[357] & b[284])^(a[356] & b[285])^(a[355] & b[286])^(a[354] & b[287])^(a[353] & b[288])^(a[352] & b[289])^(a[351] & b[290])^(a[350] & b[291])^(a[349] & b[292])^(a[348] & b[293])^(a[347] & b[294])^(a[346] & b[295])^(a[345] & b[296])^(a[344] & b[297])^(a[343] & b[298])^(a[342] & b[299])^(a[341] & b[300])^(a[340] & b[301])^(a[339] & b[302])^(a[338] & b[303])^(a[337] & b[304])^(a[336] & b[305])^(a[335] & b[306])^(a[334] & b[307])^(a[333] & b[308])^(a[332] & b[309])^(a[331] & b[310])^(a[330] & b[311])^(a[329] & b[312])^(a[328] & b[313])^(a[327] & b[314])^(a[326] & b[315])^(a[325] & b[316])^(a[324] & b[317])^(a[323] & b[318])^(a[322] & b[319])^(a[321] & b[320])^(a[320] & b[321])^(a[319] & b[322])^(a[318] & b[323])^(a[317] & b[324])^(a[316] & b[325])^(a[315] & b[326])^(a[314] & b[327])^(a[313] & b[328])^(a[312] & b[329])^(a[311] & b[330])^(a[310] & b[331])^(a[309] & b[332])^(a[308] & b[333])^(a[307] & b[334])^(a[306] & b[335])^(a[305] & b[336])^(a[304] & b[337])^(a[303] & b[338])^(a[302] & b[339])^(a[301] & b[340])^(a[300] & b[341])^(a[299] & b[342])^(a[298] & b[343])^(a[297] & b[344])^(a[296] & b[345])^(a[295] & b[346])^(a[294] & b[347])^(a[293] & b[348])^(a[292] & b[349])^(a[291] & b[350])^(a[290] & b[351])^(a[289] & b[352])^(a[288] & b[353])^(a[287] & b[354])^(a[286] & b[355])^(a[285] & b[356])^(a[284] & b[357])^(a[283] & b[358])^(a[282] & b[359])^(a[281] & b[360])^(a[280] & b[361])^(a[279] & b[362])^(a[278] & b[363])^(a[277] & b[364])^(a[276] & b[365])^(a[275] & b[366])^(a[274] & b[367])^(a[273] & b[368])^(a[272] & b[369])^(a[271] & b[370])^(a[270] & b[371])^(a[269] & b[372])^(a[268] & b[373])^(a[267] & b[374])^(a[266] & b[375])^(a[265] & b[376])^(a[264] & b[377])^(a[263] & b[378])^(a[262] & b[379])^(a[261] & b[380])^(a[260] & b[381])^(a[259] & b[382])^(a[258] & b[383])^(a[257] & b[384])^(a[256] & b[385])^(a[255] & b[386])^(a[254] & b[387])^(a[253] & b[388])^(a[252] & b[389])^(a[251] & b[390])^(a[250] & b[391])^(a[249] & b[392])^(a[248] & b[393])^(a[247] & b[394])^(a[246] & b[395])^(a[245] & b[396])^(a[244] & b[397])^(a[243] & b[398])^(a[242] & b[399])^(a[241] & b[400])^(a[240] & b[401])^(a[239] & b[402])^(a[238] & b[403])^(a[237] & b[404])^(a[236] & b[405])^(a[235] & b[406])^(a[234] & b[407])^(a[233] & b[408]);
assign y[642] = (a[408] & b[234])^(a[407] & b[235])^(a[406] & b[236])^(a[405] & b[237])^(a[404] & b[238])^(a[403] & b[239])^(a[402] & b[240])^(a[401] & b[241])^(a[400] & b[242])^(a[399] & b[243])^(a[398] & b[244])^(a[397] & b[245])^(a[396] & b[246])^(a[395] & b[247])^(a[394] & b[248])^(a[393] & b[249])^(a[392] & b[250])^(a[391] & b[251])^(a[390] & b[252])^(a[389] & b[253])^(a[388] & b[254])^(a[387] & b[255])^(a[386] & b[256])^(a[385] & b[257])^(a[384] & b[258])^(a[383] & b[259])^(a[382] & b[260])^(a[381] & b[261])^(a[380] & b[262])^(a[379] & b[263])^(a[378] & b[264])^(a[377] & b[265])^(a[376] & b[266])^(a[375] & b[267])^(a[374] & b[268])^(a[373] & b[269])^(a[372] & b[270])^(a[371] & b[271])^(a[370] & b[272])^(a[369] & b[273])^(a[368] & b[274])^(a[367] & b[275])^(a[366] & b[276])^(a[365] & b[277])^(a[364] & b[278])^(a[363] & b[279])^(a[362] & b[280])^(a[361] & b[281])^(a[360] & b[282])^(a[359] & b[283])^(a[358] & b[284])^(a[357] & b[285])^(a[356] & b[286])^(a[355] & b[287])^(a[354] & b[288])^(a[353] & b[289])^(a[352] & b[290])^(a[351] & b[291])^(a[350] & b[292])^(a[349] & b[293])^(a[348] & b[294])^(a[347] & b[295])^(a[346] & b[296])^(a[345] & b[297])^(a[344] & b[298])^(a[343] & b[299])^(a[342] & b[300])^(a[341] & b[301])^(a[340] & b[302])^(a[339] & b[303])^(a[338] & b[304])^(a[337] & b[305])^(a[336] & b[306])^(a[335] & b[307])^(a[334] & b[308])^(a[333] & b[309])^(a[332] & b[310])^(a[331] & b[311])^(a[330] & b[312])^(a[329] & b[313])^(a[328] & b[314])^(a[327] & b[315])^(a[326] & b[316])^(a[325] & b[317])^(a[324] & b[318])^(a[323] & b[319])^(a[322] & b[320])^(a[321] & b[321])^(a[320] & b[322])^(a[319] & b[323])^(a[318] & b[324])^(a[317] & b[325])^(a[316] & b[326])^(a[315] & b[327])^(a[314] & b[328])^(a[313] & b[329])^(a[312] & b[330])^(a[311] & b[331])^(a[310] & b[332])^(a[309] & b[333])^(a[308] & b[334])^(a[307] & b[335])^(a[306] & b[336])^(a[305] & b[337])^(a[304] & b[338])^(a[303] & b[339])^(a[302] & b[340])^(a[301] & b[341])^(a[300] & b[342])^(a[299] & b[343])^(a[298] & b[344])^(a[297] & b[345])^(a[296] & b[346])^(a[295] & b[347])^(a[294] & b[348])^(a[293] & b[349])^(a[292] & b[350])^(a[291] & b[351])^(a[290] & b[352])^(a[289] & b[353])^(a[288] & b[354])^(a[287] & b[355])^(a[286] & b[356])^(a[285] & b[357])^(a[284] & b[358])^(a[283] & b[359])^(a[282] & b[360])^(a[281] & b[361])^(a[280] & b[362])^(a[279] & b[363])^(a[278] & b[364])^(a[277] & b[365])^(a[276] & b[366])^(a[275] & b[367])^(a[274] & b[368])^(a[273] & b[369])^(a[272] & b[370])^(a[271] & b[371])^(a[270] & b[372])^(a[269] & b[373])^(a[268] & b[374])^(a[267] & b[375])^(a[266] & b[376])^(a[265] & b[377])^(a[264] & b[378])^(a[263] & b[379])^(a[262] & b[380])^(a[261] & b[381])^(a[260] & b[382])^(a[259] & b[383])^(a[258] & b[384])^(a[257] & b[385])^(a[256] & b[386])^(a[255] & b[387])^(a[254] & b[388])^(a[253] & b[389])^(a[252] & b[390])^(a[251] & b[391])^(a[250] & b[392])^(a[249] & b[393])^(a[248] & b[394])^(a[247] & b[395])^(a[246] & b[396])^(a[245] & b[397])^(a[244] & b[398])^(a[243] & b[399])^(a[242] & b[400])^(a[241] & b[401])^(a[240] & b[402])^(a[239] & b[403])^(a[238] & b[404])^(a[237] & b[405])^(a[236] & b[406])^(a[235] & b[407])^(a[234] & b[408]);
assign y[643] = (a[408] & b[235])^(a[407] & b[236])^(a[406] & b[237])^(a[405] & b[238])^(a[404] & b[239])^(a[403] & b[240])^(a[402] & b[241])^(a[401] & b[242])^(a[400] & b[243])^(a[399] & b[244])^(a[398] & b[245])^(a[397] & b[246])^(a[396] & b[247])^(a[395] & b[248])^(a[394] & b[249])^(a[393] & b[250])^(a[392] & b[251])^(a[391] & b[252])^(a[390] & b[253])^(a[389] & b[254])^(a[388] & b[255])^(a[387] & b[256])^(a[386] & b[257])^(a[385] & b[258])^(a[384] & b[259])^(a[383] & b[260])^(a[382] & b[261])^(a[381] & b[262])^(a[380] & b[263])^(a[379] & b[264])^(a[378] & b[265])^(a[377] & b[266])^(a[376] & b[267])^(a[375] & b[268])^(a[374] & b[269])^(a[373] & b[270])^(a[372] & b[271])^(a[371] & b[272])^(a[370] & b[273])^(a[369] & b[274])^(a[368] & b[275])^(a[367] & b[276])^(a[366] & b[277])^(a[365] & b[278])^(a[364] & b[279])^(a[363] & b[280])^(a[362] & b[281])^(a[361] & b[282])^(a[360] & b[283])^(a[359] & b[284])^(a[358] & b[285])^(a[357] & b[286])^(a[356] & b[287])^(a[355] & b[288])^(a[354] & b[289])^(a[353] & b[290])^(a[352] & b[291])^(a[351] & b[292])^(a[350] & b[293])^(a[349] & b[294])^(a[348] & b[295])^(a[347] & b[296])^(a[346] & b[297])^(a[345] & b[298])^(a[344] & b[299])^(a[343] & b[300])^(a[342] & b[301])^(a[341] & b[302])^(a[340] & b[303])^(a[339] & b[304])^(a[338] & b[305])^(a[337] & b[306])^(a[336] & b[307])^(a[335] & b[308])^(a[334] & b[309])^(a[333] & b[310])^(a[332] & b[311])^(a[331] & b[312])^(a[330] & b[313])^(a[329] & b[314])^(a[328] & b[315])^(a[327] & b[316])^(a[326] & b[317])^(a[325] & b[318])^(a[324] & b[319])^(a[323] & b[320])^(a[322] & b[321])^(a[321] & b[322])^(a[320] & b[323])^(a[319] & b[324])^(a[318] & b[325])^(a[317] & b[326])^(a[316] & b[327])^(a[315] & b[328])^(a[314] & b[329])^(a[313] & b[330])^(a[312] & b[331])^(a[311] & b[332])^(a[310] & b[333])^(a[309] & b[334])^(a[308] & b[335])^(a[307] & b[336])^(a[306] & b[337])^(a[305] & b[338])^(a[304] & b[339])^(a[303] & b[340])^(a[302] & b[341])^(a[301] & b[342])^(a[300] & b[343])^(a[299] & b[344])^(a[298] & b[345])^(a[297] & b[346])^(a[296] & b[347])^(a[295] & b[348])^(a[294] & b[349])^(a[293] & b[350])^(a[292] & b[351])^(a[291] & b[352])^(a[290] & b[353])^(a[289] & b[354])^(a[288] & b[355])^(a[287] & b[356])^(a[286] & b[357])^(a[285] & b[358])^(a[284] & b[359])^(a[283] & b[360])^(a[282] & b[361])^(a[281] & b[362])^(a[280] & b[363])^(a[279] & b[364])^(a[278] & b[365])^(a[277] & b[366])^(a[276] & b[367])^(a[275] & b[368])^(a[274] & b[369])^(a[273] & b[370])^(a[272] & b[371])^(a[271] & b[372])^(a[270] & b[373])^(a[269] & b[374])^(a[268] & b[375])^(a[267] & b[376])^(a[266] & b[377])^(a[265] & b[378])^(a[264] & b[379])^(a[263] & b[380])^(a[262] & b[381])^(a[261] & b[382])^(a[260] & b[383])^(a[259] & b[384])^(a[258] & b[385])^(a[257] & b[386])^(a[256] & b[387])^(a[255] & b[388])^(a[254] & b[389])^(a[253] & b[390])^(a[252] & b[391])^(a[251] & b[392])^(a[250] & b[393])^(a[249] & b[394])^(a[248] & b[395])^(a[247] & b[396])^(a[246] & b[397])^(a[245] & b[398])^(a[244] & b[399])^(a[243] & b[400])^(a[242] & b[401])^(a[241] & b[402])^(a[240] & b[403])^(a[239] & b[404])^(a[238] & b[405])^(a[237] & b[406])^(a[236] & b[407])^(a[235] & b[408]);
assign y[644] = (a[408] & b[236])^(a[407] & b[237])^(a[406] & b[238])^(a[405] & b[239])^(a[404] & b[240])^(a[403] & b[241])^(a[402] & b[242])^(a[401] & b[243])^(a[400] & b[244])^(a[399] & b[245])^(a[398] & b[246])^(a[397] & b[247])^(a[396] & b[248])^(a[395] & b[249])^(a[394] & b[250])^(a[393] & b[251])^(a[392] & b[252])^(a[391] & b[253])^(a[390] & b[254])^(a[389] & b[255])^(a[388] & b[256])^(a[387] & b[257])^(a[386] & b[258])^(a[385] & b[259])^(a[384] & b[260])^(a[383] & b[261])^(a[382] & b[262])^(a[381] & b[263])^(a[380] & b[264])^(a[379] & b[265])^(a[378] & b[266])^(a[377] & b[267])^(a[376] & b[268])^(a[375] & b[269])^(a[374] & b[270])^(a[373] & b[271])^(a[372] & b[272])^(a[371] & b[273])^(a[370] & b[274])^(a[369] & b[275])^(a[368] & b[276])^(a[367] & b[277])^(a[366] & b[278])^(a[365] & b[279])^(a[364] & b[280])^(a[363] & b[281])^(a[362] & b[282])^(a[361] & b[283])^(a[360] & b[284])^(a[359] & b[285])^(a[358] & b[286])^(a[357] & b[287])^(a[356] & b[288])^(a[355] & b[289])^(a[354] & b[290])^(a[353] & b[291])^(a[352] & b[292])^(a[351] & b[293])^(a[350] & b[294])^(a[349] & b[295])^(a[348] & b[296])^(a[347] & b[297])^(a[346] & b[298])^(a[345] & b[299])^(a[344] & b[300])^(a[343] & b[301])^(a[342] & b[302])^(a[341] & b[303])^(a[340] & b[304])^(a[339] & b[305])^(a[338] & b[306])^(a[337] & b[307])^(a[336] & b[308])^(a[335] & b[309])^(a[334] & b[310])^(a[333] & b[311])^(a[332] & b[312])^(a[331] & b[313])^(a[330] & b[314])^(a[329] & b[315])^(a[328] & b[316])^(a[327] & b[317])^(a[326] & b[318])^(a[325] & b[319])^(a[324] & b[320])^(a[323] & b[321])^(a[322] & b[322])^(a[321] & b[323])^(a[320] & b[324])^(a[319] & b[325])^(a[318] & b[326])^(a[317] & b[327])^(a[316] & b[328])^(a[315] & b[329])^(a[314] & b[330])^(a[313] & b[331])^(a[312] & b[332])^(a[311] & b[333])^(a[310] & b[334])^(a[309] & b[335])^(a[308] & b[336])^(a[307] & b[337])^(a[306] & b[338])^(a[305] & b[339])^(a[304] & b[340])^(a[303] & b[341])^(a[302] & b[342])^(a[301] & b[343])^(a[300] & b[344])^(a[299] & b[345])^(a[298] & b[346])^(a[297] & b[347])^(a[296] & b[348])^(a[295] & b[349])^(a[294] & b[350])^(a[293] & b[351])^(a[292] & b[352])^(a[291] & b[353])^(a[290] & b[354])^(a[289] & b[355])^(a[288] & b[356])^(a[287] & b[357])^(a[286] & b[358])^(a[285] & b[359])^(a[284] & b[360])^(a[283] & b[361])^(a[282] & b[362])^(a[281] & b[363])^(a[280] & b[364])^(a[279] & b[365])^(a[278] & b[366])^(a[277] & b[367])^(a[276] & b[368])^(a[275] & b[369])^(a[274] & b[370])^(a[273] & b[371])^(a[272] & b[372])^(a[271] & b[373])^(a[270] & b[374])^(a[269] & b[375])^(a[268] & b[376])^(a[267] & b[377])^(a[266] & b[378])^(a[265] & b[379])^(a[264] & b[380])^(a[263] & b[381])^(a[262] & b[382])^(a[261] & b[383])^(a[260] & b[384])^(a[259] & b[385])^(a[258] & b[386])^(a[257] & b[387])^(a[256] & b[388])^(a[255] & b[389])^(a[254] & b[390])^(a[253] & b[391])^(a[252] & b[392])^(a[251] & b[393])^(a[250] & b[394])^(a[249] & b[395])^(a[248] & b[396])^(a[247] & b[397])^(a[246] & b[398])^(a[245] & b[399])^(a[244] & b[400])^(a[243] & b[401])^(a[242] & b[402])^(a[241] & b[403])^(a[240] & b[404])^(a[239] & b[405])^(a[238] & b[406])^(a[237] & b[407])^(a[236] & b[408]);
assign y[645] = (a[408] & b[237])^(a[407] & b[238])^(a[406] & b[239])^(a[405] & b[240])^(a[404] & b[241])^(a[403] & b[242])^(a[402] & b[243])^(a[401] & b[244])^(a[400] & b[245])^(a[399] & b[246])^(a[398] & b[247])^(a[397] & b[248])^(a[396] & b[249])^(a[395] & b[250])^(a[394] & b[251])^(a[393] & b[252])^(a[392] & b[253])^(a[391] & b[254])^(a[390] & b[255])^(a[389] & b[256])^(a[388] & b[257])^(a[387] & b[258])^(a[386] & b[259])^(a[385] & b[260])^(a[384] & b[261])^(a[383] & b[262])^(a[382] & b[263])^(a[381] & b[264])^(a[380] & b[265])^(a[379] & b[266])^(a[378] & b[267])^(a[377] & b[268])^(a[376] & b[269])^(a[375] & b[270])^(a[374] & b[271])^(a[373] & b[272])^(a[372] & b[273])^(a[371] & b[274])^(a[370] & b[275])^(a[369] & b[276])^(a[368] & b[277])^(a[367] & b[278])^(a[366] & b[279])^(a[365] & b[280])^(a[364] & b[281])^(a[363] & b[282])^(a[362] & b[283])^(a[361] & b[284])^(a[360] & b[285])^(a[359] & b[286])^(a[358] & b[287])^(a[357] & b[288])^(a[356] & b[289])^(a[355] & b[290])^(a[354] & b[291])^(a[353] & b[292])^(a[352] & b[293])^(a[351] & b[294])^(a[350] & b[295])^(a[349] & b[296])^(a[348] & b[297])^(a[347] & b[298])^(a[346] & b[299])^(a[345] & b[300])^(a[344] & b[301])^(a[343] & b[302])^(a[342] & b[303])^(a[341] & b[304])^(a[340] & b[305])^(a[339] & b[306])^(a[338] & b[307])^(a[337] & b[308])^(a[336] & b[309])^(a[335] & b[310])^(a[334] & b[311])^(a[333] & b[312])^(a[332] & b[313])^(a[331] & b[314])^(a[330] & b[315])^(a[329] & b[316])^(a[328] & b[317])^(a[327] & b[318])^(a[326] & b[319])^(a[325] & b[320])^(a[324] & b[321])^(a[323] & b[322])^(a[322] & b[323])^(a[321] & b[324])^(a[320] & b[325])^(a[319] & b[326])^(a[318] & b[327])^(a[317] & b[328])^(a[316] & b[329])^(a[315] & b[330])^(a[314] & b[331])^(a[313] & b[332])^(a[312] & b[333])^(a[311] & b[334])^(a[310] & b[335])^(a[309] & b[336])^(a[308] & b[337])^(a[307] & b[338])^(a[306] & b[339])^(a[305] & b[340])^(a[304] & b[341])^(a[303] & b[342])^(a[302] & b[343])^(a[301] & b[344])^(a[300] & b[345])^(a[299] & b[346])^(a[298] & b[347])^(a[297] & b[348])^(a[296] & b[349])^(a[295] & b[350])^(a[294] & b[351])^(a[293] & b[352])^(a[292] & b[353])^(a[291] & b[354])^(a[290] & b[355])^(a[289] & b[356])^(a[288] & b[357])^(a[287] & b[358])^(a[286] & b[359])^(a[285] & b[360])^(a[284] & b[361])^(a[283] & b[362])^(a[282] & b[363])^(a[281] & b[364])^(a[280] & b[365])^(a[279] & b[366])^(a[278] & b[367])^(a[277] & b[368])^(a[276] & b[369])^(a[275] & b[370])^(a[274] & b[371])^(a[273] & b[372])^(a[272] & b[373])^(a[271] & b[374])^(a[270] & b[375])^(a[269] & b[376])^(a[268] & b[377])^(a[267] & b[378])^(a[266] & b[379])^(a[265] & b[380])^(a[264] & b[381])^(a[263] & b[382])^(a[262] & b[383])^(a[261] & b[384])^(a[260] & b[385])^(a[259] & b[386])^(a[258] & b[387])^(a[257] & b[388])^(a[256] & b[389])^(a[255] & b[390])^(a[254] & b[391])^(a[253] & b[392])^(a[252] & b[393])^(a[251] & b[394])^(a[250] & b[395])^(a[249] & b[396])^(a[248] & b[397])^(a[247] & b[398])^(a[246] & b[399])^(a[245] & b[400])^(a[244] & b[401])^(a[243] & b[402])^(a[242] & b[403])^(a[241] & b[404])^(a[240] & b[405])^(a[239] & b[406])^(a[238] & b[407])^(a[237] & b[408]);
assign y[646] = (a[408] & b[238])^(a[407] & b[239])^(a[406] & b[240])^(a[405] & b[241])^(a[404] & b[242])^(a[403] & b[243])^(a[402] & b[244])^(a[401] & b[245])^(a[400] & b[246])^(a[399] & b[247])^(a[398] & b[248])^(a[397] & b[249])^(a[396] & b[250])^(a[395] & b[251])^(a[394] & b[252])^(a[393] & b[253])^(a[392] & b[254])^(a[391] & b[255])^(a[390] & b[256])^(a[389] & b[257])^(a[388] & b[258])^(a[387] & b[259])^(a[386] & b[260])^(a[385] & b[261])^(a[384] & b[262])^(a[383] & b[263])^(a[382] & b[264])^(a[381] & b[265])^(a[380] & b[266])^(a[379] & b[267])^(a[378] & b[268])^(a[377] & b[269])^(a[376] & b[270])^(a[375] & b[271])^(a[374] & b[272])^(a[373] & b[273])^(a[372] & b[274])^(a[371] & b[275])^(a[370] & b[276])^(a[369] & b[277])^(a[368] & b[278])^(a[367] & b[279])^(a[366] & b[280])^(a[365] & b[281])^(a[364] & b[282])^(a[363] & b[283])^(a[362] & b[284])^(a[361] & b[285])^(a[360] & b[286])^(a[359] & b[287])^(a[358] & b[288])^(a[357] & b[289])^(a[356] & b[290])^(a[355] & b[291])^(a[354] & b[292])^(a[353] & b[293])^(a[352] & b[294])^(a[351] & b[295])^(a[350] & b[296])^(a[349] & b[297])^(a[348] & b[298])^(a[347] & b[299])^(a[346] & b[300])^(a[345] & b[301])^(a[344] & b[302])^(a[343] & b[303])^(a[342] & b[304])^(a[341] & b[305])^(a[340] & b[306])^(a[339] & b[307])^(a[338] & b[308])^(a[337] & b[309])^(a[336] & b[310])^(a[335] & b[311])^(a[334] & b[312])^(a[333] & b[313])^(a[332] & b[314])^(a[331] & b[315])^(a[330] & b[316])^(a[329] & b[317])^(a[328] & b[318])^(a[327] & b[319])^(a[326] & b[320])^(a[325] & b[321])^(a[324] & b[322])^(a[323] & b[323])^(a[322] & b[324])^(a[321] & b[325])^(a[320] & b[326])^(a[319] & b[327])^(a[318] & b[328])^(a[317] & b[329])^(a[316] & b[330])^(a[315] & b[331])^(a[314] & b[332])^(a[313] & b[333])^(a[312] & b[334])^(a[311] & b[335])^(a[310] & b[336])^(a[309] & b[337])^(a[308] & b[338])^(a[307] & b[339])^(a[306] & b[340])^(a[305] & b[341])^(a[304] & b[342])^(a[303] & b[343])^(a[302] & b[344])^(a[301] & b[345])^(a[300] & b[346])^(a[299] & b[347])^(a[298] & b[348])^(a[297] & b[349])^(a[296] & b[350])^(a[295] & b[351])^(a[294] & b[352])^(a[293] & b[353])^(a[292] & b[354])^(a[291] & b[355])^(a[290] & b[356])^(a[289] & b[357])^(a[288] & b[358])^(a[287] & b[359])^(a[286] & b[360])^(a[285] & b[361])^(a[284] & b[362])^(a[283] & b[363])^(a[282] & b[364])^(a[281] & b[365])^(a[280] & b[366])^(a[279] & b[367])^(a[278] & b[368])^(a[277] & b[369])^(a[276] & b[370])^(a[275] & b[371])^(a[274] & b[372])^(a[273] & b[373])^(a[272] & b[374])^(a[271] & b[375])^(a[270] & b[376])^(a[269] & b[377])^(a[268] & b[378])^(a[267] & b[379])^(a[266] & b[380])^(a[265] & b[381])^(a[264] & b[382])^(a[263] & b[383])^(a[262] & b[384])^(a[261] & b[385])^(a[260] & b[386])^(a[259] & b[387])^(a[258] & b[388])^(a[257] & b[389])^(a[256] & b[390])^(a[255] & b[391])^(a[254] & b[392])^(a[253] & b[393])^(a[252] & b[394])^(a[251] & b[395])^(a[250] & b[396])^(a[249] & b[397])^(a[248] & b[398])^(a[247] & b[399])^(a[246] & b[400])^(a[245] & b[401])^(a[244] & b[402])^(a[243] & b[403])^(a[242] & b[404])^(a[241] & b[405])^(a[240] & b[406])^(a[239] & b[407])^(a[238] & b[408]);
assign y[647] = (a[408] & b[239])^(a[407] & b[240])^(a[406] & b[241])^(a[405] & b[242])^(a[404] & b[243])^(a[403] & b[244])^(a[402] & b[245])^(a[401] & b[246])^(a[400] & b[247])^(a[399] & b[248])^(a[398] & b[249])^(a[397] & b[250])^(a[396] & b[251])^(a[395] & b[252])^(a[394] & b[253])^(a[393] & b[254])^(a[392] & b[255])^(a[391] & b[256])^(a[390] & b[257])^(a[389] & b[258])^(a[388] & b[259])^(a[387] & b[260])^(a[386] & b[261])^(a[385] & b[262])^(a[384] & b[263])^(a[383] & b[264])^(a[382] & b[265])^(a[381] & b[266])^(a[380] & b[267])^(a[379] & b[268])^(a[378] & b[269])^(a[377] & b[270])^(a[376] & b[271])^(a[375] & b[272])^(a[374] & b[273])^(a[373] & b[274])^(a[372] & b[275])^(a[371] & b[276])^(a[370] & b[277])^(a[369] & b[278])^(a[368] & b[279])^(a[367] & b[280])^(a[366] & b[281])^(a[365] & b[282])^(a[364] & b[283])^(a[363] & b[284])^(a[362] & b[285])^(a[361] & b[286])^(a[360] & b[287])^(a[359] & b[288])^(a[358] & b[289])^(a[357] & b[290])^(a[356] & b[291])^(a[355] & b[292])^(a[354] & b[293])^(a[353] & b[294])^(a[352] & b[295])^(a[351] & b[296])^(a[350] & b[297])^(a[349] & b[298])^(a[348] & b[299])^(a[347] & b[300])^(a[346] & b[301])^(a[345] & b[302])^(a[344] & b[303])^(a[343] & b[304])^(a[342] & b[305])^(a[341] & b[306])^(a[340] & b[307])^(a[339] & b[308])^(a[338] & b[309])^(a[337] & b[310])^(a[336] & b[311])^(a[335] & b[312])^(a[334] & b[313])^(a[333] & b[314])^(a[332] & b[315])^(a[331] & b[316])^(a[330] & b[317])^(a[329] & b[318])^(a[328] & b[319])^(a[327] & b[320])^(a[326] & b[321])^(a[325] & b[322])^(a[324] & b[323])^(a[323] & b[324])^(a[322] & b[325])^(a[321] & b[326])^(a[320] & b[327])^(a[319] & b[328])^(a[318] & b[329])^(a[317] & b[330])^(a[316] & b[331])^(a[315] & b[332])^(a[314] & b[333])^(a[313] & b[334])^(a[312] & b[335])^(a[311] & b[336])^(a[310] & b[337])^(a[309] & b[338])^(a[308] & b[339])^(a[307] & b[340])^(a[306] & b[341])^(a[305] & b[342])^(a[304] & b[343])^(a[303] & b[344])^(a[302] & b[345])^(a[301] & b[346])^(a[300] & b[347])^(a[299] & b[348])^(a[298] & b[349])^(a[297] & b[350])^(a[296] & b[351])^(a[295] & b[352])^(a[294] & b[353])^(a[293] & b[354])^(a[292] & b[355])^(a[291] & b[356])^(a[290] & b[357])^(a[289] & b[358])^(a[288] & b[359])^(a[287] & b[360])^(a[286] & b[361])^(a[285] & b[362])^(a[284] & b[363])^(a[283] & b[364])^(a[282] & b[365])^(a[281] & b[366])^(a[280] & b[367])^(a[279] & b[368])^(a[278] & b[369])^(a[277] & b[370])^(a[276] & b[371])^(a[275] & b[372])^(a[274] & b[373])^(a[273] & b[374])^(a[272] & b[375])^(a[271] & b[376])^(a[270] & b[377])^(a[269] & b[378])^(a[268] & b[379])^(a[267] & b[380])^(a[266] & b[381])^(a[265] & b[382])^(a[264] & b[383])^(a[263] & b[384])^(a[262] & b[385])^(a[261] & b[386])^(a[260] & b[387])^(a[259] & b[388])^(a[258] & b[389])^(a[257] & b[390])^(a[256] & b[391])^(a[255] & b[392])^(a[254] & b[393])^(a[253] & b[394])^(a[252] & b[395])^(a[251] & b[396])^(a[250] & b[397])^(a[249] & b[398])^(a[248] & b[399])^(a[247] & b[400])^(a[246] & b[401])^(a[245] & b[402])^(a[244] & b[403])^(a[243] & b[404])^(a[242] & b[405])^(a[241] & b[406])^(a[240] & b[407])^(a[239] & b[408]);
assign y[648] = (a[408] & b[240])^(a[407] & b[241])^(a[406] & b[242])^(a[405] & b[243])^(a[404] & b[244])^(a[403] & b[245])^(a[402] & b[246])^(a[401] & b[247])^(a[400] & b[248])^(a[399] & b[249])^(a[398] & b[250])^(a[397] & b[251])^(a[396] & b[252])^(a[395] & b[253])^(a[394] & b[254])^(a[393] & b[255])^(a[392] & b[256])^(a[391] & b[257])^(a[390] & b[258])^(a[389] & b[259])^(a[388] & b[260])^(a[387] & b[261])^(a[386] & b[262])^(a[385] & b[263])^(a[384] & b[264])^(a[383] & b[265])^(a[382] & b[266])^(a[381] & b[267])^(a[380] & b[268])^(a[379] & b[269])^(a[378] & b[270])^(a[377] & b[271])^(a[376] & b[272])^(a[375] & b[273])^(a[374] & b[274])^(a[373] & b[275])^(a[372] & b[276])^(a[371] & b[277])^(a[370] & b[278])^(a[369] & b[279])^(a[368] & b[280])^(a[367] & b[281])^(a[366] & b[282])^(a[365] & b[283])^(a[364] & b[284])^(a[363] & b[285])^(a[362] & b[286])^(a[361] & b[287])^(a[360] & b[288])^(a[359] & b[289])^(a[358] & b[290])^(a[357] & b[291])^(a[356] & b[292])^(a[355] & b[293])^(a[354] & b[294])^(a[353] & b[295])^(a[352] & b[296])^(a[351] & b[297])^(a[350] & b[298])^(a[349] & b[299])^(a[348] & b[300])^(a[347] & b[301])^(a[346] & b[302])^(a[345] & b[303])^(a[344] & b[304])^(a[343] & b[305])^(a[342] & b[306])^(a[341] & b[307])^(a[340] & b[308])^(a[339] & b[309])^(a[338] & b[310])^(a[337] & b[311])^(a[336] & b[312])^(a[335] & b[313])^(a[334] & b[314])^(a[333] & b[315])^(a[332] & b[316])^(a[331] & b[317])^(a[330] & b[318])^(a[329] & b[319])^(a[328] & b[320])^(a[327] & b[321])^(a[326] & b[322])^(a[325] & b[323])^(a[324] & b[324])^(a[323] & b[325])^(a[322] & b[326])^(a[321] & b[327])^(a[320] & b[328])^(a[319] & b[329])^(a[318] & b[330])^(a[317] & b[331])^(a[316] & b[332])^(a[315] & b[333])^(a[314] & b[334])^(a[313] & b[335])^(a[312] & b[336])^(a[311] & b[337])^(a[310] & b[338])^(a[309] & b[339])^(a[308] & b[340])^(a[307] & b[341])^(a[306] & b[342])^(a[305] & b[343])^(a[304] & b[344])^(a[303] & b[345])^(a[302] & b[346])^(a[301] & b[347])^(a[300] & b[348])^(a[299] & b[349])^(a[298] & b[350])^(a[297] & b[351])^(a[296] & b[352])^(a[295] & b[353])^(a[294] & b[354])^(a[293] & b[355])^(a[292] & b[356])^(a[291] & b[357])^(a[290] & b[358])^(a[289] & b[359])^(a[288] & b[360])^(a[287] & b[361])^(a[286] & b[362])^(a[285] & b[363])^(a[284] & b[364])^(a[283] & b[365])^(a[282] & b[366])^(a[281] & b[367])^(a[280] & b[368])^(a[279] & b[369])^(a[278] & b[370])^(a[277] & b[371])^(a[276] & b[372])^(a[275] & b[373])^(a[274] & b[374])^(a[273] & b[375])^(a[272] & b[376])^(a[271] & b[377])^(a[270] & b[378])^(a[269] & b[379])^(a[268] & b[380])^(a[267] & b[381])^(a[266] & b[382])^(a[265] & b[383])^(a[264] & b[384])^(a[263] & b[385])^(a[262] & b[386])^(a[261] & b[387])^(a[260] & b[388])^(a[259] & b[389])^(a[258] & b[390])^(a[257] & b[391])^(a[256] & b[392])^(a[255] & b[393])^(a[254] & b[394])^(a[253] & b[395])^(a[252] & b[396])^(a[251] & b[397])^(a[250] & b[398])^(a[249] & b[399])^(a[248] & b[400])^(a[247] & b[401])^(a[246] & b[402])^(a[245] & b[403])^(a[244] & b[404])^(a[243] & b[405])^(a[242] & b[406])^(a[241] & b[407])^(a[240] & b[408]);
assign y[649] = (a[408] & b[241])^(a[407] & b[242])^(a[406] & b[243])^(a[405] & b[244])^(a[404] & b[245])^(a[403] & b[246])^(a[402] & b[247])^(a[401] & b[248])^(a[400] & b[249])^(a[399] & b[250])^(a[398] & b[251])^(a[397] & b[252])^(a[396] & b[253])^(a[395] & b[254])^(a[394] & b[255])^(a[393] & b[256])^(a[392] & b[257])^(a[391] & b[258])^(a[390] & b[259])^(a[389] & b[260])^(a[388] & b[261])^(a[387] & b[262])^(a[386] & b[263])^(a[385] & b[264])^(a[384] & b[265])^(a[383] & b[266])^(a[382] & b[267])^(a[381] & b[268])^(a[380] & b[269])^(a[379] & b[270])^(a[378] & b[271])^(a[377] & b[272])^(a[376] & b[273])^(a[375] & b[274])^(a[374] & b[275])^(a[373] & b[276])^(a[372] & b[277])^(a[371] & b[278])^(a[370] & b[279])^(a[369] & b[280])^(a[368] & b[281])^(a[367] & b[282])^(a[366] & b[283])^(a[365] & b[284])^(a[364] & b[285])^(a[363] & b[286])^(a[362] & b[287])^(a[361] & b[288])^(a[360] & b[289])^(a[359] & b[290])^(a[358] & b[291])^(a[357] & b[292])^(a[356] & b[293])^(a[355] & b[294])^(a[354] & b[295])^(a[353] & b[296])^(a[352] & b[297])^(a[351] & b[298])^(a[350] & b[299])^(a[349] & b[300])^(a[348] & b[301])^(a[347] & b[302])^(a[346] & b[303])^(a[345] & b[304])^(a[344] & b[305])^(a[343] & b[306])^(a[342] & b[307])^(a[341] & b[308])^(a[340] & b[309])^(a[339] & b[310])^(a[338] & b[311])^(a[337] & b[312])^(a[336] & b[313])^(a[335] & b[314])^(a[334] & b[315])^(a[333] & b[316])^(a[332] & b[317])^(a[331] & b[318])^(a[330] & b[319])^(a[329] & b[320])^(a[328] & b[321])^(a[327] & b[322])^(a[326] & b[323])^(a[325] & b[324])^(a[324] & b[325])^(a[323] & b[326])^(a[322] & b[327])^(a[321] & b[328])^(a[320] & b[329])^(a[319] & b[330])^(a[318] & b[331])^(a[317] & b[332])^(a[316] & b[333])^(a[315] & b[334])^(a[314] & b[335])^(a[313] & b[336])^(a[312] & b[337])^(a[311] & b[338])^(a[310] & b[339])^(a[309] & b[340])^(a[308] & b[341])^(a[307] & b[342])^(a[306] & b[343])^(a[305] & b[344])^(a[304] & b[345])^(a[303] & b[346])^(a[302] & b[347])^(a[301] & b[348])^(a[300] & b[349])^(a[299] & b[350])^(a[298] & b[351])^(a[297] & b[352])^(a[296] & b[353])^(a[295] & b[354])^(a[294] & b[355])^(a[293] & b[356])^(a[292] & b[357])^(a[291] & b[358])^(a[290] & b[359])^(a[289] & b[360])^(a[288] & b[361])^(a[287] & b[362])^(a[286] & b[363])^(a[285] & b[364])^(a[284] & b[365])^(a[283] & b[366])^(a[282] & b[367])^(a[281] & b[368])^(a[280] & b[369])^(a[279] & b[370])^(a[278] & b[371])^(a[277] & b[372])^(a[276] & b[373])^(a[275] & b[374])^(a[274] & b[375])^(a[273] & b[376])^(a[272] & b[377])^(a[271] & b[378])^(a[270] & b[379])^(a[269] & b[380])^(a[268] & b[381])^(a[267] & b[382])^(a[266] & b[383])^(a[265] & b[384])^(a[264] & b[385])^(a[263] & b[386])^(a[262] & b[387])^(a[261] & b[388])^(a[260] & b[389])^(a[259] & b[390])^(a[258] & b[391])^(a[257] & b[392])^(a[256] & b[393])^(a[255] & b[394])^(a[254] & b[395])^(a[253] & b[396])^(a[252] & b[397])^(a[251] & b[398])^(a[250] & b[399])^(a[249] & b[400])^(a[248] & b[401])^(a[247] & b[402])^(a[246] & b[403])^(a[245] & b[404])^(a[244] & b[405])^(a[243] & b[406])^(a[242] & b[407])^(a[241] & b[408]);
assign y[650] = (a[408] & b[242])^(a[407] & b[243])^(a[406] & b[244])^(a[405] & b[245])^(a[404] & b[246])^(a[403] & b[247])^(a[402] & b[248])^(a[401] & b[249])^(a[400] & b[250])^(a[399] & b[251])^(a[398] & b[252])^(a[397] & b[253])^(a[396] & b[254])^(a[395] & b[255])^(a[394] & b[256])^(a[393] & b[257])^(a[392] & b[258])^(a[391] & b[259])^(a[390] & b[260])^(a[389] & b[261])^(a[388] & b[262])^(a[387] & b[263])^(a[386] & b[264])^(a[385] & b[265])^(a[384] & b[266])^(a[383] & b[267])^(a[382] & b[268])^(a[381] & b[269])^(a[380] & b[270])^(a[379] & b[271])^(a[378] & b[272])^(a[377] & b[273])^(a[376] & b[274])^(a[375] & b[275])^(a[374] & b[276])^(a[373] & b[277])^(a[372] & b[278])^(a[371] & b[279])^(a[370] & b[280])^(a[369] & b[281])^(a[368] & b[282])^(a[367] & b[283])^(a[366] & b[284])^(a[365] & b[285])^(a[364] & b[286])^(a[363] & b[287])^(a[362] & b[288])^(a[361] & b[289])^(a[360] & b[290])^(a[359] & b[291])^(a[358] & b[292])^(a[357] & b[293])^(a[356] & b[294])^(a[355] & b[295])^(a[354] & b[296])^(a[353] & b[297])^(a[352] & b[298])^(a[351] & b[299])^(a[350] & b[300])^(a[349] & b[301])^(a[348] & b[302])^(a[347] & b[303])^(a[346] & b[304])^(a[345] & b[305])^(a[344] & b[306])^(a[343] & b[307])^(a[342] & b[308])^(a[341] & b[309])^(a[340] & b[310])^(a[339] & b[311])^(a[338] & b[312])^(a[337] & b[313])^(a[336] & b[314])^(a[335] & b[315])^(a[334] & b[316])^(a[333] & b[317])^(a[332] & b[318])^(a[331] & b[319])^(a[330] & b[320])^(a[329] & b[321])^(a[328] & b[322])^(a[327] & b[323])^(a[326] & b[324])^(a[325] & b[325])^(a[324] & b[326])^(a[323] & b[327])^(a[322] & b[328])^(a[321] & b[329])^(a[320] & b[330])^(a[319] & b[331])^(a[318] & b[332])^(a[317] & b[333])^(a[316] & b[334])^(a[315] & b[335])^(a[314] & b[336])^(a[313] & b[337])^(a[312] & b[338])^(a[311] & b[339])^(a[310] & b[340])^(a[309] & b[341])^(a[308] & b[342])^(a[307] & b[343])^(a[306] & b[344])^(a[305] & b[345])^(a[304] & b[346])^(a[303] & b[347])^(a[302] & b[348])^(a[301] & b[349])^(a[300] & b[350])^(a[299] & b[351])^(a[298] & b[352])^(a[297] & b[353])^(a[296] & b[354])^(a[295] & b[355])^(a[294] & b[356])^(a[293] & b[357])^(a[292] & b[358])^(a[291] & b[359])^(a[290] & b[360])^(a[289] & b[361])^(a[288] & b[362])^(a[287] & b[363])^(a[286] & b[364])^(a[285] & b[365])^(a[284] & b[366])^(a[283] & b[367])^(a[282] & b[368])^(a[281] & b[369])^(a[280] & b[370])^(a[279] & b[371])^(a[278] & b[372])^(a[277] & b[373])^(a[276] & b[374])^(a[275] & b[375])^(a[274] & b[376])^(a[273] & b[377])^(a[272] & b[378])^(a[271] & b[379])^(a[270] & b[380])^(a[269] & b[381])^(a[268] & b[382])^(a[267] & b[383])^(a[266] & b[384])^(a[265] & b[385])^(a[264] & b[386])^(a[263] & b[387])^(a[262] & b[388])^(a[261] & b[389])^(a[260] & b[390])^(a[259] & b[391])^(a[258] & b[392])^(a[257] & b[393])^(a[256] & b[394])^(a[255] & b[395])^(a[254] & b[396])^(a[253] & b[397])^(a[252] & b[398])^(a[251] & b[399])^(a[250] & b[400])^(a[249] & b[401])^(a[248] & b[402])^(a[247] & b[403])^(a[246] & b[404])^(a[245] & b[405])^(a[244] & b[406])^(a[243] & b[407])^(a[242] & b[408]);
assign y[651] = (a[408] & b[243])^(a[407] & b[244])^(a[406] & b[245])^(a[405] & b[246])^(a[404] & b[247])^(a[403] & b[248])^(a[402] & b[249])^(a[401] & b[250])^(a[400] & b[251])^(a[399] & b[252])^(a[398] & b[253])^(a[397] & b[254])^(a[396] & b[255])^(a[395] & b[256])^(a[394] & b[257])^(a[393] & b[258])^(a[392] & b[259])^(a[391] & b[260])^(a[390] & b[261])^(a[389] & b[262])^(a[388] & b[263])^(a[387] & b[264])^(a[386] & b[265])^(a[385] & b[266])^(a[384] & b[267])^(a[383] & b[268])^(a[382] & b[269])^(a[381] & b[270])^(a[380] & b[271])^(a[379] & b[272])^(a[378] & b[273])^(a[377] & b[274])^(a[376] & b[275])^(a[375] & b[276])^(a[374] & b[277])^(a[373] & b[278])^(a[372] & b[279])^(a[371] & b[280])^(a[370] & b[281])^(a[369] & b[282])^(a[368] & b[283])^(a[367] & b[284])^(a[366] & b[285])^(a[365] & b[286])^(a[364] & b[287])^(a[363] & b[288])^(a[362] & b[289])^(a[361] & b[290])^(a[360] & b[291])^(a[359] & b[292])^(a[358] & b[293])^(a[357] & b[294])^(a[356] & b[295])^(a[355] & b[296])^(a[354] & b[297])^(a[353] & b[298])^(a[352] & b[299])^(a[351] & b[300])^(a[350] & b[301])^(a[349] & b[302])^(a[348] & b[303])^(a[347] & b[304])^(a[346] & b[305])^(a[345] & b[306])^(a[344] & b[307])^(a[343] & b[308])^(a[342] & b[309])^(a[341] & b[310])^(a[340] & b[311])^(a[339] & b[312])^(a[338] & b[313])^(a[337] & b[314])^(a[336] & b[315])^(a[335] & b[316])^(a[334] & b[317])^(a[333] & b[318])^(a[332] & b[319])^(a[331] & b[320])^(a[330] & b[321])^(a[329] & b[322])^(a[328] & b[323])^(a[327] & b[324])^(a[326] & b[325])^(a[325] & b[326])^(a[324] & b[327])^(a[323] & b[328])^(a[322] & b[329])^(a[321] & b[330])^(a[320] & b[331])^(a[319] & b[332])^(a[318] & b[333])^(a[317] & b[334])^(a[316] & b[335])^(a[315] & b[336])^(a[314] & b[337])^(a[313] & b[338])^(a[312] & b[339])^(a[311] & b[340])^(a[310] & b[341])^(a[309] & b[342])^(a[308] & b[343])^(a[307] & b[344])^(a[306] & b[345])^(a[305] & b[346])^(a[304] & b[347])^(a[303] & b[348])^(a[302] & b[349])^(a[301] & b[350])^(a[300] & b[351])^(a[299] & b[352])^(a[298] & b[353])^(a[297] & b[354])^(a[296] & b[355])^(a[295] & b[356])^(a[294] & b[357])^(a[293] & b[358])^(a[292] & b[359])^(a[291] & b[360])^(a[290] & b[361])^(a[289] & b[362])^(a[288] & b[363])^(a[287] & b[364])^(a[286] & b[365])^(a[285] & b[366])^(a[284] & b[367])^(a[283] & b[368])^(a[282] & b[369])^(a[281] & b[370])^(a[280] & b[371])^(a[279] & b[372])^(a[278] & b[373])^(a[277] & b[374])^(a[276] & b[375])^(a[275] & b[376])^(a[274] & b[377])^(a[273] & b[378])^(a[272] & b[379])^(a[271] & b[380])^(a[270] & b[381])^(a[269] & b[382])^(a[268] & b[383])^(a[267] & b[384])^(a[266] & b[385])^(a[265] & b[386])^(a[264] & b[387])^(a[263] & b[388])^(a[262] & b[389])^(a[261] & b[390])^(a[260] & b[391])^(a[259] & b[392])^(a[258] & b[393])^(a[257] & b[394])^(a[256] & b[395])^(a[255] & b[396])^(a[254] & b[397])^(a[253] & b[398])^(a[252] & b[399])^(a[251] & b[400])^(a[250] & b[401])^(a[249] & b[402])^(a[248] & b[403])^(a[247] & b[404])^(a[246] & b[405])^(a[245] & b[406])^(a[244] & b[407])^(a[243] & b[408]);
assign y[652] = (a[408] & b[244])^(a[407] & b[245])^(a[406] & b[246])^(a[405] & b[247])^(a[404] & b[248])^(a[403] & b[249])^(a[402] & b[250])^(a[401] & b[251])^(a[400] & b[252])^(a[399] & b[253])^(a[398] & b[254])^(a[397] & b[255])^(a[396] & b[256])^(a[395] & b[257])^(a[394] & b[258])^(a[393] & b[259])^(a[392] & b[260])^(a[391] & b[261])^(a[390] & b[262])^(a[389] & b[263])^(a[388] & b[264])^(a[387] & b[265])^(a[386] & b[266])^(a[385] & b[267])^(a[384] & b[268])^(a[383] & b[269])^(a[382] & b[270])^(a[381] & b[271])^(a[380] & b[272])^(a[379] & b[273])^(a[378] & b[274])^(a[377] & b[275])^(a[376] & b[276])^(a[375] & b[277])^(a[374] & b[278])^(a[373] & b[279])^(a[372] & b[280])^(a[371] & b[281])^(a[370] & b[282])^(a[369] & b[283])^(a[368] & b[284])^(a[367] & b[285])^(a[366] & b[286])^(a[365] & b[287])^(a[364] & b[288])^(a[363] & b[289])^(a[362] & b[290])^(a[361] & b[291])^(a[360] & b[292])^(a[359] & b[293])^(a[358] & b[294])^(a[357] & b[295])^(a[356] & b[296])^(a[355] & b[297])^(a[354] & b[298])^(a[353] & b[299])^(a[352] & b[300])^(a[351] & b[301])^(a[350] & b[302])^(a[349] & b[303])^(a[348] & b[304])^(a[347] & b[305])^(a[346] & b[306])^(a[345] & b[307])^(a[344] & b[308])^(a[343] & b[309])^(a[342] & b[310])^(a[341] & b[311])^(a[340] & b[312])^(a[339] & b[313])^(a[338] & b[314])^(a[337] & b[315])^(a[336] & b[316])^(a[335] & b[317])^(a[334] & b[318])^(a[333] & b[319])^(a[332] & b[320])^(a[331] & b[321])^(a[330] & b[322])^(a[329] & b[323])^(a[328] & b[324])^(a[327] & b[325])^(a[326] & b[326])^(a[325] & b[327])^(a[324] & b[328])^(a[323] & b[329])^(a[322] & b[330])^(a[321] & b[331])^(a[320] & b[332])^(a[319] & b[333])^(a[318] & b[334])^(a[317] & b[335])^(a[316] & b[336])^(a[315] & b[337])^(a[314] & b[338])^(a[313] & b[339])^(a[312] & b[340])^(a[311] & b[341])^(a[310] & b[342])^(a[309] & b[343])^(a[308] & b[344])^(a[307] & b[345])^(a[306] & b[346])^(a[305] & b[347])^(a[304] & b[348])^(a[303] & b[349])^(a[302] & b[350])^(a[301] & b[351])^(a[300] & b[352])^(a[299] & b[353])^(a[298] & b[354])^(a[297] & b[355])^(a[296] & b[356])^(a[295] & b[357])^(a[294] & b[358])^(a[293] & b[359])^(a[292] & b[360])^(a[291] & b[361])^(a[290] & b[362])^(a[289] & b[363])^(a[288] & b[364])^(a[287] & b[365])^(a[286] & b[366])^(a[285] & b[367])^(a[284] & b[368])^(a[283] & b[369])^(a[282] & b[370])^(a[281] & b[371])^(a[280] & b[372])^(a[279] & b[373])^(a[278] & b[374])^(a[277] & b[375])^(a[276] & b[376])^(a[275] & b[377])^(a[274] & b[378])^(a[273] & b[379])^(a[272] & b[380])^(a[271] & b[381])^(a[270] & b[382])^(a[269] & b[383])^(a[268] & b[384])^(a[267] & b[385])^(a[266] & b[386])^(a[265] & b[387])^(a[264] & b[388])^(a[263] & b[389])^(a[262] & b[390])^(a[261] & b[391])^(a[260] & b[392])^(a[259] & b[393])^(a[258] & b[394])^(a[257] & b[395])^(a[256] & b[396])^(a[255] & b[397])^(a[254] & b[398])^(a[253] & b[399])^(a[252] & b[400])^(a[251] & b[401])^(a[250] & b[402])^(a[249] & b[403])^(a[248] & b[404])^(a[247] & b[405])^(a[246] & b[406])^(a[245] & b[407])^(a[244] & b[408]);
assign y[653] = (a[408] & b[245])^(a[407] & b[246])^(a[406] & b[247])^(a[405] & b[248])^(a[404] & b[249])^(a[403] & b[250])^(a[402] & b[251])^(a[401] & b[252])^(a[400] & b[253])^(a[399] & b[254])^(a[398] & b[255])^(a[397] & b[256])^(a[396] & b[257])^(a[395] & b[258])^(a[394] & b[259])^(a[393] & b[260])^(a[392] & b[261])^(a[391] & b[262])^(a[390] & b[263])^(a[389] & b[264])^(a[388] & b[265])^(a[387] & b[266])^(a[386] & b[267])^(a[385] & b[268])^(a[384] & b[269])^(a[383] & b[270])^(a[382] & b[271])^(a[381] & b[272])^(a[380] & b[273])^(a[379] & b[274])^(a[378] & b[275])^(a[377] & b[276])^(a[376] & b[277])^(a[375] & b[278])^(a[374] & b[279])^(a[373] & b[280])^(a[372] & b[281])^(a[371] & b[282])^(a[370] & b[283])^(a[369] & b[284])^(a[368] & b[285])^(a[367] & b[286])^(a[366] & b[287])^(a[365] & b[288])^(a[364] & b[289])^(a[363] & b[290])^(a[362] & b[291])^(a[361] & b[292])^(a[360] & b[293])^(a[359] & b[294])^(a[358] & b[295])^(a[357] & b[296])^(a[356] & b[297])^(a[355] & b[298])^(a[354] & b[299])^(a[353] & b[300])^(a[352] & b[301])^(a[351] & b[302])^(a[350] & b[303])^(a[349] & b[304])^(a[348] & b[305])^(a[347] & b[306])^(a[346] & b[307])^(a[345] & b[308])^(a[344] & b[309])^(a[343] & b[310])^(a[342] & b[311])^(a[341] & b[312])^(a[340] & b[313])^(a[339] & b[314])^(a[338] & b[315])^(a[337] & b[316])^(a[336] & b[317])^(a[335] & b[318])^(a[334] & b[319])^(a[333] & b[320])^(a[332] & b[321])^(a[331] & b[322])^(a[330] & b[323])^(a[329] & b[324])^(a[328] & b[325])^(a[327] & b[326])^(a[326] & b[327])^(a[325] & b[328])^(a[324] & b[329])^(a[323] & b[330])^(a[322] & b[331])^(a[321] & b[332])^(a[320] & b[333])^(a[319] & b[334])^(a[318] & b[335])^(a[317] & b[336])^(a[316] & b[337])^(a[315] & b[338])^(a[314] & b[339])^(a[313] & b[340])^(a[312] & b[341])^(a[311] & b[342])^(a[310] & b[343])^(a[309] & b[344])^(a[308] & b[345])^(a[307] & b[346])^(a[306] & b[347])^(a[305] & b[348])^(a[304] & b[349])^(a[303] & b[350])^(a[302] & b[351])^(a[301] & b[352])^(a[300] & b[353])^(a[299] & b[354])^(a[298] & b[355])^(a[297] & b[356])^(a[296] & b[357])^(a[295] & b[358])^(a[294] & b[359])^(a[293] & b[360])^(a[292] & b[361])^(a[291] & b[362])^(a[290] & b[363])^(a[289] & b[364])^(a[288] & b[365])^(a[287] & b[366])^(a[286] & b[367])^(a[285] & b[368])^(a[284] & b[369])^(a[283] & b[370])^(a[282] & b[371])^(a[281] & b[372])^(a[280] & b[373])^(a[279] & b[374])^(a[278] & b[375])^(a[277] & b[376])^(a[276] & b[377])^(a[275] & b[378])^(a[274] & b[379])^(a[273] & b[380])^(a[272] & b[381])^(a[271] & b[382])^(a[270] & b[383])^(a[269] & b[384])^(a[268] & b[385])^(a[267] & b[386])^(a[266] & b[387])^(a[265] & b[388])^(a[264] & b[389])^(a[263] & b[390])^(a[262] & b[391])^(a[261] & b[392])^(a[260] & b[393])^(a[259] & b[394])^(a[258] & b[395])^(a[257] & b[396])^(a[256] & b[397])^(a[255] & b[398])^(a[254] & b[399])^(a[253] & b[400])^(a[252] & b[401])^(a[251] & b[402])^(a[250] & b[403])^(a[249] & b[404])^(a[248] & b[405])^(a[247] & b[406])^(a[246] & b[407])^(a[245] & b[408]);
assign y[654] = (a[408] & b[246])^(a[407] & b[247])^(a[406] & b[248])^(a[405] & b[249])^(a[404] & b[250])^(a[403] & b[251])^(a[402] & b[252])^(a[401] & b[253])^(a[400] & b[254])^(a[399] & b[255])^(a[398] & b[256])^(a[397] & b[257])^(a[396] & b[258])^(a[395] & b[259])^(a[394] & b[260])^(a[393] & b[261])^(a[392] & b[262])^(a[391] & b[263])^(a[390] & b[264])^(a[389] & b[265])^(a[388] & b[266])^(a[387] & b[267])^(a[386] & b[268])^(a[385] & b[269])^(a[384] & b[270])^(a[383] & b[271])^(a[382] & b[272])^(a[381] & b[273])^(a[380] & b[274])^(a[379] & b[275])^(a[378] & b[276])^(a[377] & b[277])^(a[376] & b[278])^(a[375] & b[279])^(a[374] & b[280])^(a[373] & b[281])^(a[372] & b[282])^(a[371] & b[283])^(a[370] & b[284])^(a[369] & b[285])^(a[368] & b[286])^(a[367] & b[287])^(a[366] & b[288])^(a[365] & b[289])^(a[364] & b[290])^(a[363] & b[291])^(a[362] & b[292])^(a[361] & b[293])^(a[360] & b[294])^(a[359] & b[295])^(a[358] & b[296])^(a[357] & b[297])^(a[356] & b[298])^(a[355] & b[299])^(a[354] & b[300])^(a[353] & b[301])^(a[352] & b[302])^(a[351] & b[303])^(a[350] & b[304])^(a[349] & b[305])^(a[348] & b[306])^(a[347] & b[307])^(a[346] & b[308])^(a[345] & b[309])^(a[344] & b[310])^(a[343] & b[311])^(a[342] & b[312])^(a[341] & b[313])^(a[340] & b[314])^(a[339] & b[315])^(a[338] & b[316])^(a[337] & b[317])^(a[336] & b[318])^(a[335] & b[319])^(a[334] & b[320])^(a[333] & b[321])^(a[332] & b[322])^(a[331] & b[323])^(a[330] & b[324])^(a[329] & b[325])^(a[328] & b[326])^(a[327] & b[327])^(a[326] & b[328])^(a[325] & b[329])^(a[324] & b[330])^(a[323] & b[331])^(a[322] & b[332])^(a[321] & b[333])^(a[320] & b[334])^(a[319] & b[335])^(a[318] & b[336])^(a[317] & b[337])^(a[316] & b[338])^(a[315] & b[339])^(a[314] & b[340])^(a[313] & b[341])^(a[312] & b[342])^(a[311] & b[343])^(a[310] & b[344])^(a[309] & b[345])^(a[308] & b[346])^(a[307] & b[347])^(a[306] & b[348])^(a[305] & b[349])^(a[304] & b[350])^(a[303] & b[351])^(a[302] & b[352])^(a[301] & b[353])^(a[300] & b[354])^(a[299] & b[355])^(a[298] & b[356])^(a[297] & b[357])^(a[296] & b[358])^(a[295] & b[359])^(a[294] & b[360])^(a[293] & b[361])^(a[292] & b[362])^(a[291] & b[363])^(a[290] & b[364])^(a[289] & b[365])^(a[288] & b[366])^(a[287] & b[367])^(a[286] & b[368])^(a[285] & b[369])^(a[284] & b[370])^(a[283] & b[371])^(a[282] & b[372])^(a[281] & b[373])^(a[280] & b[374])^(a[279] & b[375])^(a[278] & b[376])^(a[277] & b[377])^(a[276] & b[378])^(a[275] & b[379])^(a[274] & b[380])^(a[273] & b[381])^(a[272] & b[382])^(a[271] & b[383])^(a[270] & b[384])^(a[269] & b[385])^(a[268] & b[386])^(a[267] & b[387])^(a[266] & b[388])^(a[265] & b[389])^(a[264] & b[390])^(a[263] & b[391])^(a[262] & b[392])^(a[261] & b[393])^(a[260] & b[394])^(a[259] & b[395])^(a[258] & b[396])^(a[257] & b[397])^(a[256] & b[398])^(a[255] & b[399])^(a[254] & b[400])^(a[253] & b[401])^(a[252] & b[402])^(a[251] & b[403])^(a[250] & b[404])^(a[249] & b[405])^(a[248] & b[406])^(a[247] & b[407])^(a[246] & b[408]);
assign y[655] = (a[408] & b[247])^(a[407] & b[248])^(a[406] & b[249])^(a[405] & b[250])^(a[404] & b[251])^(a[403] & b[252])^(a[402] & b[253])^(a[401] & b[254])^(a[400] & b[255])^(a[399] & b[256])^(a[398] & b[257])^(a[397] & b[258])^(a[396] & b[259])^(a[395] & b[260])^(a[394] & b[261])^(a[393] & b[262])^(a[392] & b[263])^(a[391] & b[264])^(a[390] & b[265])^(a[389] & b[266])^(a[388] & b[267])^(a[387] & b[268])^(a[386] & b[269])^(a[385] & b[270])^(a[384] & b[271])^(a[383] & b[272])^(a[382] & b[273])^(a[381] & b[274])^(a[380] & b[275])^(a[379] & b[276])^(a[378] & b[277])^(a[377] & b[278])^(a[376] & b[279])^(a[375] & b[280])^(a[374] & b[281])^(a[373] & b[282])^(a[372] & b[283])^(a[371] & b[284])^(a[370] & b[285])^(a[369] & b[286])^(a[368] & b[287])^(a[367] & b[288])^(a[366] & b[289])^(a[365] & b[290])^(a[364] & b[291])^(a[363] & b[292])^(a[362] & b[293])^(a[361] & b[294])^(a[360] & b[295])^(a[359] & b[296])^(a[358] & b[297])^(a[357] & b[298])^(a[356] & b[299])^(a[355] & b[300])^(a[354] & b[301])^(a[353] & b[302])^(a[352] & b[303])^(a[351] & b[304])^(a[350] & b[305])^(a[349] & b[306])^(a[348] & b[307])^(a[347] & b[308])^(a[346] & b[309])^(a[345] & b[310])^(a[344] & b[311])^(a[343] & b[312])^(a[342] & b[313])^(a[341] & b[314])^(a[340] & b[315])^(a[339] & b[316])^(a[338] & b[317])^(a[337] & b[318])^(a[336] & b[319])^(a[335] & b[320])^(a[334] & b[321])^(a[333] & b[322])^(a[332] & b[323])^(a[331] & b[324])^(a[330] & b[325])^(a[329] & b[326])^(a[328] & b[327])^(a[327] & b[328])^(a[326] & b[329])^(a[325] & b[330])^(a[324] & b[331])^(a[323] & b[332])^(a[322] & b[333])^(a[321] & b[334])^(a[320] & b[335])^(a[319] & b[336])^(a[318] & b[337])^(a[317] & b[338])^(a[316] & b[339])^(a[315] & b[340])^(a[314] & b[341])^(a[313] & b[342])^(a[312] & b[343])^(a[311] & b[344])^(a[310] & b[345])^(a[309] & b[346])^(a[308] & b[347])^(a[307] & b[348])^(a[306] & b[349])^(a[305] & b[350])^(a[304] & b[351])^(a[303] & b[352])^(a[302] & b[353])^(a[301] & b[354])^(a[300] & b[355])^(a[299] & b[356])^(a[298] & b[357])^(a[297] & b[358])^(a[296] & b[359])^(a[295] & b[360])^(a[294] & b[361])^(a[293] & b[362])^(a[292] & b[363])^(a[291] & b[364])^(a[290] & b[365])^(a[289] & b[366])^(a[288] & b[367])^(a[287] & b[368])^(a[286] & b[369])^(a[285] & b[370])^(a[284] & b[371])^(a[283] & b[372])^(a[282] & b[373])^(a[281] & b[374])^(a[280] & b[375])^(a[279] & b[376])^(a[278] & b[377])^(a[277] & b[378])^(a[276] & b[379])^(a[275] & b[380])^(a[274] & b[381])^(a[273] & b[382])^(a[272] & b[383])^(a[271] & b[384])^(a[270] & b[385])^(a[269] & b[386])^(a[268] & b[387])^(a[267] & b[388])^(a[266] & b[389])^(a[265] & b[390])^(a[264] & b[391])^(a[263] & b[392])^(a[262] & b[393])^(a[261] & b[394])^(a[260] & b[395])^(a[259] & b[396])^(a[258] & b[397])^(a[257] & b[398])^(a[256] & b[399])^(a[255] & b[400])^(a[254] & b[401])^(a[253] & b[402])^(a[252] & b[403])^(a[251] & b[404])^(a[250] & b[405])^(a[249] & b[406])^(a[248] & b[407])^(a[247] & b[408]);
assign y[656] = (a[408] & b[248])^(a[407] & b[249])^(a[406] & b[250])^(a[405] & b[251])^(a[404] & b[252])^(a[403] & b[253])^(a[402] & b[254])^(a[401] & b[255])^(a[400] & b[256])^(a[399] & b[257])^(a[398] & b[258])^(a[397] & b[259])^(a[396] & b[260])^(a[395] & b[261])^(a[394] & b[262])^(a[393] & b[263])^(a[392] & b[264])^(a[391] & b[265])^(a[390] & b[266])^(a[389] & b[267])^(a[388] & b[268])^(a[387] & b[269])^(a[386] & b[270])^(a[385] & b[271])^(a[384] & b[272])^(a[383] & b[273])^(a[382] & b[274])^(a[381] & b[275])^(a[380] & b[276])^(a[379] & b[277])^(a[378] & b[278])^(a[377] & b[279])^(a[376] & b[280])^(a[375] & b[281])^(a[374] & b[282])^(a[373] & b[283])^(a[372] & b[284])^(a[371] & b[285])^(a[370] & b[286])^(a[369] & b[287])^(a[368] & b[288])^(a[367] & b[289])^(a[366] & b[290])^(a[365] & b[291])^(a[364] & b[292])^(a[363] & b[293])^(a[362] & b[294])^(a[361] & b[295])^(a[360] & b[296])^(a[359] & b[297])^(a[358] & b[298])^(a[357] & b[299])^(a[356] & b[300])^(a[355] & b[301])^(a[354] & b[302])^(a[353] & b[303])^(a[352] & b[304])^(a[351] & b[305])^(a[350] & b[306])^(a[349] & b[307])^(a[348] & b[308])^(a[347] & b[309])^(a[346] & b[310])^(a[345] & b[311])^(a[344] & b[312])^(a[343] & b[313])^(a[342] & b[314])^(a[341] & b[315])^(a[340] & b[316])^(a[339] & b[317])^(a[338] & b[318])^(a[337] & b[319])^(a[336] & b[320])^(a[335] & b[321])^(a[334] & b[322])^(a[333] & b[323])^(a[332] & b[324])^(a[331] & b[325])^(a[330] & b[326])^(a[329] & b[327])^(a[328] & b[328])^(a[327] & b[329])^(a[326] & b[330])^(a[325] & b[331])^(a[324] & b[332])^(a[323] & b[333])^(a[322] & b[334])^(a[321] & b[335])^(a[320] & b[336])^(a[319] & b[337])^(a[318] & b[338])^(a[317] & b[339])^(a[316] & b[340])^(a[315] & b[341])^(a[314] & b[342])^(a[313] & b[343])^(a[312] & b[344])^(a[311] & b[345])^(a[310] & b[346])^(a[309] & b[347])^(a[308] & b[348])^(a[307] & b[349])^(a[306] & b[350])^(a[305] & b[351])^(a[304] & b[352])^(a[303] & b[353])^(a[302] & b[354])^(a[301] & b[355])^(a[300] & b[356])^(a[299] & b[357])^(a[298] & b[358])^(a[297] & b[359])^(a[296] & b[360])^(a[295] & b[361])^(a[294] & b[362])^(a[293] & b[363])^(a[292] & b[364])^(a[291] & b[365])^(a[290] & b[366])^(a[289] & b[367])^(a[288] & b[368])^(a[287] & b[369])^(a[286] & b[370])^(a[285] & b[371])^(a[284] & b[372])^(a[283] & b[373])^(a[282] & b[374])^(a[281] & b[375])^(a[280] & b[376])^(a[279] & b[377])^(a[278] & b[378])^(a[277] & b[379])^(a[276] & b[380])^(a[275] & b[381])^(a[274] & b[382])^(a[273] & b[383])^(a[272] & b[384])^(a[271] & b[385])^(a[270] & b[386])^(a[269] & b[387])^(a[268] & b[388])^(a[267] & b[389])^(a[266] & b[390])^(a[265] & b[391])^(a[264] & b[392])^(a[263] & b[393])^(a[262] & b[394])^(a[261] & b[395])^(a[260] & b[396])^(a[259] & b[397])^(a[258] & b[398])^(a[257] & b[399])^(a[256] & b[400])^(a[255] & b[401])^(a[254] & b[402])^(a[253] & b[403])^(a[252] & b[404])^(a[251] & b[405])^(a[250] & b[406])^(a[249] & b[407])^(a[248] & b[408]);
assign y[657] = (a[408] & b[249])^(a[407] & b[250])^(a[406] & b[251])^(a[405] & b[252])^(a[404] & b[253])^(a[403] & b[254])^(a[402] & b[255])^(a[401] & b[256])^(a[400] & b[257])^(a[399] & b[258])^(a[398] & b[259])^(a[397] & b[260])^(a[396] & b[261])^(a[395] & b[262])^(a[394] & b[263])^(a[393] & b[264])^(a[392] & b[265])^(a[391] & b[266])^(a[390] & b[267])^(a[389] & b[268])^(a[388] & b[269])^(a[387] & b[270])^(a[386] & b[271])^(a[385] & b[272])^(a[384] & b[273])^(a[383] & b[274])^(a[382] & b[275])^(a[381] & b[276])^(a[380] & b[277])^(a[379] & b[278])^(a[378] & b[279])^(a[377] & b[280])^(a[376] & b[281])^(a[375] & b[282])^(a[374] & b[283])^(a[373] & b[284])^(a[372] & b[285])^(a[371] & b[286])^(a[370] & b[287])^(a[369] & b[288])^(a[368] & b[289])^(a[367] & b[290])^(a[366] & b[291])^(a[365] & b[292])^(a[364] & b[293])^(a[363] & b[294])^(a[362] & b[295])^(a[361] & b[296])^(a[360] & b[297])^(a[359] & b[298])^(a[358] & b[299])^(a[357] & b[300])^(a[356] & b[301])^(a[355] & b[302])^(a[354] & b[303])^(a[353] & b[304])^(a[352] & b[305])^(a[351] & b[306])^(a[350] & b[307])^(a[349] & b[308])^(a[348] & b[309])^(a[347] & b[310])^(a[346] & b[311])^(a[345] & b[312])^(a[344] & b[313])^(a[343] & b[314])^(a[342] & b[315])^(a[341] & b[316])^(a[340] & b[317])^(a[339] & b[318])^(a[338] & b[319])^(a[337] & b[320])^(a[336] & b[321])^(a[335] & b[322])^(a[334] & b[323])^(a[333] & b[324])^(a[332] & b[325])^(a[331] & b[326])^(a[330] & b[327])^(a[329] & b[328])^(a[328] & b[329])^(a[327] & b[330])^(a[326] & b[331])^(a[325] & b[332])^(a[324] & b[333])^(a[323] & b[334])^(a[322] & b[335])^(a[321] & b[336])^(a[320] & b[337])^(a[319] & b[338])^(a[318] & b[339])^(a[317] & b[340])^(a[316] & b[341])^(a[315] & b[342])^(a[314] & b[343])^(a[313] & b[344])^(a[312] & b[345])^(a[311] & b[346])^(a[310] & b[347])^(a[309] & b[348])^(a[308] & b[349])^(a[307] & b[350])^(a[306] & b[351])^(a[305] & b[352])^(a[304] & b[353])^(a[303] & b[354])^(a[302] & b[355])^(a[301] & b[356])^(a[300] & b[357])^(a[299] & b[358])^(a[298] & b[359])^(a[297] & b[360])^(a[296] & b[361])^(a[295] & b[362])^(a[294] & b[363])^(a[293] & b[364])^(a[292] & b[365])^(a[291] & b[366])^(a[290] & b[367])^(a[289] & b[368])^(a[288] & b[369])^(a[287] & b[370])^(a[286] & b[371])^(a[285] & b[372])^(a[284] & b[373])^(a[283] & b[374])^(a[282] & b[375])^(a[281] & b[376])^(a[280] & b[377])^(a[279] & b[378])^(a[278] & b[379])^(a[277] & b[380])^(a[276] & b[381])^(a[275] & b[382])^(a[274] & b[383])^(a[273] & b[384])^(a[272] & b[385])^(a[271] & b[386])^(a[270] & b[387])^(a[269] & b[388])^(a[268] & b[389])^(a[267] & b[390])^(a[266] & b[391])^(a[265] & b[392])^(a[264] & b[393])^(a[263] & b[394])^(a[262] & b[395])^(a[261] & b[396])^(a[260] & b[397])^(a[259] & b[398])^(a[258] & b[399])^(a[257] & b[400])^(a[256] & b[401])^(a[255] & b[402])^(a[254] & b[403])^(a[253] & b[404])^(a[252] & b[405])^(a[251] & b[406])^(a[250] & b[407])^(a[249] & b[408]);
assign y[658] = (a[408] & b[250])^(a[407] & b[251])^(a[406] & b[252])^(a[405] & b[253])^(a[404] & b[254])^(a[403] & b[255])^(a[402] & b[256])^(a[401] & b[257])^(a[400] & b[258])^(a[399] & b[259])^(a[398] & b[260])^(a[397] & b[261])^(a[396] & b[262])^(a[395] & b[263])^(a[394] & b[264])^(a[393] & b[265])^(a[392] & b[266])^(a[391] & b[267])^(a[390] & b[268])^(a[389] & b[269])^(a[388] & b[270])^(a[387] & b[271])^(a[386] & b[272])^(a[385] & b[273])^(a[384] & b[274])^(a[383] & b[275])^(a[382] & b[276])^(a[381] & b[277])^(a[380] & b[278])^(a[379] & b[279])^(a[378] & b[280])^(a[377] & b[281])^(a[376] & b[282])^(a[375] & b[283])^(a[374] & b[284])^(a[373] & b[285])^(a[372] & b[286])^(a[371] & b[287])^(a[370] & b[288])^(a[369] & b[289])^(a[368] & b[290])^(a[367] & b[291])^(a[366] & b[292])^(a[365] & b[293])^(a[364] & b[294])^(a[363] & b[295])^(a[362] & b[296])^(a[361] & b[297])^(a[360] & b[298])^(a[359] & b[299])^(a[358] & b[300])^(a[357] & b[301])^(a[356] & b[302])^(a[355] & b[303])^(a[354] & b[304])^(a[353] & b[305])^(a[352] & b[306])^(a[351] & b[307])^(a[350] & b[308])^(a[349] & b[309])^(a[348] & b[310])^(a[347] & b[311])^(a[346] & b[312])^(a[345] & b[313])^(a[344] & b[314])^(a[343] & b[315])^(a[342] & b[316])^(a[341] & b[317])^(a[340] & b[318])^(a[339] & b[319])^(a[338] & b[320])^(a[337] & b[321])^(a[336] & b[322])^(a[335] & b[323])^(a[334] & b[324])^(a[333] & b[325])^(a[332] & b[326])^(a[331] & b[327])^(a[330] & b[328])^(a[329] & b[329])^(a[328] & b[330])^(a[327] & b[331])^(a[326] & b[332])^(a[325] & b[333])^(a[324] & b[334])^(a[323] & b[335])^(a[322] & b[336])^(a[321] & b[337])^(a[320] & b[338])^(a[319] & b[339])^(a[318] & b[340])^(a[317] & b[341])^(a[316] & b[342])^(a[315] & b[343])^(a[314] & b[344])^(a[313] & b[345])^(a[312] & b[346])^(a[311] & b[347])^(a[310] & b[348])^(a[309] & b[349])^(a[308] & b[350])^(a[307] & b[351])^(a[306] & b[352])^(a[305] & b[353])^(a[304] & b[354])^(a[303] & b[355])^(a[302] & b[356])^(a[301] & b[357])^(a[300] & b[358])^(a[299] & b[359])^(a[298] & b[360])^(a[297] & b[361])^(a[296] & b[362])^(a[295] & b[363])^(a[294] & b[364])^(a[293] & b[365])^(a[292] & b[366])^(a[291] & b[367])^(a[290] & b[368])^(a[289] & b[369])^(a[288] & b[370])^(a[287] & b[371])^(a[286] & b[372])^(a[285] & b[373])^(a[284] & b[374])^(a[283] & b[375])^(a[282] & b[376])^(a[281] & b[377])^(a[280] & b[378])^(a[279] & b[379])^(a[278] & b[380])^(a[277] & b[381])^(a[276] & b[382])^(a[275] & b[383])^(a[274] & b[384])^(a[273] & b[385])^(a[272] & b[386])^(a[271] & b[387])^(a[270] & b[388])^(a[269] & b[389])^(a[268] & b[390])^(a[267] & b[391])^(a[266] & b[392])^(a[265] & b[393])^(a[264] & b[394])^(a[263] & b[395])^(a[262] & b[396])^(a[261] & b[397])^(a[260] & b[398])^(a[259] & b[399])^(a[258] & b[400])^(a[257] & b[401])^(a[256] & b[402])^(a[255] & b[403])^(a[254] & b[404])^(a[253] & b[405])^(a[252] & b[406])^(a[251] & b[407])^(a[250] & b[408]);
assign y[659] = (a[408] & b[251])^(a[407] & b[252])^(a[406] & b[253])^(a[405] & b[254])^(a[404] & b[255])^(a[403] & b[256])^(a[402] & b[257])^(a[401] & b[258])^(a[400] & b[259])^(a[399] & b[260])^(a[398] & b[261])^(a[397] & b[262])^(a[396] & b[263])^(a[395] & b[264])^(a[394] & b[265])^(a[393] & b[266])^(a[392] & b[267])^(a[391] & b[268])^(a[390] & b[269])^(a[389] & b[270])^(a[388] & b[271])^(a[387] & b[272])^(a[386] & b[273])^(a[385] & b[274])^(a[384] & b[275])^(a[383] & b[276])^(a[382] & b[277])^(a[381] & b[278])^(a[380] & b[279])^(a[379] & b[280])^(a[378] & b[281])^(a[377] & b[282])^(a[376] & b[283])^(a[375] & b[284])^(a[374] & b[285])^(a[373] & b[286])^(a[372] & b[287])^(a[371] & b[288])^(a[370] & b[289])^(a[369] & b[290])^(a[368] & b[291])^(a[367] & b[292])^(a[366] & b[293])^(a[365] & b[294])^(a[364] & b[295])^(a[363] & b[296])^(a[362] & b[297])^(a[361] & b[298])^(a[360] & b[299])^(a[359] & b[300])^(a[358] & b[301])^(a[357] & b[302])^(a[356] & b[303])^(a[355] & b[304])^(a[354] & b[305])^(a[353] & b[306])^(a[352] & b[307])^(a[351] & b[308])^(a[350] & b[309])^(a[349] & b[310])^(a[348] & b[311])^(a[347] & b[312])^(a[346] & b[313])^(a[345] & b[314])^(a[344] & b[315])^(a[343] & b[316])^(a[342] & b[317])^(a[341] & b[318])^(a[340] & b[319])^(a[339] & b[320])^(a[338] & b[321])^(a[337] & b[322])^(a[336] & b[323])^(a[335] & b[324])^(a[334] & b[325])^(a[333] & b[326])^(a[332] & b[327])^(a[331] & b[328])^(a[330] & b[329])^(a[329] & b[330])^(a[328] & b[331])^(a[327] & b[332])^(a[326] & b[333])^(a[325] & b[334])^(a[324] & b[335])^(a[323] & b[336])^(a[322] & b[337])^(a[321] & b[338])^(a[320] & b[339])^(a[319] & b[340])^(a[318] & b[341])^(a[317] & b[342])^(a[316] & b[343])^(a[315] & b[344])^(a[314] & b[345])^(a[313] & b[346])^(a[312] & b[347])^(a[311] & b[348])^(a[310] & b[349])^(a[309] & b[350])^(a[308] & b[351])^(a[307] & b[352])^(a[306] & b[353])^(a[305] & b[354])^(a[304] & b[355])^(a[303] & b[356])^(a[302] & b[357])^(a[301] & b[358])^(a[300] & b[359])^(a[299] & b[360])^(a[298] & b[361])^(a[297] & b[362])^(a[296] & b[363])^(a[295] & b[364])^(a[294] & b[365])^(a[293] & b[366])^(a[292] & b[367])^(a[291] & b[368])^(a[290] & b[369])^(a[289] & b[370])^(a[288] & b[371])^(a[287] & b[372])^(a[286] & b[373])^(a[285] & b[374])^(a[284] & b[375])^(a[283] & b[376])^(a[282] & b[377])^(a[281] & b[378])^(a[280] & b[379])^(a[279] & b[380])^(a[278] & b[381])^(a[277] & b[382])^(a[276] & b[383])^(a[275] & b[384])^(a[274] & b[385])^(a[273] & b[386])^(a[272] & b[387])^(a[271] & b[388])^(a[270] & b[389])^(a[269] & b[390])^(a[268] & b[391])^(a[267] & b[392])^(a[266] & b[393])^(a[265] & b[394])^(a[264] & b[395])^(a[263] & b[396])^(a[262] & b[397])^(a[261] & b[398])^(a[260] & b[399])^(a[259] & b[400])^(a[258] & b[401])^(a[257] & b[402])^(a[256] & b[403])^(a[255] & b[404])^(a[254] & b[405])^(a[253] & b[406])^(a[252] & b[407])^(a[251] & b[408]);
assign y[660] = (a[408] & b[252])^(a[407] & b[253])^(a[406] & b[254])^(a[405] & b[255])^(a[404] & b[256])^(a[403] & b[257])^(a[402] & b[258])^(a[401] & b[259])^(a[400] & b[260])^(a[399] & b[261])^(a[398] & b[262])^(a[397] & b[263])^(a[396] & b[264])^(a[395] & b[265])^(a[394] & b[266])^(a[393] & b[267])^(a[392] & b[268])^(a[391] & b[269])^(a[390] & b[270])^(a[389] & b[271])^(a[388] & b[272])^(a[387] & b[273])^(a[386] & b[274])^(a[385] & b[275])^(a[384] & b[276])^(a[383] & b[277])^(a[382] & b[278])^(a[381] & b[279])^(a[380] & b[280])^(a[379] & b[281])^(a[378] & b[282])^(a[377] & b[283])^(a[376] & b[284])^(a[375] & b[285])^(a[374] & b[286])^(a[373] & b[287])^(a[372] & b[288])^(a[371] & b[289])^(a[370] & b[290])^(a[369] & b[291])^(a[368] & b[292])^(a[367] & b[293])^(a[366] & b[294])^(a[365] & b[295])^(a[364] & b[296])^(a[363] & b[297])^(a[362] & b[298])^(a[361] & b[299])^(a[360] & b[300])^(a[359] & b[301])^(a[358] & b[302])^(a[357] & b[303])^(a[356] & b[304])^(a[355] & b[305])^(a[354] & b[306])^(a[353] & b[307])^(a[352] & b[308])^(a[351] & b[309])^(a[350] & b[310])^(a[349] & b[311])^(a[348] & b[312])^(a[347] & b[313])^(a[346] & b[314])^(a[345] & b[315])^(a[344] & b[316])^(a[343] & b[317])^(a[342] & b[318])^(a[341] & b[319])^(a[340] & b[320])^(a[339] & b[321])^(a[338] & b[322])^(a[337] & b[323])^(a[336] & b[324])^(a[335] & b[325])^(a[334] & b[326])^(a[333] & b[327])^(a[332] & b[328])^(a[331] & b[329])^(a[330] & b[330])^(a[329] & b[331])^(a[328] & b[332])^(a[327] & b[333])^(a[326] & b[334])^(a[325] & b[335])^(a[324] & b[336])^(a[323] & b[337])^(a[322] & b[338])^(a[321] & b[339])^(a[320] & b[340])^(a[319] & b[341])^(a[318] & b[342])^(a[317] & b[343])^(a[316] & b[344])^(a[315] & b[345])^(a[314] & b[346])^(a[313] & b[347])^(a[312] & b[348])^(a[311] & b[349])^(a[310] & b[350])^(a[309] & b[351])^(a[308] & b[352])^(a[307] & b[353])^(a[306] & b[354])^(a[305] & b[355])^(a[304] & b[356])^(a[303] & b[357])^(a[302] & b[358])^(a[301] & b[359])^(a[300] & b[360])^(a[299] & b[361])^(a[298] & b[362])^(a[297] & b[363])^(a[296] & b[364])^(a[295] & b[365])^(a[294] & b[366])^(a[293] & b[367])^(a[292] & b[368])^(a[291] & b[369])^(a[290] & b[370])^(a[289] & b[371])^(a[288] & b[372])^(a[287] & b[373])^(a[286] & b[374])^(a[285] & b[375])^(a[284] & b[376])^(a[283] & b[377])^(a[282] & b[378])^(a[281] & b[379])^(a[280] & b[380])^(a[279] & b[381])^(a[278] & b[382])^(a[277] & b[383])^(a[276] & b[384])^(a[275] & b[385])^(a[274] & b[386])^(a[273] & b[387])^(a[272] & b[388])^(a[271] & b[389])^(a[270] & b[390])^(a[269] & b[391])^(a[268] & b[392])^(a[267] & b[393])^(a[266] & b[394])^(a[265] & b[395])^(a[264] & b[396])^(a[263] & b[397])^(a[262] & b[398])^(a[261] & b[399])^(a[260] & b[400])^(a[259] & b[401])^(a[258] & b[402])^(a[257] & b[403])^(a[256] & b[404])^(a[255] & b[405])^(a[254] & b[406])^(a[253] & b[407])^(a[252] & b[408]);
assign y[661] = (a[408] & b[253])^(a[407] & b[254])^(a[406] & b[255])^(a[405] & b[256])^(a[404] & b[257])^(a[403] & b[258])^(a[402] & b[259])^(a[401] & b[260])^(a[400] & b[261])^(a[399] & b[262])^(a[398] & b[263])^(a[397] & b[264])^(a[396] & b[265])^(a[395] & b[266])^(a[394] & b[267])^(a[393] & b[268])^(a[392] & b[269])^(a[391] & b[270])^(a[390] & b[271])^(a[389] & b[272])^(a[388] & b[273])^(a[387] & b[274])^(a[386] & b[275])^(a[385] & b[276])^(a[384] & b[277])^(a[383] & b[278])^(a[382] & b[279])^(a[381] & b[280])^(a[380] & b[281])^(a[379] & b[282])^(a[378] & b[283])^(a[377] & b[284])^(a[376] & b[285])^(a[375] & b[286])^(a[374] & b[287])^(a[373] & b[288])^(a[372] & b[289])^(a[371] & b[290])^(a[370] & b[291])^(a[369] & b[292])^(a[368] & b[293])^(a[367] & b[294])^(a[366] & b[295])^(a[365] & b[296])^(a[364] & b[297])^(a[363] & b[298])^(a[362] & b[299])^(a[361] & b[300])^(a[360] & b[301])^(a[359] & b[302])^(a[358] & b[303])^(a[357] & b[304])^(a[356] & b[305])^(a[355] & b[306])^(a[354] & b[307])^(a[353] & b[308])^(a[352] & b[309])^(a[351] & b[310])^(a[350] & b[311])^(a[349] & b[312])^(a[348] & b[313])^(a[347] & b[314])^(a[346] & b[315])^(a[345] & b[316])^(a[344] & b[317])^(a[343] & b[318])^(a[342] & b[319])^(a[341] & b[320])^(a[340] & b[321])^(a[339] & b[322])^(a[338] & b[323])^(a[337] & b[324])^(a[336] & b[325])^(a[335] & b[326])^(a[334] & b[327])^(a[333] & b[328])^(a[332] & b[329])^(a[331] & b[330])^(a[330] & b[331])^(a[329] & b[332])^(a[328] & b[333])^(a[327] & b[334])^(a[326] & b[335])^(a[325] & b[336])^(a[324] & b[337])^(a[323] & b[338])^(a[322] & b[339])^(a[321] & b[340])^(a[320] & b[341])^(a[319] & b[342])^(a[318] & b[343])^(a[317] & b[344])^(a[316] & b[345])^(a[315] & b[346])^(a[314] & b[347])^(a[313] & b[348])^(a[312] & b[349])^(a[311] & b[350])^(a[310] & b[351])^(a[309] & b[352])^(a[308] & b[353])^(a[307] & b[354])^(a[306] & b[355])^(a[305] & b[356])^(a[304] & b[357])^(a[303] & b[358])^(a[302] & b[359])^(a[301] & b[360])^(a[300] & b[361])^(a[299] & b[362])^(a[298] & b[363])^(a[297] & b[364])^(a[296] & b[365])^(a[295] & b[366])^(a[294] & b[367])^(a[293] & b[368])^(a[292] & b[369])^(a[291] & b[370])^(a[290] & b[371])^(a[289] & b[372])^(a[288] & b[373])^(a[287] & b[374])^(a[286] & b[375])^(a[285] & b[376])^(a[284] & b[377])^(a[283] & b[378])^(a[282] & b[379])^(a[281] & b[380])^(a[280] & b[381])^(a[279] & b[382])^(a[278] & b[383])^(a[277] & b[384])^(a[276] & b[385])^(a[275] & b[386])^(a[274] & b[387])^(a[273] & b[388])^(a[272] & b[389])^(a[271] & b[390])^(a[270] & b[391])^(a[269] & b[392])^(a[268] & b[393])^(a[267] & b[394])^(a[266] & b[395])^(a[265] & b[396])^(a[264] & b[397])^(a[263] & b[398])^(a[262] & b[399])^(a[261] & b[400])^(a[260] & b[401])^(a[259] & b[402])^(a[258] & b[403])^(a[257] & b[404])^(a[256] & b[405])^(a[255] & b[406])^(a[254] & b[407])^(a[253] & b[408]);
assign y[662] = (a[408] & b[254])^(a[407] & b[255])^(a[406] & b[256])^(a[405] & b[257])^(a[404] & b[258])^(a[403] & b[259])^(a[402] & b[260])^(a[401] & b[261])^(a[400] & b[262])^(a[399] & b[263])^(a[398] & b[264])^(a[397] & b[265])^(a[396] & b[266])^(a[395] & b[267])^(a[394] & b[268])^(a[393] & b[269])^(a[392] & b[270])^(a[391] & b[271])^(a[390] & b[272])^(a[389] & b[273])^(a[388] & b[274])^(a[387] & b[275])^(a[386] & b[276])^(a[385] & b[277])^(a[384] & b[278])^(a[383] & b[279])^(a[382] & b[280])^(a[381] & b[281])^(a[380] & b[282])^(a[379] & b[283])^(a[378] & b[284])^(a[377] & b[285])^(a[376] & b[286])^(a[375] & b[287])^(a[374] & b[288])^(a[373] & b[289])^(a[372] & b[290])^(a[371] & b[291])^(a[370] & b[292])^(a[369] & b[293])^(a[368] & b[294])^(a[367] & b[295])^(a[366] & b[296])^(a[365] & b[297])^(a[364] & b[298])^(a[363] & b[299])^(a[362] & b[300])^(a[361] & b[301])^(a[360] & b[302])^(a[359] & b[303])^(a[358] & b[304])^(a[357] & b[305])^(a[356] & b[306])^(a[355] & b[307])^(a[354] & b[308])^(a[353] & b[309])^(a[352] & b[310])^(a[351] & b[311])^(a[350] & b[312])^(a[349] & b[313])^(a[348] & b[314])^(a[347] & b[315])^(a[346] & b[316])^(a[345] & b[317])^(a[344] & b[318])^(a[343] & b[319])^(a[342] & b[320])^(a[341] & b[321])^(a[340] & b[322])^(a[339] & b[323])^(a[338] & b[324])^(a[337] & b[325])^(a[336] & b[326])^(a[335] & b[327])^(a[334] & b[328])^(a[333] & b[329])^(a[332] & b[330])^(a[331] & b[331])^(a[330] & b[332])^(a[329] & b[333])^(a[328] & b[334])^(a[327] & b[335])^(a[326] & b[336])^(a[325] & b[337])^(a[324] & b[338])^(a[323] & b[339])^(a[322] & b[340])^(a[321] & b[341])^(a[320] & b[342])^(a[319] & b[343])^(a[318] & b[344])^(a[317] & b[345])^(a[316] & b[346])^(a[315] & b[347])^(a[314] & b[348])^(a[313] & b[349])^(a[312] & b[350])^(a[311] & b[351])^(a[310] & b[352])^(a[309] & b[353])^(a[308] & b[354])^(a[307] & b[355])^(a[306] & b[356])^(a[305] & b[357])^(a[304] & b[358])^(a[303] & b[359])^(a[302] & b[360])^(a[301] & b[361])^(a[300] & b[362])^(a[299] & b[363])^(a[298] & b[364])^(a[297] & b[365])^(a[296] & b[366])^(a[295] & b[367])^(a[294] & b[368])^(a[293] & b[369])^(a[292] & b[370])^(a[291] & b[371])^(a[290] & b[372])^(a[289] & b[373])^(a[288] & b[374])^(a[287] & b[375])^(a[286] & b[376])^(a[285] & b[377])^(a[284] & b[378])^(a[283] & b[379])^(a[282] & b[380])^(a[281] & b[381])^(a[280] & b[382])^(a[279] & b[383])^(a[278] & b[384])^(a[277] & b[385])^(a[276] & b[386])^(a[275] & b[387])^(a[274] & b[388])^(a[273] & b[389])^(a[272] & b[390])^(a[271] & b[391])^(a[270] & b[392])^(a[269] & b[393])^(a[268] & b[394])^(a[267] & b[395])^(a[266] & b[396])^(a[265] & b[397])^(a[264] & b[398])^(a[263] & b[399])^(a[262] & b[400])^(a[261] & b[401])^(a[260] & b[402])^(a[259] & b[403])^(a[258] & b[404])^(a[257] & b[405])^(a[256] & b[406])^(a[255] & b[407])^(a[254] & b[408]);
assign y[663] = (a[408] & b[255])^(a[407] & b[256])^(a[406] & b[257])^(a[405] & b[258])^(a[404] & b[259])^(a[403] & b[260])^(a[402] & b[261])^(a[401] & b[262])^(a[400] & b[263])^(a[399] & b[264])^(a[398] & b[265])^(a[397] & b[266])^(a[396] & b[267])^(a[395] & b[268])^(a[394] & b[269])^(a[393] & b[270])^(a[392] & b[271])^(a[391] & b[272])^(a[390] & b[273])^(a[389] & b[274])^(a[388] & b[275])^(a[387] & b[276])^(a[386] & b[277])^(a[385] & b[278])^(a[384] & b[279])^(a[383] & b[280])^(a[382] & b[281])^(a[381] & b[282])^(a[380] & b[283])^(a[379] & b[284])^(a[378] & b[285])^(a[377] & b[286])^(a[376] & b[287])^(a[375] & b[288])^(a[374] & b[289])^(a[373] & b[290])^(a[372] & b[291])^(a[371] & b[292])^(a[370] & b[293])^(a[369] & b[294])^(a[368] & b[295])^(a[367] & b[296])^(a[366] & b[297])^(a[365] & b[298])^(a[364] & b[299])^(a[363] & b[300])^(a[362] & b[301])^(a[361] & b[302])^(a[360] & b[303])^(a[359] & b[304])^(a[358] & b[305])^(a[357] & b[306])^(a[356] & b[307])^(a[355] & b[308])^(a[354] & b[309])^(a[353] & b[310])^(a[352] & b[311])^(a[351] & b[312])^(a[350] & b[313])^(a[349] & b[314])^(a[348] & b[315])^(a[347] & b[316])^(a[346] & b[317])^(a[345] & b[318])^(a[344] & b[319])^(a[343] & b[320])^(a[342] & b[321])^(a[341] & b[322])^(a[340] & b[323])^(a[339] & b[324])^(a[338] & b[325])^(a[337] & b[326])^(a[336] & b[327])^(a[335] & b[328])^(a[334] & b[329])^(a[333] & b[330])^(a[332] & b[331])^(a[331] & b[332])^(a[330] & b[333])^(a[329] & b[334])^(a[328] & b[335])^(a[327] & b[336])^(a[326] & b[337])^(a[325] & b[338])^(a[324] & b[339])^(a[323] & b[340])^(a[322] & b[341])^(a[321] & b[342])^(a[320] & b[343])^(a[319] & b[344])^(a[318] & b[345])^(a[317] & b[346])^(a[316] & b[347])^(a[315] & b[348])^(a[314] & b[349])^(a[313] & b[350])^(a[312] & b[351])^(a[311] & b[352])^(a[310] & b[353])^(a[309] & b[354])^(a[308] & b[355])^(a[307] & b[356])^(a[306] & b[357])^(a[305] & b[358])^(a[304] & b[359])^(a[303] & b[360])^(a[302] & b[361])^(a[301] & b[362])^(a[300] & b[363])^(a[299] & b[364])^(a[298] & b[365])^(a[297] & b[366])^(a[296] & b[367])^(a[295] & b[368])^(a[294] & b[369])^(a[293] & b[370])^(a[292] & b[371])^(a[291] & b[372])^(a[290] & b[373])^(a[289] & b[374])^(a[288] & b[375])^(a[287] & b[376])^(a[286] & b[377])^(a[285] & b[378])^(a[284] & b[379])^(a[283] & b[380])^(a[282] & b[381])^(a[281] & b[382])^(a[280] & b[383])^(a[279] & b[384])^(a[278] & b[385])^(a[277] & b[386])^(a[276] & b[387])^(a[275] & b[388])^(a[274] & b[389])^(a[273] & b[390])^(a[272] & b[391])^(a[271] & b[392])^(a[270] & b[393])^(a[269] & b[394])^(a[268] & b[395])^(a[267] & b[396])^(a[266] & b[397])^(a[265] & b[398])^(a[264] & b[399])^(a[263] & b[400])^(a[262] & b[401])^(a[261] & b[402])^(a[260] & b[403])^(a[259] & b[404])^(a[258] & b[405])^(a[257] & b[406])^(a[256] & b[407])^(a[255] & b[408]);
assign y[664] = (a[408] & b[256])^(a[407] & b[257])^(a[406] & b[258])^(a[405] & b[259])^(a[404] & b[260])^(a[403] & b[261])^(a[402] & b[262])^(a[401] & b[263])^(a[400] & b[264])^(a[399] & b[265])^(a[398] & b[266])^(a[397] & b[267])^(a[396] & b[268])^(a[395] & b[269])^(a[394] & b[270])^(a[393] & b[271])^(a[392] & b[272])^(a[391] & b[273])^(a[390] & b[274])^(a[389] & b[275])^(a[388] & b[276])^(a[387] & b[277])^(a[386] & b[278])^(a[385] & b[279])^(a[384] & b[280])^(a[383] & b[281])^(a[382] & b[282])^(a[381] & b[283])^(a[380] & b[284])^(a[379] & b[285])^(a[378] & b[286])^(a[377] & b[287])^(a[376] & b[288])^(a[375] & b[289])^(a[374] & b[290])^(a[373] & b[291])^(a[372] & b[292])^(a[371] & b[293])^(a[370] & b[294])^(a[369] & b[295])^(a[368] & b[296])^(a[367] & b[297])^(a[366] & b[298])^(a[365] & b[299])^(a[364] & b[300])^(a[363] & b[301])^(a[362] & b[302])^(a[361] & b[303])^(a[360] & b[304])^(a[359] & b[305])^(a[358] & b[306])^(a[357] & b[307])^(a[356] & b[308])^(a[355] & b[309])^(a[354] & b[310])^(a[353] & b[311])^(a[352] & b[312])^(a[351] & b[313])^(a[350] & b[314])^(a[349] & b[315])^(a[348] & b[316])^(a[347] & b[317])^(a[346] & b[318])^(a[345] & b[319])^(a[344] & b[320])^(a[343] & b[321])^(a[342] & b[322])^(a[341] & b[323])^(a[340] & b[324])^(a[339] & b[325])^(a[338] & b[326])^(a[337] & b[327])^(a[336] & b[328])^(a[335] & b[329])^(a[334] & b[330])^(a[333] & b[331])^(a[332] & b[332])^(a[331] & b[333])^(a[330] & b[334])^(a[329] & b[335])^(a[328] & b[336])^(a[327] & b[337])^(a[326] & b[338])^(a[325] & b[339])^(a[324] & b[340])^(a[323] & b[341])^(a[322] & b[342])^(a[321] & b[343])^(a[320] & b[344])^(a[319] & b[345])^(a[318] & b[346])^(a[317] & b[347])^(a[316] & b[348])^(a[315] & b[349])^(a[314] & b[350])^(a[313] & b[351])^(a[312] & b[352])^(a[311] & b[353])^(a[310] & b[354])^(a[309] & b[355])^(a[308] & b[356])^(a[307] & b[357])^(a[306] & b[358])^(a[305] & b[359])^(a[304] & b[360])^(a[303] & b[361])^(a[302] & b[362])^(a[301] & b[363])^(a[300] & b[364])^(a[299] & b[365])^(a[298] & b[366])^(a[297] & b[367])^(a[296] & b[368])^(a[295] & b[369])^(a[294] & b[370])^(a[293] & b[371])^(a[292] & b[372])^(a[291] & b[373])^(a[290] & b[374])^(a[289] & b[375])^(a[288] & b[376])^(a[287] & b[377])^(a[286] & b[378])^(a[285] & b[379])^(a[284] & b[380])^(a[283] & b[381])^(a[282] & b[382])^(a[281] & b[383])^(a[280] & b[384])^(a[279] & b[385])^(a[278] & b[386])^(a[277] & b[387])^(a[276] & b[388])^(a[275] & b[389])^(a[274] & b[390])^(a[273] & b[391])^(a[272] & b[392])^(a[271] & b[393])^(a[270] & b[394])^(a[269] & b[395])^(a[268] & b[396])^(a[267] & b[397])^(a[266] & b[398])^(a[265] & b[399])^(a[264] & b[400])^(a[263] & b[401])^(a[262] & b[402])^(a[261] & b[403])^(a[260] & b[404])^(a[259] & b[405])^(a[258] & b[406])^(a[257] & b[407])^(a[256] & b[408]);
assign y[665] = (a[408] & b[257])^(a[407] & b[258])^(a[406] & b[259])^(a[405] & b[260])^(a[404] & b[261])^(a[403] & b[262])^(a[402] & b[263])^(a[401] & b[264])^(a[400] & b[265])^(a[399] & b[266])^(a[398] & b[267])^(a[397] & b[268])^(a[396] & b[269])^(a[395] & b[270])^(a[394] & b[271])^(a[393] & b[272])^(a[392] & b[273])^(a[391] & b[274])^(a[390] & b[275])^(a[389] & b[276])^(a[388] & b[277])^(a[387] & b[278])^(a[386] & b[279])^(a[385] & b[280])^(a[384] & b[281])^(a[383] & b[282])^(a[382] & b[283])^(a[381] & b[284])^(a[380] & b[285])^(a[379] & b[286])^(a[378] & b[287])^(a[377] & b[288])^(a[376] & b[289])^(a[375] & b[290])^(a[374] & b[291])^(a[373] & b[292])^(a[372] & b[293])^(a[371] & b[294])^(a[370] & b[295])^(a[369] & b[296])^(a[368] & b[297])^(a[367] & b[298])^(a[366] & b[299])^(a[365] & b[300])^(a[364] & b[301])^(a[363] & b[302])^(a[362] & b[303])^(a[361] & b[304])^(a[360] & b[305])^(a[359] & b[306])^(a[358] & b[307])^(a[357] & b[308])^(a[356] & b[309])^(a[355] & b[310])^(a[354] & b[311])^(a[353] & b[312])^(a[352] & b[313])^(a[351] & b[314])^(a[350] & b[315])^(a[349] & b[316])^(a[348] & b[317])^(a[347] & b[318])^(a[346] & b[319])^(a[345] & b[320])^(a[344] & b[321])^(a[343] & b[322])^(a[342] & b[323])^(a[341] & b[324])^(a[340] & b[325])^(a[339] & b[326])^(a[338] & b[327])^(a[337] & b[328])^(a[336] & b[329])^(a[335] & b[330])^(a[334] & b[331])^(a[333] & b[332])^(a[332] & b[333])^(a[331] & b[334])^(a[330] & b[335])^(a[329] & b[336])^(a[328] & b[337])^(a[327] & b[338])^(a[326] & b[339])^(a[325] & b[340])^(a[324] & b[341])^(a[323] & b[342])^(a[322] & b[343])^(a[321] & b[344])^(a[320] & b[345])^(a[319] & b[346])^(a[318] & b[347])^(a[317] & b[348])^(a[316] & b[349])^(a[315] & b[350])^(a[314] & b[351])^(a[313] & b[352])^(a[312] & b[353])^(a[311] & b[354])^(a[310] & b[355])^(a[309] & b[356])^(a[308] & b[357])^(a[307] & b[358])^(a[306] & b[359])^(a[305] & b[360])^(a[304] & b[361])^(a[303] & b[362])^(a[302] & b[363])^(a[301] & b[364])^(a[300] & b[365])^(a[299] & b[366])^(a[298] & b[367])^(a[297] & b[368])^(a[296] & b[369])^(a[295] & b[370])^(a[294] & b[371])^(a[293] & b[372])^(a[292] & b[373])^(a[291] & b[374])^(a[290] & b[375])^(a[289] & b[376])^(a[288] & b[377])^(a[287] & b[378])^(a[286] & b[379])^(a[285] & b[380])^(a[284] & b[381])^(a[283] & b[382])^(a[282] & b[383])^(a[281] & b[384])^(a[280] & b[385])^(a[279] & b[386])^(a[278] & b[387])^(a[277] & b[388])^(a[276] & b[389])^(a[275] & b[390])^(a[274] & b[391])^(a[273] & b[392])^(a[272] & b[393])^(a[271] & b[394])^(a[270] & b[395])^(a[269] & b[396])^(a[268] & b[397])^(a[267] & b[398])^(a[266] & b[399])^(a[265] & b[400])^(a[264] & b[401])^(a[263] & b[402])^(a[262] & b[403])^(a[261] & b[404])^(a[260] & b[405])^(a[259] & b[406])^(a[258] & b[407])^(a[257] & b[408]);
assign y[666] = (a[408] & b[258])^(a[407] & b[259])^(a[406] & b[260])^(a[405] & b[261])^(a[404] & b[262])^(a[403] & b[263])^(a[402] & b[264])^(a[401] & b[265])^(a[400] & b[266])^(a[399] & b[267])^(a[398] & b[268])^(a[397] & b[269])^(a[396] & b[270])^(a[395] & b[271])^(a[394] & b[272])^(a[393] & b[273])^(a[392] & b[274])^(a[391] & b[275])^(a[390] & b[276])^(a[389] & b[277])^(a[388] & b[278])^(a[387] & b[279])^(a[386] & b[280])^(a[385] & b[281])^(a[384] & b[282])^(a[383] & b[283])^(a[382] & b[284])^(a[381] & b[285])^(a[380] & b[286])^(a[379] & b[287])^(a[378] & b[288])^(a[377] & b[289])^(a[376] & b[290])^(a[375] & b[291])^(a[374] & b[292])^(a[373] & b[293])^(a[372] & b[294])^(a[371] & b[295])^(a[370] & b[296])^(a[369] & b[297])^(a[368] & b[298])^(a[367] & b[299])^(a[366] & b[300])^(a[365] & b[301])^(a[364] & b[302])^(a[363] & b[303])^(a[362] & b[304])^(a[361] & b[305])^(a[360] & b[306])^(a[359] & b[307])^(a[358] & b[308])^(a[357] & b[309])^(a[356] & b[310])^(a[355] & b[311])^(a[354] & b[312])^(a[353] & b[313])^(a[352] & b[314])^(a[351] & b[315])^(a[350] & b[316])^(a[349] & b[317])^(a[348] & b[318])^(a[347] & b[319])^(a[346] & b[320])^(a[345] & b[321])^(a[344] & b[322])^(a[343] & b[323])^(a[342] & b[324])^(a[341] & b[325])^(a[340] & b[326])^(a[339] & b[327])^(a[338] & b[328])^(a[337] & b[329])^(a[336] & b[330])^(a[335] & b[331])^(a[334] & b[332])^(a[333] & b[333])^(a[332] & b[334])^(a[331] & b[335])^(a[330] & b[336])^(a[329] & b[337])^(a[328] & b[338])^(a[327] & b[339])^(a[326] & b[340])^(a[325] & b[341])^(a[324] & b[342])^(a[323] & b[343])^(a[322] & b[344])^(a[321] & b[345])^(a[320] & b[346])^(a[319] & b[347])^(a[318] & b[348])^(a[317] & b[349])^(a[316] & b[350])^(a[315] & b[351])^(a[314] & b[352])^(a[313] & b[353])^(a[312] & b[354])^(a[311] & b[355])^(a[310] & b[356])^(a[309] & b[357])^(a[308] & b[358])^(a[307] & b[359])^(a[306] & b[360])^(a[305] & b[361])^(a[304] & b[362])^(a[303] & b[363])^(a[302] & b[364])^(a[301] & b[365])^(a[300] & b[366])^(a[299] & b[367])^(a[298] & b[368])^(a[297] & b[369])^(a[296] & b[370])^(a[295] & b[371])^(a[294] & b[372])^(a[293] & b[373])^(a[292] & b[374])^(a[291] & b[375])^(a[290] & b[376])^(a[289] & b[377])^(a[288] & b[378])^(a[287] & b[379])^(a[286] & b[380])^(a[285] & b[381])^(a[284] & b[382])^(a[283] & b[383])^(a[282] & b[384])^(a[281] & b[385])^(a[280] & b[386])^(a[279] & b[387])^(a[278] & b[388])^(a[277] & b[389])^(a[276] & b[390])^(a[275] & b[391])^(a[274] & b[392])^(a[273] & b[393])^(a[272] & b[394])^(a[271] & b[395])^(a[270] & b[396])^(a[269] & b[397])^(a[268] & b[398])^(a[267] & b[399])^(a[266] & b[400])^(a[265] & b[401])^(a[264] & b[402])^(a[263] & b[403])^(a[262] & b[404])^(a[261] & b[405])^(a[260] & b[406])^(a[259] & b[407])^(a[258] & b[408]);
assign y[667] = (a[408] & b[259])^(a[407] & b[260])^(a[406] & b[261])^(a[405] & b[262])^(a[404] & b[263])^(a[403] & b[264])^(a[402] & b[265])^(a[401] & b[266])^(a[400] & b[267])^(a[399] & b[268])^(a[398] & b[269])^(a[397] & b[270])^(a[396] & b[271])^(a[395] & b[272])^(a[394] & b[273])^(a[393] & b[274])^(a[392] & b[275])^(a[391] & b[276])^(a[390] & b[277])^(a[389] & b[278])^(a[388] & b[279])^(a[387] & b[280])^(a[386] & b[281])^(a[385] & b[282])^(a[384] & b[283])^(a[383] & b[284])^(a[382] & b[285])^(a[381] & b[286])^(a[380] & b[287])^(a[379] & b[288])^(a[378] & b[289])^(a[377] & b[290])^(a[376] & b[291])^(a[375] & b[292])^(a[374] & b[293])^(a[373] & b[294])^(a[372] & b[295])^(a[371] & b[296])^(a[370] & b[297])^(a[369] & b[298])^(a[368] & b[299])^(a[367] & b[300])^(a[366] & b[301])^(a[365] & b[302])^(a[364] & b[303])^(a[363] & b[304])^(a[362] & b[305])^(a[361] & b[306])^(a[360] & b[307])^(a[359] & b[308])^(a[358] & b[309])^(a[357] & b[310])^(a[356] & b[311])^(a[355] & b[312])^(a[354] & b[313])^(a[353] & b[314])^(a[352] & b[315])^(a[351] & b[316])^(a[350] & b[317])^(a[349] & b[318])^(a[348] & b[319])^(a[347] & b[320])^(a[346] & b[321])^(a[345] & b[322])^(a[344] & b[323])^(a[343] & b[324])^(a[342] & b[325])^(a[341] & b[326])^(a[340] & b[327])^(a[339] & b[328])^(a[338] & b[329])^(a[337] & b[330])^(a[336] & b[331])^(a[335] & b[332])^(a[334] & b[333])^(a[333] & b[334])^(a[332] & b[335])^(a[331] & b[336])^(a[330] & b[337])^(a[329] & b[338])^(a[328] & b[339])^(a[327] & b[340])^(a[326] & b[341])^(a[325] & b[342])^(a[324] & b[343])^(a[323] & b[344])^(a[322] & b[345])^(a[321] & b[346])^(a[320] & b[347])^(a[319] & b[348])^(a[318] & b[349])^(a[317] & b[350])^(a[316] & b[351])^(a[315] & b[352])^(a[314] & b[353])^(a[313] & b[354])^(a[312] & b[355])^(a[311] & b[356])^(a[310] & b[357])^(a[309] & b[358])^(a[308] & b[359])^(a[307] & b[360])^(a[306] & b[361])^(a[305] & b[362])^(a[304] & b[363])^(a[303] & b[364])^(a[302] & b[365])^(a[301] & b[366])^(a[300] & b[367])^(a[299] & b[368])^(a[298] & b[369])^(a[297] & b[370])^(a[296] & b[371])^(a[295] & b[372])^(a[294] & b[373])^(a[293] & b[374])^(a[292] & b[375])^(a[291] & b[376])^(a[290] & b[377])^(a[289] & b[378])^(a[288] & b[379])^(a[287] & b[380])^(a[286] & b[381])^(a[285] & b[382])^(a[284] & b[383])^(a[283] & b[384])^(a[282] & b[385])^(a[281] & b[386])^(a[280] & b[387])^(a[279] & b[388])^(a[278] & b[389])^(a[277] & b[390])^(a[276] & b[391])^(a[275] & b[392])^(a[274] & b[393])^(a[273] & b[394])^(a[272] & b[395])^(a[271] & b[396])^(a[270] & b[397])^(a[269] & b[398])^(a[268] & b[399])^(a[267] & b[400])^(a[266] & b[401])^(a[265] & b[402])^(a[264] & b[403])^(a[263] & b[404])^(a[262] & b[405])^(a[261] & b[406])^(a[260] & b[407])^(a[259] & b[408]);
assign y[668] = (a[408] & b[260])^(a[407] & b[261])^(a[406] & b[262])^(a[405] & b[263])^(a[404] & b[264])^(a[403] & b[265])^(a[402] & b[266])^(a[401] & b[267])^(a[400] & b[268])^(a[399] & b[269])^(a[398] & b[270])^(a[397] & b[271])^(a[396] & b[272])^(a[395] & b[273])^(a[394] & b[274])^(a[393] & b[275])^(a[392] & b[276])^(a[391] & b[277])^(a[390] & b[278])^(a[389] & b[279])^(a[388] & b[280])^(a[387] & b[281])^(a[386] & b[282])^(a[385] & b[283])^(a[384] & b[284])^(a[383] & b[285])^(a[382] & b[286])^(a[381] & b[287])^(a[380] & b[288])^(a[379] & b[289])^(a[378] & b[290])^(a[377] & b[291])^(a[376] & b[292])^(a[375] & b[293])^(a[374] & b[294])^(a[373] & b[295])^(a[372] & b[296])^(a[371] & b[297])^(a[370] & b[298])^(a[369] & b[299])^(a[368] & b[300])^(a[367] & b[301])^(a[366] & b[302])^(a[365] & b[303])^(a[364] & b[304])^(a[363] & b[305])^(a[362] & b[306])^(a[361] & b[307])^(a[360] & b[308])^(a[359] & b[309])^(a[358] & b[310])^(a[357] & b[311])^(a[356] & b[312])^(a[355] & b[313])^(a[354] & b[314])^(a[353] & b[315])^(a[352] & b[316])^(a[351] & b[317])^(a[350] & b[318])^(a[349] & b[319])^(a[348] & b[320])^(a[347] & b[321])^(a[346] & b[322])^(a[345] & b[323])^(a[344] & b[324])^(a[343] & b[325])^(a[342] & b[326])^(a[341] & b[327])^(a[340] & b[328])^(a[339] & b[329])^(a[338] & b[330])^(a[337] & b[331])^(a[336] & b[332])^(a[335] & b[333])^(a[334] & b[334])^(a[333] & b[335])^(a[332] & b[336])^(a[331] & b[337])^(a[330] & b[338])^(a[329] & b[339])^(a[328] & b[340])^(a[327] & b[341])^(a[326] & b[342])^(a[325] & b[343])^(a[324] & b[344])^(a[323] & b[345])^(a[322] & b[346])^(a[321] & b[347])^(a[320] & b[348])^(a[319] & b[349])^(a[318] & b[350])^(a[317] & b[351])^(a[316] & b[352])^(a[315] & b[353])^(a[314] & b[354])^(a[313] & b[355])^(a[312] & b[356])^(a[311] & b[357])^(a[310] & b[358])^(a[309] & b[359])^(a[308] & b[360])^(a[307] & b[361])^(a[306] & b[362])^(a[305] & b[363])^(a[304] & b[364])^(a[303] & b[365])^(a[302] & b[366])^(a[301] & b[367])^(a[300] & b[368])^(a[299] & b[369])^(a[298] & b[370])^(a[297] & b[371])^(a[296] & b[372])^(a[295] & b[373])^(a[294] & b[374])^(a[293] & b[375])^(a[292] & b[376])^(a[291] & b[377])^(a[290] & b[378])^(a[289] & b[379])^(a[288] & b[380])^(a[287] & b[381])^(a[286] & b[382])^(a[285] & b[383])^(a[284] & b[384])^(a[283] & b[385])^(a[282] & b[386])^(a[281] & b[387])^(a[280] & b[388])^(a[279] & b[389])^(a[278] & b[390])^(a[277] & b[391])^(a[276] & b[392])^(a[275] & b[393])^(a[274] & b[394])^(a[273] & b[395])^(a[272] & b[396])^(a[271] & b[397])^(a[270] & b[398])^(a[269] & b[399])^(a[268] & b[400])^(a[267] & b[401])^(a[266] & b[402])^(a[265] & b[403])^(a[264] & b[404])^(a[263] & b[405])^(a[262] & b[406])^(a[261] & b[407])^(a[260] & b[408]);
assign y[669] = (a[408] & b[261])^(a[407] & b[262])^(a[406] & b[263])^(a[405] & b[264])^(a[404] & b[265])^(a[403] & b[266])^(a[402] & b[267])^(a[401] & b[268])^(a[400] & b[269])^(a[399] & b[270])^(a[398] & b[271])^(a[397] & b[272])^(a[396] & b[273])^(a[395] & b[274])^(a[394] & b[275])^(a[393] & b[276])^(a[392] & b[277])^(a[391] & b[278])^(a[390] & b[279])^(a[389] & b[280])^(a[388] & b[281])^(a[387] & b[282])^(a[386] & b[283])^(a[385] & b[284])^(a[384] & b[285])^(a[383] & b[286])^(a[382] & b[287])^(a[381] & b[288])^(a[380] & b[289])^(a[379] & b[290])^(a[378] & b[291])^(a[377] & b[292])^(a[376] & b[293])^(a[375] & b[294])^(a[374] & b[295])^(a[373] & b[296])^(a[372] & b[297])^(a[371] & b[298])^(a[370] & b[299])^(a[369] & b[300])^(a[368] & b[301])^(a[367] & b[302])^(a[366] & b[303])^(a[365] & b[304])^(a[364] & b[305])^(a[363] & b[306])^(a[362] & b[307])^(a[361] & b[308])^(a[360] & b[309])^(a[359] & b[310])^(a[358] & b[311])^(a[357] & b[312])^(a[356] & b[313])^(a[355] & b[314])^(a[354] & b[315])^(a[353] & b[316])^(a[352] & b[317])^(a[351] & b[318])^(a[350] & b[319])^(a[349] & b[320])^(a[348] & b[321])^(a[347] & b[322])^(a[346] & b[323])^(a[345] & b[324])^(a[344] & b[325])^(a[343] & b[326])^(a[342] & b[327])^(a[341] & b[328])^(a[340] & b[329])^(a[339] & b[330])^(a[338] & b[331])^(a[337] & b[332])^(a[336] & b[333])^(a[335] & b[334])^(a[334] & b[335])^(a[333] & b[336])^(a[332] & b[337])^(a[331] & b[338])^(a[330] & b[339])^(a[329] & b[340])^(a[328] & b[341])^(a[327] & b[342])^(a[326] & b[343])^(a[325] & b[344])^(a[324] & b[345])^(a[323] & b[346])^(a[322] & b[347])^(a[321] & b[348])^(a[320] & b[349])^(a[319] & b[350])^(a[318] & b[351])^(a[317] & b[352])^(a[316] & b[353])^(a[315] & b[354])^(a[314] & b[355])^(a[313] & b[356])^(a[312] & b[357])^(a[311] & b[358])^(a[310] & b[359])^(a[309] & b[360])^(a[308] & b[361])^(a[307] & b[362])^(a[306] & b[363])^(a[305] & b[364])^(a[304] & b[365])^(a[303] & b[366])^(a[302] & b[367])^(a[301] & b[368])^(a[300] & b[369])^(a[299] & b[370])^(a[298] & b[371])^(a[297] & b[372])^(a[296] & b[373])^(a[295] & b[374])^(a[294] & b[375])^(a[293] & b[376])^(a[292] & b[377])^(a[291] & b[378])^(a[290] & b[379])^(a[289] & b[380])^(a[288] & b[381])^(a[287] & b[382])^(a[286] & b[383])^(a[285] & b[384])^(a[284] & b[385])^(a[283] & b[386])^(a[282] & b[387])^(a[281] & b[388])^(a[280] & b[389])^(a[279] & b[390])^(a[278] & b[391])^(a[277] & b[392])^(a[276] & b[393])^(a[275] & b[394])^(a[274] & b[395])^(a[273] & b[396])^(a[272] & b[397])^(a[271] & b[398])^(a[270] & b[399])^(a[269] & b[400])^(a[268] & b[401])^(a[267] & b[402])^(a[266] & b[403])^(a[265] & b[404])^(a[264] & b[405])^(a[263] & b[406])^(a[262] & b[407])^(a[261] & b[408]);
assign y[670] = (a[408] & b[262])^(a[407] & b[263])^(a[406] & b[264])^(a[405] & b[265])^(a[404] & b[266])^(a[403] & b[267])^(a[402] & b[268])^(a[401] & b[269])^(a[400] & b[270])^(a[399] & b[271])^(a[398] & b[272])^(a[397] & b[273])^(a[396] & b[274])^(a[395] & b[275])^(a[394] & b[276])^(a[393] & b[277])^(a[392] & b[278])^(a[391] & b[279])^(a[390] & b[280])^(a[389] & b[281])^(a[388] & b[282])^(a[387] & b[283])^(a[386] & b[284])^(a[385] & b[285])^(a[384] & b[286])^(a[383] & b[287])^(a[382] & b[288])^(a[381] & b[289])^(a[380] & b[290])^(a[379] & b[291])^(a[378] & b[292])^(a[377] & b[293])^(a[376] & b[294])^(a[375] & b[295])^(a[374] & b[296])^(a[373] & b[297])^(a[372] & b[298])^(a[371] & b[299])^(a[370] & b[300])^(a[369] & b[301])^(a[368] & b[302])^(a[367] & b[303])^(a[366] & b[304])^(a[365] & b[305])^(a[364] & b[306])^(a[363] & b[307])^(a[362] & b[308])^(a[361] & b[309])^(a[360] & b[310])^(a[359] & b[311])^(a[358] & b[312])^(a[357] & b[313])^(a[356] & b[314])^(a[355] & b[315])^(a[354] & b[316])^(a[353] & b[317])^(a[352] & b[318])^(a[351] & b[319])^(a[350] & b[320])^(a[349] & b[321])^(a[348] & b[322])^(a[347] & b[323])^(a[346] & b[324])^(a[345] & b[325])^(a[344] & b[326])^(a[343] & b[327])^(a[342] & b[328])^(a[341] & b[329])^(a[340] & b[330])^(a[339] & b[331])^(a[338] & b[332])^(a[337] & b[333])^(a[336] & b[334])^(a[335] & b[335])^(a[334] & b[336])^(a[333] & b[337])^(a[332] & b[338])^(a[331] & b[339])^(a[330] & b[340])^(a[329] & b[341])^(a[328] & b[342])^(a[327] & b[343])^(a[326] & b[344])^(a[325] & b[345])^(a[324] & b[346])^(a[323] & b[347])^(a[322] & b[348])^(a[321] & b[349])^(a[320] & b[350])^(a[319] & b[351])^(a[318] & b[352])^(a[317] & b[353])^(a[316] & b[354])^(a[315] & b[355])^(a[314] & b[356])^(a[313] & b[357])^(a[312] & b[358])^(a[311] & b[359])^(a[310] & b[360])^(a[309] & b[361])^(a[308] & b[362])^(a[307] & b[363])^(a[306] & b[364])^(a[305] & b[365])^(a[304] & b[366])^(a[303] & b[367])^(a[302] & b[368])^(a[301] & b[369])^(a[300] & b[370])^(a[299] & b[371])^(a[298] & b[372])^(a[297] & b[373])^(a[296] & b[374])^(a[295] & b[375])^(a[294] & b[376])^(a[293] & b[377])^(a[292] & b[378])^(a[291] & b[379])^(a[290] & b[380])^(a[289] & b[381])^(a[288] & b[382])^(a[287] & b[383])^(a[286] & b[384])^(a[285] & b[385])^(a[284] & b[386])^(a[283] & b[387])^(a[282] & b[388])^(a[281] & b[389])^(a[280] & b[390])^(a[279] & b[391])^(a[278] & b[392])^(a[277] & b[393])^(a[276] & b[394])^(a[275] & b[395])^(a[274] & b[396])^(a[273] & b[397])^(a[272] & b[398])^(a[271] & b[399])^(a[270] & b[400])^(a[269] & b[401])^(a[268] & b[402])^(a[267] & b[403])^(a[266] & b[404])^(a[265] & b[405])^(a[264] & b[406])^(a[263] & b[407])^(a[262] & b[408]);
assign y[671] = (a[408] & b[263])^(a[407] & b[264])^(a[406] & b[265])^(a[405] & b[266])^(a[404] & b[267])^(a[403] & b[268])^(a[402] & b[269])^(a[401] & b[270])^(a[400] & b[271])^(a[399] & b[272])^(a[398] & b[273])^(a[397] & b[274])^(a[396] & b[275])^(a[395] & b[276])^(a[394] & b[277])^(a[393] & b[278])^(a[392] & b[279])^(a[391] & b[280])^(a[390] & b[281])^(a[389] & b[282])^(a[388] & b[283])^(a[387] & b[284])^(a[386] & b[285])^(a[385] & b[286])^(a[384] & b[287])^(a[383] & b[288])^(a[382] & b[289])^(a[381] & b[290])^(a[380] & b[291])^(a[379] & b[292])^(a[378] & b[293])^(a[377] & b[294])^(a[376] & b[295])^(a[375] & b[296])^(a[374] & b[297])^(a[373] & b[298])^(a[372] & b[299])^(a[371] & b[300])^(a[370] & b[301])^(a[369] & b[302])^(a[368] & b[303])^(a[367] & b[304])^(a[366] & b[305])^(a[365] & b[306])^(a[364] & b[307])^(a[363] & b[308])^(a[362] & b[309])^(a[361] & b[310])^(a[360] & b[311])^(a[359] & b[312])^(a[358] & b[313])^(a[357] & b[314])^(a[356] & b[315])^(a[355] & b[316])^(a[354] & b[317])^(a[353] & b[318])^(a[352] & b[319])^(a[351] & b[320])^(a[350] & b[321])^(a[349] & b[322])^(a[348] & b[323])^(a[347] & b[324])^(a[346] & b[325])^(a[345] & b[326])^(a[344] & b[327])^(a[343] & b[328])^(a[342] & b[329])^(a[341] & b[330])^(a[340] & b[331])^(a[339] & b[332])^(a[338] & b[333])^(a[337] & b[334])^(a[336] & b[335])^(a[335] & b[336])^(a[334] & b[337])^(a[333] & b[338])^(a[332] & b[339])^(a[331] & b[340])^(a[330] & b[341])^(a[329] & b[342])^(a[328] & b[343])^(a[327] & b[344])^(a[326] & b[345])^(a[325] & b[346])^(a[324] & b[347])^(a[323] & b[348])^(a[322] & b[349])^(a[321] & b[350])^(a[320] & b[351])^(a[319] & b[352])^(a[318] & b[353])^(a[317] & b[354])^(a[316] & b[355])^(a[315] & b[356])^(a[314] & b[357])^(a[313] & b[358])^(a[312] & b[359])^(a[311] & b[360])^(a[310] & b[361])^(a[309] & b[362])^(a[308] & b[363])^(a[307] & b[364])^(a[306] & b[365])^(a[305] & b[366])^(a[304] & b[367])^(a[303] & b[368])^(a[302] & b[369])^(a[301] & b[370])^(a[300] & b[371])^(a[299] & b[372])^(a[298] & b[373])^(a[297] & b[374])^(a[296] & b[375])^(a[295] & b[376])^(a[294] & b[377])^(a[293] & b[378])^(a[292] & b[379])^(a[291] & b[380])^(a[290] & b[381])^(a[289] & b[382])^(a[288] & b[383])^(a[287] & b[384])^(a[286] & b[385])^(a[285] & b[386])^(a[284] & b[387])^(a[283] & b[388])^(a[282] & b[389])^(a[281] & b[390])^(a[280] & b[391])^(a[279] & b[392])^(a[278] & b[393])^(a[277] & b[394])^(a[276] & b[395])^(a[275] & b[396])^(a[274] & b[397])^(a[273] & b[398])^(a[272] & b[399])^(a[271] & b[400])^(a[270] & b[401])^(a[269] & b[402])^(a[268] & b[403])^(a[267] & b[404])^(a[266] & b[405])^(a[265] & b[406])^(a[264] & b[407])^(a[263] & b[408]);
assign y[672] = (a[408] & b[264])^(a[407] & b[265])^(a[406] & b[266])^(a[405] & b[267])^(a[404] & b[268])^(a[403] & b[269])^(a[402] & b[270])^(a[401] & b[271])^(a[400] & b[272])^(a[399] & b[273])^(a[398] & b[274])^(a[397] & b[275])^(a[396] & b[276])^(a[395] & b[277])^(a[394] & b[278])^(a[393] & b[279])^(a[392] & b[280])^(a[391] & b[281])^(a[390] & b[282])^(a[389] & b[283])^(a[388] & b[284])^(a[387] & b[285])^(a[386] & b[286])^(a[385] & b[287])^(a[384] & b[288])^(a[383] & b[289])^(a[382] & b[290])^(a[381] & b[291])^(a[380] & b[292])^(a[379] & b[293])^(a[378] & b[294])^(a[377] & b[295])^(a[376] & b[296])^(a[375] & b[297])^(a[374] & b[298])^(a[373] & b[299])^(a[372] & b[300])^(a[371] & b[301])^(a[370] & b[302])^(a[369] & b[303])^(a[368] & b[304])^(a[367] & b[305])^(a[366] & b[306])^(a[365] & b[307])^(a[364] & b[308])^(a[363] & b[309])^(a[362] & b[310])^(a[361] & b[311])^(a[360] & b[312])^(a[359] & b[313])^(a[358] & b[314])^(a[357] & b[315])^(a[356] & b[316])^(a[355] & b[317])^(a[354] & b[318])^(a[353] & b[319])^(a[352] & b[320])^(a[351] & b[321])^(a[350] & b[322])^(a[349] & b[323])^(a[348] & b[324])^(a[347] & b[325])^(a[346] & b[326])^(a[345] & b[327])^(a[344] & b[328])^(a[343] & b[329])^(a[342] & b[330])^(a[341] & b[331])^(a[340] & b[332])^(a[339] & b[333])^(a[338] & b[334])^(a[337] & b[335])^(a[336] & b[336])^(a[335] & b[337])^(a[334] & b[338])^(a[333] & b[339])^(a[332] & b[340])^(a[331] & b[341])^(a[330] & b[342])^(a[329] & b[343])^(a[328] & b[344])^(a[327] & b[345])^(a[326] & b[346])^(a[325] & b[347])^(a[324] & b[348])^(a[323] & b[349])^(a[322] & b[350])^(a[321] & b[351])^(a[320] & b[352])^(a[319] & b[353])^(a[318] & b[354])^(a[317] & b[355])^(a[316] & b[356])^(a[315] & b[357])^(a[314] & b[358])^(a[313] & b[359])^(a[312] & b[360])^(a[311] & b[361])^(a[310] & b[362])^(a[309] & b[363])^(a[308] & b[364])^(a[307] & b[365])^(a[306] & b[366])^(a[305] & b[367])^(a[304] & b[368])^(a[303] & b[369])^(a[302] & b[370])^(a[301] & b[371])^(a[300] & b[372])^(a[299] & b[373])^(a[298] & b[374])^(a[297] & b[375])^(a[296] & b[376])^(a[295] & b[377])^(a[294] & b[378])^(a[293] & b[379])^(a[292] & b[380])^(a[291] & b[381])^(a[290] & b[382])^(a[289] & b[383])^(a[288] & b[384])^(a[287] & b[385])^(a[286] & b[386])^(a[285] & b[387])^(a[284] & b[388])^(a[283] & b[389])^(a[282] & b[390])^(a[281] & b[391])^(a[280] & b[392])^(a[279] & b[393])^(a[278] & b[394])^(a[277] & b[395])^(a[276] & b[396])^(a[275] & b[397])^(a[274] & b[398])^(a[273] & b[399])^(a[272] & b[400])^(a[271] & b[401])^(a[270] & b[402])^(a[269] & b[403])^(a[268] & b[404])^(a[267] & b[405])^(a[266] & b[406])^(a[265] & b[407])^(a[264] & b[408]);
assign y[673] = (a[408] & b[265])^(a[407] & b[266])^(a[406] & b[267])^(a[405] & b[268])^(a[404] & b[269])^(a[403] & b[270])^(a[402] & b[271])^(a[401] & b[272])^(a[400] & b[273])^(a[399] & b[274])^(a[398] & b[275])^(a[397] & b[276])^(a[396] & b[277])^(a[395] & b[278])^(a[394] & b[279])^(a[393] & b[280])^(a[392] & b[281])^(a[391] & b[282])^(a[390] & b[283])^(a[389] & b[284])^(a[388] & b[285])^(a[387] & b[286])^(a[386] & b[287])^(a[385] & b[288])^(a[384] & b[289])^(a[383] & b[290])^(a[382] & b[291])^(a[381] & b[292])^(a[380] & b[293])^(a[379] & b[294])^(a[378] & b[295])^(a[377] & b[296])^(a[376] & b[297])^(a[375] & b[298])^(a[374] & b[299])^(a[373] & b[300])^(a[372] & b[301])^(a[371] & b[302])^(a[370] & b[303])^(a[369] & b[304])^(a[368] & b[305])^(a[367] & b[306])^(a[366] & b[307])^(a[365] & b[308])^(a[364] & b[309])^(a[363] & b[310])^(a[362] & b[311])^(a[361] & b[312])^(a[360] & b[313])^(a[359] & b[314])^(a[358] & b[315])^(a[357] & b[316])^(a[356] & b[317])^(a[355] & b[318])^(a[354] & b[319])^(a[353] & b[320])^(a[352] & b[321])^(a[351] & b[322])^(a[350] & b[323])^(a[349] & b[324])^(a[348] & b[325])^(a[347] & b[326])^(a[346] & b[327])^(a[345] & b[328])^(a[344] & b[329])^(a[343] & b[330])^(a[342] & b[331])^(a[341] & b[332])^(a[340] & b[333])^(a[339] & b[334])^(a[338] & b[335])^(a[337] & b[336])^(a[336] & b[337])^(a[335] & b[338])^(a[334] & b[339])^(a[333] & b[340])^(a[332] & b[341])^(a[331] & b[342])^(a[330] & b[343])^(a[329] & b[344])^(a[328] & b[345])^(a[327] & b[346])^(a[326] & b[347])^(a[325] & b[348])^(a[324] & b[349])^(a[323] & b[350])^(a[322] & b[351])^(a[321] & b[352])^(a[320] & b[353])^(a[319] & b[354])^(a[318] & b[355])^(a[317] & b[356])^(a[316] & b[357])^(a[315] & b[358])^(a[314] & b[359])^(a[313] & b[360])^(a[312] & b[361])^(a[311] & b[362])^(a[310] & b[363])^(a[309] & b[364])^(a[308] & b[365])^(a[307] & b[366])^(a[306] & b[367])^(a[305] & b[368])^(a[304] & b[369])^(a[303] & b[370])^(a[302] & b[371])^(a[301] & b[372])^(a[300] & b[373])^(a[299] & b[374])^(a[298] & b[375])^(a[297] & b[376])^(a[296] & b[377])^(a[295] & b[378])^(a[294] & b[379])^(a[293] & b[380])^(a[292] & b[381])^(a[291] & b[382])^(a[290] & b[383])^(a[289] & b[384])^(a[288] & b[385])^(a[287] & b[386])^(a[286] & b[387])^(a[285] & b[388])^(a[284] & b[389])^(a[283] & b[390])^(a[282] & b[391])^(a[281] & b[392])^(a[280] & b[393])^(a[279] & b[394])^(a[278] & b[395])^(a[277] & b[396])^(a[276] & b[397])^(a[275] & b[398])^(a[274] & b[399])^(a[273] & b[400])^(a[272] & b[401])^(a[271] & b[402])^(a[270] & b[403])^(a[269] & b[404])^(a[268] & b[405])^(a[267] & b[406])^(a[266] & b[407])^(a[265] & b[408]);
assign y[674] = (a[408] & b[266])^(a[407] & b[267])^(a[406] & b[268])^(a[405] & b[269])^(a[404] & b[270])^(a[403] & b[271])^(a[402] & b[272])^(a[401] & b[273])^(a[400] & b[274])^(a[399] & b[275])^(a[398] & b[276])^(a[397] & b[277])^(a[396] & b[278])^(a[395] & b[279])^(a[394] & b[280])^(a[393] & b[281])^(a[392] & b[282])^(a[391] & b[283])^(a[390] & b[284])^(a[389] & b[285])^(a[388] & b[286])^(a[387] & b[287])^(a[386] & b[288])^(a[385] & b[289])^(a[384] & b[290])^(a[383] & b[291])^(a[382] & b[292])^(a[381] & b[293])^(a[380] & b[294])^(a[379] & b[295])^(a[378] & b[296])^(a[377] & b[297])^(a[376] & b[298])^(a[375] & b[299])^(a[374] & b[300])^(a[373] & b[301])^(a[372] & b[302])^(a[371] & b[303])^(a[370] & b[304])^(a[369] & b[305])^(a[368] & b[306])^(a[367] & b[307])^(a[366] & b[308])^(a[365] & b[309])^(a[364] & b[310])^(a[363] & b[311])^(a[362] & b[312])^(a[361] & b[313])^(a[360] & b[314])^(a[359] & b[315])^(a[358] & b[316])^(a[357] & b[317])^(a[356] & b[318])^(a[355] & b[319])^(a[354] & b[320])^(a[353] & b[321])^(a[352] & b[322])^(a[351] & b[323])^(a[350] & b[324])^(a[349] & b[325])^(a[348] & b[326])^(a[347] & b[327])^(a[346] & b[328])^(a[345] & b[329])^(a[344] & b[330])^(a[343] & b[331])^(a[342] & b[332])^(a[341] & b[333])^(a[340] & b[334])^(a[339] & b[335])^(a[338] & b[336])^(a[337] & b[337])^(a[336] & b[338])^(a[335] & b[339])^(a[334] & b[340])^(a[333] & b[341])^(a[332] & b[342])^(a[331] & b[343])^(a[330] & b[344])^(a[329] & b[345])^(a[328] & b[346])^(a[327] & b[347])^(a[326] & b[348])^(a[325] & b[349])^(a[324] & b[350])^(a[323] & b[351])^(a[322] & b[352])^(a[321] & b[353])^(a[320] & b[354])^(a[319] & b[355])^(a[318] & b[356])^(a[317] & b[357])^(a[316] & b[358])^(a[315] & b[359])^(a[314] & b[360])^(a[313] & b[361])^(a[312] & b[362])^(a[311] & b[363])^(a[310] & b[364])^(a[309] & b[365])^(a[308] & b[366])^(a[307] & b[367])^(a[306] & b[368])^(a[305] & b[369])^(a[304] & b[370])^(a[303] & b[371])^(a[302] & b[372])^(a[301] & b[373])^(a[300] & b[374])^(a[299] & b[375])^(a[298] & b[376])^(a[297] & b[377])^(a[296] & b[378])^(a[295] & b[379])^(a[294] & b[380])^(a[293] & b[381])^(a[292] & b[382])^(a[291] & b[383])^(a[290] & b[384])^(a[289] & b[385])^(a[288] & b[386])^(a[287] & b[387])^(a[286] & b[388])^(a[285] & b[389])^(a[284] & b[390])^(a[283] & b[391])^(a[282] & b[392])^(a[281] & b[393])^(a[280] & b[394])^(a[279] & b[395])^(a[278] & b[396])^(a[277] & b[397])^(a[276] & b[398])^(a[275] & b[399])^(a[274] & b[400])^(a[273] & b[401])^(a[272] & b[402])^(a[271] & b[403])^(a[270] & b[404])^(a[269] & b[405])^(a[268] & b[406])^(a[267] & b[407])^(a[266] & b[408]);
assign y[675] = (a[408] & b[267])^(a[407] & b[268])^(a[406] & b[269])^(a[405] & b[270])^(a[404] & b[271])^(a[403] & b[272])^(a[402] & b[273])^(a[401] & b[274])^(a[400] & b[275])^(a[399] & b[276])^(a[398] & b[277])^(a[397] & b[278])^(a[396] & b[279])^(a[395] & b[280])^(a[394] & b[281])^(a[393] & b[282])^(a[392] & b[283])^(a[391] & b[284])^(a[390] & b[285])^(a[389] & b[286])^(a[388] & b[287])^(a[387] & b[288])^(a[386] & b[289])^(a[385] & b[290])^(a[384] & b[291])^(a[383] & b[292])^(a[382] & b[293])^(a[381] & b[294])^(a[380] & b[295])^(a[379] & b[296])^(a[378] & b[297])^(a[377] & b[298])^(a[376] & b[299])^(a[375] & b[300])^(a[374] & b[301])^(a[373] & b[302])^(a[372] & b[303])^(a[371] & b[304])^(a[370] & b[305])^(a[369] & b[306])^(a[368] & b[307])^(a[367] & b[308])^(a[366] & b[309])^(a[365] & b[310])^(a[364] & b[311])^(a[363] & b[312])^(a[362] & b[313])^(a[361] & b[314])^(a[360] & b[315])^(a[359] & b[316])^(a[358] & b[317])^(a[357] & b[318])^(a[356] & b[319])^(a[355] & b[320])^(a[354] & b[321])^(a[353] & b[322])^(a[352] & b[323])^(a[351] & b[324])^(a[350] & b[325])^(a[349] & b[326])^(a[348] & b[327])^(a[347] & b[328])^(a[346] & b[329])^(a[345] & b[330])^(a[344] & b[331])^(a[343] & b[332])^(a[342] & b[333])^(a[341] & b[334])^(a[340] & b[335])^(a[339] & b[336])^(a[338] & b[337])^(a[337] & b[338])^(a[336] & b[339])^(a[335] & b[340])^(a[334] & b[341])^(a[333] & b[342])^(a[332] & b[343])^(a[331] & b[344])^(a[330] & b[345])^(a[329] & b[346])^(a[328] & b[347])^(a[327] & b[348])^(a[326] & b[349])^(a[325] & b[350])^(a[324] & b[351])^(a[323] & b[352])^(a[322] & b[353])^(a[321] & b[354])^(a[320] & b[355])^(a[319] & b[356])^(a[318] & b[357])^(a[317] & b[358])^(a[316] & b[359])^(a[315] & b[360])^(a[314] & b[361])^(a[313] & b[362])^(a[312] & b[363])^(a[311] & b[364])^(a[310] & b[365])^(a[309] & b[366])^(a[308] & b[367])^(a[307] & b[368])^(a[306] & b[369])^(a[305] & b[370])^(a[304] & b[371])^(a[303] & b[372])^(a[302] & b[373])^(a[301] & b[374])^(a[300] & b[375])^(a[299] & b[376])^(a[298] & b[377])^(a[297] & b[378])^(a[296] & b[379])^(a[295] & b[380])^(a[294] & b[381])^(a[293] & b[382])^(a[292] & b[383])^(a[291] & b[384])^(a[290] & b[385])^(a[289] & b[386])^(a[288] & b[387])^(a[287] & b[388])^(a[286] & b[389])^(a[285] & b[390])^(a[284] & b[391])^(a[283] & b[392])^(a[282] & b[393])^(a[281] & b[394])^(a[280] & b[395])^(a[279] & b[396])^(a[278] & b[397])^(a[277] & b[398])^(a[276] & b[399])^(a[275] & b[400])^(a[274] & b[401])^(a[273] & b[402])^(a[272] & b[403])^(a[271] & b[404])^(a[270] & b[405])^(a[269] & b[406])^(a[268] & b[407])^(a[267] & b[408]);
assign y[676] = (a[408] & b[268])^(a[407] & b[269])^(a[406] & b[270])^(a[405] & b[271])^(a[404] & b[272])^(a[403] & b[273])^(a[402] & b[274])^(a[401] & b[275])^(a[400] & b[276])^(a[399] & b[277])^(a[398] & b[278])^(a[397] & b[279])^(a[396] & b[280])^(a[395] & b[281])^(a[394] & b[282])^(a[393] & b[283])^(a[392] & b[284])^(a[391] & b[285])^(a[390] & b[286])^(a[389] & b[287])^(a[388] & b[288])^(a[387] & b[289])^(a[386] & b[290])^(a[385] & b[291])^(a[384] & b[292])^(a[383] & b[293])^(a[382] & b[294])^(a[381] & b[295])^(a[380] & b[296])^(a[379] & b[297])^(a[378] & b[298])^(a[377] & b[299])^(a[376] & b[300])^(a[375] & b[301])^(a[374] & b[302])^(a[373] & b[303])^(a[372] & b[304])^(a[371] & b[305])^(a[370] & b[306])^(a[369] & b[307])^(a[368] & b[308])^(a[367] & b[309])^(a[366] & b[310])^(a[365] & b[311])^(a[364] & b[312])^(a[363] & b[313])^(a[362] & b[314])^(a[361] & b[315])^(a[360] & b[316])^(a[359] & b[317])^(a[358] & b[318])^(a[357] & b[319])^(a[356] & b[320])^(a[355] & b[321])^(a[354] & b[322])^(a[353] & b[323])^(a[352] & b[324])^(a[351] & b[325])^(a[350] & b[326])^(a[349] & b[327])^(a[348] & b[328])^(a[347] & b[329])^(a[346] & b[330])^(a[345] & b[331])^(a[344] & b[332])^(a[343] & b[333])^(a[342] & b[334])^(a[341] & b[335])^(a[340] & b[336])^(a[339] & b[337])^(a[338] & b[338])^(a[337] & b[339])^(a[336] & b[340])^(a[335] & b[341])^(a[334] & b[342])^(a[333] & b[343])^(a[332] & b[344])^(a[331] & b[345])^(a[330] & b[346])^(a[329] & b[347])^(a[328] & b[348])^(a[327] & b[349])^(a[326] & b[350])^(a[325] & b[351])^(a[324] & b[352])^(a[323] & b[353])^(a[322] & b[354])^(a[321] & b[355])^(a[320] & b[356])^(a[319] & b[357])^(a[318] & b[358])^(a[317] & b[359])^(a[316] & b[360])^(a[315] & b[361])^(a[314] & b[362])^(a[313] & b[363])^(a[312] & b[364])^(a[311] & b[365])^(a[310] & b[366])^(a[309] & b[367])^(a[308] & b[368])^(a[307] & b[369])^(a[306] & b[370])^(a[305] & b[371])^(a[304] & b[372])^(a[303] & b[373])^(a[302] & b[374])^(a[301] & b[375])^(a[300] & b[376])^(a[299] & b[377])^(a[298] & b[378])^(a[297] & b[379])^(a[296] & b[380])^(a[295] & b[381])^(a[294] & b[382])^(a[293] & b[383])^(a[292] & b[384])^(a[291] & b[385])^(a[290] & b[386])^(a[289] & b[387])^(a[288] & b[388])^(a[287] & b[389])^(a[286] & b[390])^(a[285] & b[391])^(a[284] & b[392])^(a[283] & b[393])^(a[282] & b[394])^(a[281] & b[395])^(a[280] & b[396])^(a[279] & b[397])^(a[278] & b[398])^(a[277] & b[399])^(a[276] & b[400])^(a[275] & b[401])^(a[274] & b[402])^(a[273] & b[403])^(a[272] & b[404])^(a[271] & b[405])^(a[270] & b[406])^(a[269] & b[407])^(a[268] & b[408]);
assign y[677] = (a[408] & b[269])^(a[407] & b[270])^(a[406] & b[271])^(a[405] & b[272])^(a[404] & b[273])^(a[403] & b[274])^(a[402] & b[275])^(a[401] & b[276])^(a[400] & b[277])^(a[399] & b[278])^(a[398] & b[279])^(a[397] & b[280])^(a[396] & b[281])^(a[395] & b[282])^(a[394] & b[283])^(a[393] & b[284])^(a[392] & b[285])^(a[391] & b[286])^(a[390] & b[287])^(a[389] & b[288])^(a[388] & b[289])^(a[387] & b[290])^(a[386] & b[291])^(a[385] & b[292])^(a[384] & b[293])^(a[383] & b[294])^(a[382] & b[295])^(a[381] & b[296])^(a[380] & b[297])^(a[379] & b[298])^(a[378] & b[299])^(a[377] & b[300])^(a[376] & b[301])^(a[375] & b[302])^(a[374] & b[303])^(a[373] & b[304])^(a[372] & b[305])^(a[371] & b[306])^(a[370] & b[307])^(a[369] & b[308])^(a[368] & b[309])^(a[367] & b[310])^(a[366] & b[311])^(a[365] & b[312])^(a[364] & b[313])^(a[363] & b[314])^(a[362] & b[315])^(a[361] & b[316])^(a[360] & b[317])^(a[359] & b[318])^(a[358] & b[319])^(a[357] & b[320])^(a[356] & b[321])^(a[355] & b[322])^(a[354] & b[323])^(a[353] & b[324])^(a[352] & b[325])^(a[351] & b[326])^(a[350] & b[327])^(a[349] & b[328])^(a[348] & b[329])^(a[347] & b[330])^(a[346] & b[331])^(a[345] & b[332])^(a[344] & b[333])^(a[343] & b[334])^(a[342] & b[335])^(a[341] & b[336])^(a[340] & b[337])^(a[339] & b[338])^(a[338] & b[339])^(a[337] & b[340])^(a[336] & b[341])^(a[335] & b[342])^(a[334] & b[343])^(a[333] & b[344])^(a[332] & b[345])^(a[331] & b[346])^(a[330] & b[347])^(a[329] & b[348])^(a[328] & b[349])^(a[327] & b[350])^(a[326] & b[351])^(a[325] & b[352])^(a[324] & b[353])^(a[323] & b[354])^(a[322] & b[355])^(a[321] & b[356])^(a[320] & b[357])^(a[319] & b[358])^(a[318] & b[359])^(a[317] & b[360])^(a[316] & b[361])^(a[315] & b[362])^(a[314] & b[363])^(a[313] & b[364])^(a[312] & b[365])^(a[311] & b[366])^(a[310] & b[367])^(a[309] & b[368])^(a[308] & b[369])^(a[307] & b[370])^(a[306] & b[371])^(a[305] & b[372])^(a[304] & b[373])^(a[303] & b[374])^(a[302] & b[375])^(a[301] & b[376])^(a[300] & b[377])^(a[299] & b[378])^(a[298] & b[379])^(a[297] & b[380])^(a[296] & b[381])^(a[295] & b[382])^(a[294] & b[383])^(a[293] & b[384])^(a[292] & b[385])^(a[291] & b[386])^(a[290] & b[387])^(a[289] & b[388])^(a[288] & b[389])^(a[287] & b[390])^(a[286] & b[391])^(a[285] & b[392])^(a[284] & b[393])^(a[283] & b[394])^(a[282] & b[395])^(a[281] & b[396])^(a[280] & b[397])^(a[279] & b[398])^(a[278] & b[399])^(a[277] & b[400])^(a[276] & b[401])^(a[275] & b[402])^(a[274] & b[403])^(a[273] & b[404])^(a[272] & b[405])^(a[271] & b[406])^(a[270] & b[407])^(a[269] & b[408]);
assign y[678] = (a[408] & b[270])^(a[407] & b[271])^(a[406] & b[272])^(a[405] & b[273])^(a[404] & b[274])^(a[403] & b[275])^(a[402] & b[276])^(a[401] & b[277])^(a[400] & b[278])^(a[399] & b[279])^(a[398] & b[280])^(a[397] & b[281])^(a[396] & b[282])^(a[395] & b[283])^(a[394] & b[284])^(a[393] & b[285])^(a[392] & b[286])^(a[391] & b[287])^(a[390] & b[288])^(a[389] & b[289])^(a[388] & b[290])^(a[387] & b[291])^(a[386] & b[292])^(a[385] & b[293])^(a[384] & b[294])^(a[383] & b[295])^(a[382] & b[296])^(a[381] & b[297])^(a[380] & b[298])^(a[379] & b[299])^(a[378] & b[300])^(a[377] & b[301])^(a[376] & b[302])^(a[375] & b[303])^(a[374] & b[304])^(a[373] & b[305])^(a[372] & b[306])^(a[371] & b[307])^(a[370] & b[308])^(a[369] & b[309])^(a[368] & b[310])^(a[367] & b[311])^(a[366] & b[312])^(a[365] & b[313])^(a[364] & b[314])^(a[363] & b[315])^(a[362] & b[316])^(a[361] & b[317])^(a[360] & b[318])^(a[359] & b[319])^(a[358] & b[320])^(a[357] & b[321])^(a[356] & b[322])^(a[355] & b[323])^(a[354] & b[324])^(a[353] & b[325])^(a[352] & b[326])^(a[351] & b[327])^(a[350] & b[328])^(a[349] & b[329])^(a[348] & b[330])^(a[347] & b[331])^(a[346] & b[332])^(a[345] & b[333])^(a[344] & b[334])^(a[343] & b[335])^(a[342] & b[336])^(a[341] & b[337])^(a[340] & b[338])^(a[339] & b[339])^(a[338] & b[340])^(a[337] & b[341])^(a[336] & b[342])^(a[335] & b[343])^(a[334] & b[344])^(a[333] & b[345])^(a[332] & b[346])^(a[331] & b[347])^(a[330] & b[348])^(a[329] & b[349])^(a[328] & b[350])^(a[327] & b[351])^(a[326] & b[352])^(a[325] & b[353])^(a[324] & b[354])^(a[323] & b[355])^(a[322] & b[356])^(a[321] & b[357])^(a[320] & b[358])^(a[319] & b[359])^(a[318] & b[360])^(a[317] & b[361])^(a[316] & b[362])^(a[315] & b[363])^(a[314] & b[364])^(a[313] & b[365])^(a[312] & b[366])^(a[311] & b[367])^(a[310] & b[368])^(a[309] & b[369])^(a[308] & b[370])^(a[307] & b[371])^(a[306] & b[372])^(a[305] & b[373])^(a[304] & b[374])^(a[303] & b[375])^(a[302] & b[376])^(a[301] & b[377])^(a[300] & b[378])^(a[299] & b[379])^(a[298] & b[380])^(a[297] & b[381])^(a[296] & b[382])^(a[295] & b[383])^(a[294] & b[384])^(a[293] & b[385])^(a[292] & b[386])^(a[291] & b[387])^(a[290] & b[388])^(a[289] & b[389])^(a[288] & b[390])^(a[287] & b[391])^(a[286] & b[392])^(a[285] & b[393])^(a[284] & b[394])^(a[283] & b[395])^(a[282] & b[396])^(a[281] & b[397])^(a[280] & b[398])^(a[279] & b[399])^(a[278] & b[400])^(a[277] & b[401])^(a[276] & b[402])^(a[275] & b[403])^(a[274] & b[404])^(a[273] & b[405])^(a[272] & b[406])^(a[271] & b[407])^(a[270] & b[408]);
assign y[679] = (a[408] & b[271])^(a[407] & b[272])^(a[406] & b[273])^(a[405] & b[274])^(a[404] & b[275])^(a[403] & b[276])^(a[402] & b[277])^(a[401] & b[278])^(a[400] & b[279])^(a[399] & b[280])^(a[398] & b[281])^(a[397] & b[282])^(a[396] & b[283])^(a[395] & b[284])^(a[394] & b[285])^(a[393] & b[286])^(a[392] & b[287])^(a[391] & b[288])^(a[390] & b[289])^(a[389] & b[290])^(a[388] & b[291])^(a[387] & b[292])^(a[386] & b[293])^(a[385] & b[294])^(a[384] & b[295])^(a[383] & b[296])^(a[382] & b[297])^(a[381] & b[298])^(a[380] & b[299])^(a[379] & b[300])^(a[378] & b[301])^(a[377] & b[302])^(a[376] & b[303])^(a[375] & b[304])^(a[374] & b[305])^(a[373] & b[306])^(a[372] & b[307])^(a[371] & b[308])^(a[370] & b[309])^(a[369] & b[310])^(a[368] & b[311])^(a[367] & b[312])^(a[366] & b[313])^(a[365] & b[314])^(a[364] & b[315])^(a[363] & b[316])^(a[362] & b[317])^(a[361] & b[318])^(a[360] & b[319])^(a[359] & b[320])^(a[358] & b[321])^(a[357] & b[322])^(a[356] & b[323])^(a[355] & b[324])^(a[354] & b[325])^(a[353] & b[326])^(a[352] & b[327])^(a[351] & b[328])^(a[350] & b[329])^(a[349] & b[330])^(a[348] & b[331])^(a[347] & b[332])^(a[346] & b[333])^(a[345] & b[334])^(a[344] & b[335])^(a[343] & b[336])^(a[342] & b[337])^(a[341] & b[338])^(a[340] & b[339])^(a[339] & b[340])^(a[338] & b[341])^(a[337] & b[342])^(a[336] & b[343])^(a[335] & b[344])^(a[334] & b[345])^(a[333] & b[346])^(a[332] & b[347])^(a[331] & b[348])^(a[330] & b[349])^(a[329] & b[350])^(a[328] & b[351])^(a[327] & b[352])^(a[326] & b[353])^(a[325] & b[354])^(a[324] & b[355])^(a[323] & b[356])^(a[322] & b[357])^(a[321] & b[358])^(a[320] & b[359])^(a[319] & b[360])^(a[318] & b[361])^(a[317] & b[362])^(a[316] & b[363])^(a[315] & b[364])^(a[314] & b[365])^(a[313] & b[366])^(a[312] & b[367])^(a[311] & b[368])^(a[310] & b[369])^(a[309] & b[370])^(a[308] & b[371])^(a[307] & b[372])^(a[306] & b[373])^(a[305] & b[374])^(a[304] & b[375])^(a[303] & b[376])^(a[302] & b[377])^(a[301] & b[378])^(a[300] & b[379])^(a[299] & b[380])^(a[298] & b[381])^(a[297] & b[382])^(a[296] & b[383])^(a[295] & b[384])^(a[294] & b[385])^(a[293] & b[386])^(a[292] & b[387])^(a[291] & b[388])^(a[290] & b[389])^(a[289] & b[390])^(a[288] & b[391])^(a[287] & b[392])^(a[286] & b[393])^(a[285] & b[394])^(a[284] & b[395])^(a[283] & b[396])^(a[282] & b[397])^(a[281] & b[398])^(a[280] & b[399])^(a[279] & b[400])^(a[278] & b[401])^(a[277] & b[402])^(a[276] & b[403])^(a[275] & b[404])^(a[274] & b[405])^(a[273] & b[406])^(a[272] & b[407])^(a[271] & b[408]);
assign y[680] = (a[408] & b[272])^(a[407] & b[273])^(a[406] & b[274])^(a[405] & b[275])^(a[404] & b[276])^(a[403] & b[277])^(a[402] & b[278])^(a[401] & b[279])^(a[400] & b[280])^(a[399] & b[281])^(a[398] & b[282])^(a[397] & b[283])^(a[396] & b[284])^(a[395] & b[285])^(a[394] & b[286])^(a[393] & b[287])^(a[392] & b[288])^(a[391] & b[289])^(a[390] & b[290])^(a[389] & b[291])^(a[388] & b[292])^(a[387] & b[293])^(a[386] & b[294])^(a[385] & b[295])^(a[384] & b[296])^(a[383] & b[297])^(a[382] & b[298])^(a[381] & b[299])^(a[380] & b[300])^(a[379] & b[301])^(a[378] & b[302])^(a[377] & b[303])^(a[376] & b[304])^(a[375] & b[305])^(a[374] & b[306])^(a[373] & b[307])^(a[372] & b[308])^(a[371] & b[309])^(a[370] & b[310])^(a[369] & b[311])^(a[368] & b[312])^(a[367] & b[313])^(a[366] & b[314])^(a[365] & b[315])^(a[364] & b[316])^(a[363] & b[317])^(a[362] & b[318])^(a[361] & b[319])^(a[360] & b[320])^(a[359] & b[321])^(a[358] & b[322])^(a[357] & b[323])^(a[356] & b[324])^(a[355] & b[325])^(a[354] & b[326])^(a[353] & b[327])^(a[352] & b[328])^(a[351] & b[329])^(a[350] & b[330])^(a[349] & b[331])^(a[348] & b[332])^(a[347] & b[333])^(a[346] & b[334])^(a[345] & b[335])^(a[344] & b[336])^(a[343] & b[337])^(a[342] & b[338])^(a[341] & b[339])^(a[340] & b[340])^(a[339] & b[341])^(a[338] & b[342])^(a[337] & b[343])^(a[336] & b[344])^(a[335] & b[345])^(a[334] & b[346])^(a[333] & b[347])^(a[332] & b[348])^(a[331] & b[349])^(a[330] & b[350])^(a[329] & b[351])^(a[328] & b[352])^(a[327] & b[353])^(a[326] & b[354])^(a[325] & b[355])^(a[324] & b[356])^(a[323] & b[357])^(a[322] & b[358])^(a[321] & b[359])^(a[320] & b[360])^(a[319] & b[361])^(a[318] & b[362])^(a[317] & b[363])^(a[316] & b[364])^(a[315] & b[365])^(a[314] & b[366])^(a[313] & b[367])^(a[312] & b[368])^(a[311] & b[369])^(a[310] & b[370])^(a[309] & b[371])^(a[308] & b[372])^(a[307] & b[373])^(a[306] & b[374])^(a[305] & b[375])^(a[304] & b[376])^(a[303] & b[377])^(a[302] & b[378])^(a[301] & b[379])^(a[300] & b[380])^(a[299] & b[381])^(a[298] & b[382])^(a[297] & b[383])^(a[296] & b[384])^(a[295] & b[385])^(a[294] & b[386])^(a[293] & b[387])^(a[292] & b[388])^(a[291] & b[389])^(a[290] & b[390])^(a[289] & b[391])^(a[288] & b[392])^(a[287] & b[393])^(a[286] & b[394])^(a[285] & b[395])^(a[284] & b[396])^(a[283] & b[397])^(a[282] & b[398])^(a[281] & b[399])^(a[280] & b[400])^(a[279] & b[401])^(a[278] & b[402])^(a[277] & b[403])^(a[276] & b[404])^(a[275] & b[405])^(a[274] & b[406])^(a[273] & b[407])^(a[272] & b[408]);
assign y[681] = (a[408] & b[273])^(a[407] & b[274])^(a[406] & b[275])^(a[405] & b[276])^(a[404] & b[277])^(a[403] & b[278])^(a[402] & b[279])^(a[401] & b[280])^(a[400] & b[281])^(a[399] & b[282])^(a[398] & b[283])^(a[397] & b[284])^(a[396] & b[285])^(a[395] & b[286])^(a[394] & b[287])^(a[393] & b[288])^(a[392] & b[289])^(a[391] & b[290])^(a[390] & b[291])^(a[389] & b[292])^(a[388] & b[293])^(a[387] & b[294])^(a[386] & b[295])^(a[385] & b[296])^(a[384] & b[297])^(a[383] & b[298])^(a[382] & b[299])^(a[381] & b[300])^(a[380] & b[301])^(a[379] & b[302])^(a[378] & b[303])^(a[377] & b[304])^(a[376] & b[305])^(a[375] & b[306])^(a[374] & b[307])^(a[373] & b[308])^(a[372] & b[309])^(a[371] & b[310])^(a[370] & b[311])^(a[369] & b[312])^(a[368] & b[313])^(a[367] & b[314])^(a[366] & b[315])^(a[365] & b[316])^(a[364] & b[317])^(a[363] & b[318])^(a[362] & b[319])^(a[361] & b[320])^(a[360] & b[321])^(a[359] & b[322])^(a[358] & b[323])^(a[357] & b[324])^(a[356] & b[325])^(a[355] & b[326])^(a[354] & b[327])^(a[353] & b[328])^(a[352] & b[329])^(a[351] & b[330])^(a[350] & b[331])^(a[349] & b[332])^(a[348] & b[333])^(a[347] & b[334])^(a[346] & b[335])^(a[345] & b[336])^(a[344] & b[337])^(a[343] & b[338])^(a[342] & b[339])^(a[341] & b[340])^(a[340] & b[341])^(a[339] & b[342])^(a[338] & b[343])^(a[337] & b[344])^(a[336] & b[345])^(a[335] & b[346])^(a[334] & b[347])^(a[333] & b[348])^(a[332] & b[349])^(a[331] & b[350])^(a[330] & b[351])^(a[329] & b[352])^(a[328] & b[353])^(a[327] & b[354])^(a[326] & b[355])^(a[325] & b[356])^(a[324] & b[357])^(a[323] & b[358])^(a[322] & b[359])^(a[321] & b[360])^(a[320] & b[361])^(a[319] & b[362])^(a[318] & b[363])^(a[317] & b[364])^(a[316] & b[365])^(a[315] & b[366])^(a[314] & b[367])^(a[313] & b[368])^(a[312] & b[369])^(a[311] & b[370])^(a[310] & b[371])^(a[309] & b[372])^(a[308] & b[373])^(a[307] & b[374])^(a[306] & b[375])^(a[305] & b[376])^(a[304] & b[377])^(a[303] & b[378])^(a[302] & b[379])^(a[301] & b[380])^(a[300] & b[381])^(a[299] & b[382])^(a[298] & b[383])^(a[297] & b[384])^(a[296] & b[385])^(a[295] & b[386])^(a[294] & b[387])^(a[293] & b[388])^(a[292] & b[389])^(a[291] & b[390])^(a[290] & b[391])^(a[289] & b[392])^(a[288] & b[393])^(a[287] & b[394])^(a[286] & b[395])^(a[285] & b[396])^(a[284] & b[397])^(a[283] & b[398])^(a[282] & b[399])^(a[281] & b[400])^(a[280] & b[401])^(a[279] & b[402])^(a[278] & b[403])^(a[277] & b[404])^(a[276] & b[405])^(a[275] & b[406])^(a[274] & b[407])^(a[273] & b[408]);
assign y[682] = (a[408] & b[274])^(a[407] & b[275])^(a[406] & b[276])^(a[405] & b[277])^(a[404] & b[278])^(a[403] & b[279])^(a[402] & b[280])^(a[401] & b[281])^(a[400] & b[282])^(a[399] & b[283])^(a[398] & b[284])^(a[397] & b[285])^(a[396] & b[286])^(a[395] & b[287])^(a[394] & b[288])^(a[393] & b[289])^(a[392] & b[290])^(a[391] & b[291])^(a[390] & b[292])^(a[389] & b[293])^(a[388] & b[294])^(a[387] & b[295])^(a[386] & b[296])^(a[385] & b[297])^(a[384] & b[298])^(a[383] & b[299])^(a[382] & b[300])^(a[381] & b[301])^(a[380] & b[302])^(a[379] & b[303])^(a[378] & b[304])^(a[377] & b[305])^(a[376] & b[306])^(a[375] & b[307])^(a[374] & b[308])^(a[373] & b[309])^(a[372] & b[310])^(a[371] & b[311])^(a[370] & b[312])^(a[369] & b[313])^(a[368] & b[314])^(a[367] & b[315])^(a[366] & b[316])^(a[365] & b[317])^(a[364] & b[318])^(a[363] & b[319])^(a[362] & b[320])^(a[361] & b[321])^(a[360] & b[322])^(a[359] & b[323])^(a[358] & b[324])^(a[357] & b[325])^(a[356] & b[326])^(a[355] & b[327])^(a[354] & b[328])^(a[353] & b[329])^(a[352] & b[330])^(a[351] & b[331])^(a[350] & b[332])^(a[349] & b[333])^(a[348] & b[334])^(a[347] & b[335])^(a[346] & b[336])^(a[345] & b[337])^(a[344] & b[338])^(a[343] & b[339])^(a[342] & b[340])^(a[341] & b[341])^(a[340] & b[342])^(a[339] & b[343])^(a[338] & b[344])^(a[337] & b[345])^(a[336] & b[346])^(a[335] & b[347])^(a[334] & b[348])^(a[333] & b[349])^(a[332] & b[350])^(a[331] & b[351])^(a[330] & b[352])^(a[329] & b[353])^(a[328] & b[354])^(a[327] & b[355])^(a[326] & b[356])^(a[325] & b[357])^(a[324] & b[358])^(a[323] & b[359])^(a[322] & b[360])^(a[321] & b[361])^(a[320] & b[362])^(a[319] & b[363])^(a[318] & b[364])^(a[317] & b[365])^(a[316] & b[366])^(a[315] & b[367])^(a[314] & b[368])^(a[313] & b[369])^(a[312] & b[370])^(a[311] & b[371])^(a[310] & b[372])^(a[309] & b[373])^(a[308] & b[374])^(a[307] & b[375])^(a[306] & b[376])^(a[305] & b[377])^(a[304] & b[378])^(a[303] & b[379])^(a[302] & b[380])^(a[301] & b[381])^(a[300] & b[382])^(a[299] & b[383])^(a[298] & b[384])^(a[297] & b[385])^(a[296] & b[386])^(a[295] & b[387])^(a[294] & b[388])^(a[293] & b[389])^(a[292] & b[390])^(a[291] & b[391])^(a[290] & b[392])^(a[289] & b[393])^(a[288] & b[394])^(a[287] & b[395])^(a[286] & b[396])^(a[285] & b[397])^(a[284] & b[398])^(a[283] & b[399])^(a[282] & b[400])^(a[281] & b[401])^(a[280] & b[402])^(a[279] & b[403])^(a[278] & b[404])^(a[277] & b[405])^(a[276] & b[406])^(a[275] & b[407])^(a[274] & b[408]);
assign y[683] = (a[408] & b[275])^(a[407] & b[276])^(a[406] & b[277])^(a[405] & b[278])^(a[404] & b[279])^(a[403] & b[280])^(a[402] & b[281])^(a[401] & b[282])^(a[400] & b[283])^(a[399] & b[284])^(a[398] & b[285])^(a[397] & b[286])^(a[396] & b[287])^(a[395] & b[288])^(a[394] & b[289])^(a[393] & b[290])^(a[392] & b[291])^(a[391] & b[292])^(a[390] & b[293])^(a[389] & b[294])^(a[388] & b[295])^(a[387] & b[296])^(a[386] & b[297])^(a[385] & b[298])^(a[384] & b[299])^(a[383] & b[300])^(a[382] & b[301])^(a[381] & b[302])^(a[380] & b[303])^(a[379] & b[304])^(a[378] & b[305])^(a[377] & b[306])^(a[376] & b[307])^(a[375] & b[308])^(a[374] & b[309])^(a[373] & b[310])^(a[372] & b[311])^(a[371] & b[312])^(a[370] & b[313])^(a[369] & b[314])^(a[368] & b[315])^(a[367] & b[316])^(a[366] & b[317])^(a[365] & b[318])^(a[364] & b[319])^(a[363] & b[320])^(a[362] & b[321])^(a[361] & b[322])^(a[360] & b[323])^(a[359] & b[324])^(a[358] & b[325])^(a[357] & b[326])^(a[356] & b[327])^(a[355] & b[328])^(a[354] & b[329])^(a[353] & b[330])^(a[352] & b[331])^(a[351] & b[332])^(a[350] & b[333])^(a[349] & b[334])^(a[348] & b[335])^(a[347] & b[336])^(a[346] & b[337])^(a[345] & b[338])^(a[344] & b[339])^(a[343] & b[340])^(a[342] & b[341])^(a[341] & b[342])^(a[340] & b[343])^(a[339] & b[344])^(a[338] & b[345])^(a[337] & b[346])^(a[336] & b[347])^(a[335] & b[348])^(a[334] & b[349])^(a[333] & b[350])^(a[332] & b[351])^(a[331] & b[352])^(a[330] & b[353])^(a[329] & b[354])^(a[328] & b[355])^(a[327] & b[356])^(a[326] & b[357])^(a[325] & b[358])^(a[324] & b[359])^(a[323] & b[360])^(a[322] & b[361])^(a[321] & b[362])^(a[320] & b[363])^(a[319] & b[364])^(a[318] & b[365])^(a[317] & b[366])^(a[316] & b[367])^(a[315] & b[368])^(a[314] & b[369])^(a[313] & b[370])^(a[312] & b[371])^(a[311] & b[372])^(a[310] & b[373])^(a[309] & b[374])^(a[308] & b[375])^(a[307] & b[376])^(a[306] & b[377])^(a[305] & b[378])^(a[304] & b[379])^(a[303] & b[380])^(a[302] & b[381])^(a[301] & b[382])^(a[300] & b[383])^(a[299] & b[384])^(a[298] & b[385])^(a[297] & b[386])^(a[296] & b[387])^(a[295] & b[388])^(a[294] & b[389])^(a[293] & b[390])^(a[292] & b[391])^(a[291] & b[392])^(a[290] & b[393])^(a[289] & b[394])^(a[288] & b[395])^(a[287] & b[396])^(a[286] & b[397])^(a[285] & b[398])^(a[284] & b[399])^(a[283] & b[400])^(a[282] & b[401])^(a[281] & b[402])^(a[280] & b[403])^(a[279] & b[404])^(a[278] & b[405])^(a[277] & b[406])^(a[276] & b[407])^(a[275] & b[408]);
assign y[684] = (a[408] & b[276])^(a[407] & b[277])^(a[406] & b[278])^(a[405] & b[279])^(a[404] & b[280])^(a[403] & b[281])^(a[402] & b[282])^(a[401] & b[283])^(a[400] & b[284])^(a[399] & b[285])^(a[398] & b[286])^(a[397] & b[287])^(a[396] & b[288])^(a[395] & b[289])^(a[394] & b[290])^(a[393] & b[291])^(a[392] & b[292])^(a[391] & b[293])^(a[390] & b[294])^(a[389] & b[295])^(a[388] & b[296])^(a[387] & b[297])^(a[386] & b[298])^(a[385] & b[299])^(a[384] & b[300])^(a[383] & b[301])^(a[382] & b[302])^(a[381] & b[303])^(a[380] & b[304])^(a[379] & b[305])^(a[378] & b[306])^(a[377] & b[307])^(a[376] & b[308])^(a[375] & b[309])^(a[374] & b[310])^(a[373] & b[311])^(a[372] & b[312])^(a[371] & b[313])^(a[370] & b[314])^(a[369] & b[315])^(a[368] & b[316])^(a[367] & b[317])^(a[366] & b[318])^(a[365] & b[319])^(a[364] & b[320])^(a[363] & b[321])^(a[362] & b[322])^(a[361] & b[323])^(a[360] & b[324])^(a[359] & b[325])^(a[358] & b[326])^(a[357] & b[327])^(a[356] & b[328])^(a[355] & b[329])^(a[354] & b[330])^(a[353] & b[331])^(a[352] & b[332])^(a[351] & b[333])^(a[350] & b[334])^(a[349] & b[335])^(a[348] & b[336])^(a[347] & b[337])^(a[346] & b[338])^(a[345] & b[339])^(a[344] & b[340])^(a[343] & b[341])^(a[342] & b[342])^(a[341] & b[343])^(a[340] & b[344])^(a[339] & b[345])^(a[338] & b[346])^(a[337] & b[347])^(a[336] & b[348])^(a[335] & b[349])^(a[334] & b[350])^(a[333] & b[351])^(a[332] & b[352])^(a[331] & b[353])^(a[330] & b[354])^(a[329] & b[355])^(a[328] & b[356])^(a[327] & b[357])^(a[326] & b[358])^(a[325] & b[359])^(a[324] & b[360])^(a[323] & b[361])^(a[322] & b[362])^(a[321] & b[363])^(a[320] & b[364])^(a[319] & b[365])^(a[318] & b[366])^(a[317] & b[367])^(a[316] & b[368])^(a[315] & b[369])^(a[314] & b[370])^(a[313] & b[371])^(a[312] & b[372])^(a[311] & b[373])^(a[310] & b[374])^(a[309] & b[375])^(a[308] & b[376])^(a[307] & b[377])^(a[306] & b[378])^(a[305] & b[379])^(a[304] & b[380])^(a[303] & b[381])^(a[302] & b[382])^(a[301] & b[383])^(a[300] & b[384])^(a[299] & b[385])^(a[298] & b[386])^(a[297] & b[387])^(a[296] & b[388])^(a[295] & b[389])^(a[294] & b[390])^(a[293] & b[391])^(a[292] & b[392])^(a[291] & b[393])^(a[290] & b[394])^(a[289] & b[395])^(a[288] & b[396])^(a[287] & b[397])^(a[286] & b[398])^(a[285] & b[399])^(a[284] & b[400])^(a[283] & b[401])^(a[282] & b[402])^(a[281] & b[403])^(a[280] & b[404])^(a[279] & b[405])^(a[278] & b[406])^(a[277] & b[407])^(a[276] & b[408]);
assign y[685] = (a[408] & b[277])^(a[407] & b[278])^(a[406] & b[279])^(a[405] & b[280])^(a[404] & b[281])^(a[403] & b[282])^(a[402] & b[283])^(a[401] & b[284])^(a[400] & b[285])^(a[399] & b[286])^(a[398] & b[287])^(a[397] & b[288])^(a[396] & b[289])^(a[395] & b[290])^(a[394] & b[291])^(a[393] & b[292])^(a[392] & b[293])^(a[391] & b[294])^(a[390] & b[295])^(a[389] & b[296])^(a[388] & b[297])^(a[387] & b[298])^(a[386] & b[299])^(a[385] & b[300])^(a[384] & b[301])^(a[383] & b[302])^(a[382] & b[303])^(a[381] & b[304])^(a[380] & b[305])^(a[379] & b[306])^(a[378] & b[307])^(a[377] & b[308])^(a[376] & b[309])^(a[375] & b[310])^(a[374] & b[311])^(a[373] & b[312])^(a[372] & b[313])^(a[371] & b[314])^(a[370] & b[315])^(a[369] & b[316])^(a[368] & b[317])^(a[367] & b[318])^(a[366] & b[319])^(a[365] & b[320])^(a[364] & b[321])^(a[363] & b[322])^(a[362] & b[323])^(a[361] & b[324])^(a[360] & b[325])^(a[359] & b[326])^(a[358] & b[327])^(a[357] & b[328])^(a[356] & b[329])^(a[355] & b[330])^(a[354] & b[331])^(a[353] & b[332])^(a[352] & b[333])^(a[351] & b[334])^(a[350] & b[335])^(a[349] & b[336])^(a[348] & b[337])^(a[347] & b[338])^(a[346] & b[339])^(a[345] & b[340])^(a[344] & b[341])^(a[343] & b[342])^(a[342] & b[343])^(a[341] & b[344])^(a[340] & b[345])^(a[339] & b[346])^(a[338] & b[347])^(a[337] & b[348])^(a[336] & b[349])^(a[335] & b[350])^(a[334] & b[351])^(a[333] & b[352])^(a[332] & b[353])^(a[331] & b[354])^(a[330] & b[355])^(a[329] & b[356])^(a[328] & b[357])^(a[327] & b[358])^(a[326] & b[359])^(a[325] & b[360])^(a[324] & b[361])^(a[323] & b[362])^(a[322] & b[363])^(a[321] & b[364])^(a[320] & b[365])^(a[319] & b[366])^(a[318] & b[367])^(a[317] & b[368])^(a[316] & b[369])^(a[315] & b[370])^(a[314] & b[371])^(a[313] & b[372])^(a[312] & b[373])^(a[311] & b[374])^(a[310] & b[375])^(a[309] & b[376])^(a[308] & b[377])^(a[307] & b[378])^(a[306] & b[379])^(a[305] & b[380])^(a[304] & b[381])^(a[303] & b[382])^(a[302] & b[383])^(a[301] & b[384])^(a[300] & b[385])^(a[299] & b[386])^(a[298] & b[387])^(a[297] & b[388])^(a[296] & b[389])^(a[295] & b[390])^(a[294] & b[391])^(a[293] & b[392])^(a[292] & b[393])^(a[291] & b[394])^(a[290] & b[395])^(a[289] & b[396])^(a[288] & b[397])^(a[287] & b[398])^(a[286] & b[399])^(a[285] & b[400])^(a[284] & b[401])^(a[283] & b[402])^(a[282] & b[403])^(a[281] & b[404])^(a[280] & b[405])^(a[279] & b[406])^(a[278] & b[407])^(a[277] & b[408]);
assign y[686] = (a[408] & b[278])^(a[407] & b[279])^(a[406] & b[280])^(a[405] & b[281])^(a[404] & b[282])^(a[403] & b[283])^(a[402] & b[284])^(a[401] & b[285])^(a[400] & b[286])^(a[399] & b[287])^(a[398] & b[288])^(a[397] & b[289])^(a[396] & b[290])^(a[395] & b[291])^(a[394] & b[292])^(a[393] & b[293])^(a[392] & b[294])^(a[391] & b[295])^(a[390] & b[296])^(a[389] & b[297])^(a[388] & b[298])^(a[387] & b[299])^(a[386] & b[300])^(a[385] & b[301])^(a[384] & b[302])^(a[383] & b[303])^(a[382] & b[304])^(a[381] & b[305])^(a[380] & b[306])^(a[379] & b[307])^(a[378] & b[308])^(a[377] & b[309])^(a[376] & b[310])^(a[375] & b[311])^(a[374] & b[312])^(a[373] & b[313])^(a[372] & b[314])^(a[371] & b[315])^(a[370] & b[316])^(a[369] & b[317])^(a[368] & b[318])^(a[367] & b[319])^(a[366] & b[320])^(a[365] & b[321])^(a[364] & b[322])^(a[363] & b[323])^(a[362] & b[324])^(a[361] & b[325])^(a[360] & b[326])^(a[359] & b[327])^(a[358] & b[328])^(a[357] & b[329])^(a[356] & b[330])^(a[355] & b[331])^(a[354] & b[332])^(a[353] & b[333])^(a[352] & b[334])^(a[351] & b[335])^(a[350] & b[336])^(a[349] & b[337])^(a[348] & b[338])^(a[347] & b[339])^(a[346] & b[340])^(a[345] & b[341])^(a[344] & b[342])^(a[343] & b[343])^(a[342] & b[344])^(a[341] & b[345])^(a[340] & b[346])^(a[339] & b[347])^(a[338] & b[348])^(a[337] & b[349])^(a[336] & b[350])^(a[335] & b[351])^(a[334] & b[352])^(a[333] & b[353])^(a[332] & b[354])^(a[331] & b[355])^(a[330] & b[356])^(a[329] & b[357])^(a[328] & b[358])^(a[327] & b[359])^(a[326] & b[360])^(a[325] & b[361])^(a[324] & b[362])^(a[323] & b[363])^(a[322] & b[364])^(a[321] & b[365])^(a[320] & b[366])^(a[319] & b[367])^(a[318] & b[368])^(a[317] & b[369])^(a[316] & b[370])^(a[315] & b[371])^(a[314] & b[372])^(a[313] & b[373])^(a[312] & b[374])^(a[311] & b[375])^(a[310] & b[376])^(a[309] & b[377])^(a[308] & b[378])^(a[307] & b[379])^(a[306] & b[380])^(a[305] & b[381])^(a[304] & b[382])^(a[303] & b[383])^(a[302] & b[384])^(a[301] & b[385])^(a[300] & b[386])^(a[299] & b[387])^(a[298] & b[388])^(a[297] & b[389])^(a[296] & b[390])^(a[295] & b[391])^(a[294] & b[392])^(a[293] & b[393])^(a[292] & b[394])^(a[291] & b[395])^(a[290] & b[396])^(a[289] & b[397])^(a[288] & b[398])^(a[287] & b[399])^(a[286] & b[400])^(a[285] & b[401])^(a[284] & b[402])^(a[283] & b[403])^(a[282] & b[404])^(a[281] & b[405])^(a[280] & b[406])^(a[279] & b[407])^(a[278] & b[408]);
assign y[687] = (a[408] & b[279])^(a[407] & b[280])^(a[406] & b[281])^(a[405] & b[282])^(a[404] & b[283])^(a[403] & b[284])^(a[402] & b[285])^(a[401] & b[286])^(a[400] & b[287])^(a[399] & b[288])^(a[398] & b[289])^(a[397] & b[290])^(a[396] & b[291])^(a[395] & b[292])^(a[394] & b[293])^(a[393] & b[294])^(a[392] & b[295])^(a[391] & b[296])^(a[390] & b[297])^(a[389] & b[298])^(a[388] & b[299])^(a[387] & b[300])^(a[386] & b[301])^(a[385] & b[302])^(a[384] & b[303])^(a[383] & b[304])^(a[382] & b[305])^(a[381] & b[306])^(a[380] & b[307])^(a[379] & b[308])^(a[378] & b[309])^(a[377] & b[310])^(a[376] & b[311])^(a[375] & b[312])^(a[374] & b[313])^(a[373] & b[314])^(a[372] & b[315])^(a[371] & b[316])^(a[370] & b[317])^(a[369] & b[318])^(a[368] & b[319])^(a[367] & b[320])^(a[366] & b[321])^(a[365] & b[322])^(a[364] & b[323])^(a[363] & b[324])^(a[362] & b[325])^(a[361] & b[326])^(a[360] & b[327])^(a[359] & b[328])^(a[358] & b[329])^(a[357] & b[330])^(a[356] & b[331])^(a[355] & b[332])^(a[354] & b[333])^(a[353] & b[334])^(a[352] & b[335])^(a[351] & b[336])^(a[350] & b[337])^(a[349] & b[338])^(a[348] & b[339])^(a[347] & b[340])^(a[346] & b[341])^(a[345] & b[342])^(a[344] & b[343])^(a[343] & b[344])^(a[342] & b[345])^(a[341] & b[346])^(a[340] & b[347])^(a[339] & b[348])^(a[338] & b[349])^(a[337] & b[350])^(a[336] & b[351])^(a[335] & b[352])^(a[334] & b[353])^(a[333] & b[354])^(a[332] & b[355])^(a[331] & b[356])^(a[330] & b[357])^(a[329] & b[358])^(a[328] & b[359])^(a[327] & b[360])^(a[326] & b[361])^(a[325] & b[362])^(a[324] & b[363])^(a[323] & b[364])^(a[322] & b[365])^(a[321] & b[366])^(a[320] & b[367])^(a[319] & b[368])^(a[318] & b[369])^(a[317] & b[370])^(a[316] & b[371])^(a[315] & b[372])^(a[314] & b[373])^(a[313] & b[374])^(a[312] & b[375])^(a[311] & b[376])^(a[310] & b[377])^(a[309] & b[378])^(a[308] & b[379])^(a[307] & b[380])^(a[306] & b[381])^(a[305] & b[382])^(a[304] & b[383])^(a[303] & b[384])^(a[302] & b[385])^(a[301] & b[386])^(a[300] & b[387])^(a[299] & b[388])^(a[298] & b[389])^(a[297] & b[390])^(a[296] & b[391])^(a[295] & b[392])^(a[294] & b[393])^(a[293] & b[394])^(a[292] & b[395])^(a[291] & b[396])^(a[290] & b[397])^(a[289] & b[398])^(a[288] & b[399])^(a[287] & b[400])^(a[286] & b[401])^(a[285] & b[402])^(a[284] & b[403])^(a[283] & b[404])^(a[282] & b[405])^(a[281] & b[406])^(a[280] & b[407])^(a[279] & b[408]);
assign y[688] = (a[408] & b[280])^(a[407] & b[281])^(a[406] & b[282])^(a[405] & b[283])^(a[404] & b[284])^(a[403] & b[285])^(a[402] & b[286])^(a[401] & b[287])^(a[400] & b[288])^(a[399] & b[289])^(a[398] & b[290])^(a[397] & b[291])^(a[396] & b[292])^(a[395] & b[293])^(a[394] & b[294])^(a[393] & b[295])^(a[392] & b[296])^(a[391] & b[297])^(a[390] & b[298])^(a[389] & b[299])^(a[388] & b[300])^(a[387] & b[301])^(a[386] & b[302])^(a[385] & b[303])^(a[384] & b[304])^(a[383] & b[305])^(a[382] & b[306])^(a[381] & b[307])^(a[380] & b[308])^(a[379] & b[309])^(a[378] & b[310])^(a[377] & b[311])^(a[376] & b[312])^(a[375] & b[313])^(a[374] & b[314])^(a[373] & b[315])^(a[372] & b[316])^(a[371] & b[317])^(a[370] & b[318])^(a[369] & b[319])^(a[368] & b[320])^(a[367] & b[321])^(a[366] & b[322])^(a[365] & b[323])^(a[364] & b[324])^(a[363] & b[325])^(a[362] & b[326])^(a[361] & b[327])^(a[360] & b[328])^(a[359] & b[329])^(a[358] & b[330])^(a[357] & b[331])^(a[356] & b[332])^(a[355] & b[333])^(a[354] & b[334])^(a[353] & b[335])^(a[352] & b[336])^(a[351] & b[337])^(a[350] & b[338])^(a[349] & b[339])^(a[348] & b[340])^(a[347] & b[341])^(a[346] & b[342])^(a[345] & b[343])^(a[344] & b[344])^(a[343] & b[345])^(a[342] & b[346])^(a[341] & b[347])^(a[340] & b[348])^(a[339] & b[349])^(a[338] & b[350])^(a[337] & b[351])^(a[336] & b[352])^(a[335] & b[353])^(a[334] & b[354])^(a[333] & b[355])^(a[332] & b[356])^(a[331] & b[357])^(a[330] & b[358])^(a[329] & b[359])^(a[328] & b[360])^(a[327] & b[361])^(a[326] & b[362])^(a[325] & b[363])^(a[324] & b[364])^(a[323] & b[365])^(a[322] & b[366])^(a[321] & b[367])^(a[320] & b[368])^(a[319] & b[369])^(a[318] & b[370])^(a[317] & b[371])^(a[316] & b[372])^(a[315] & b[373])^(a[314] & b[374])^(a[313] & b[375])^(a[312] & b[376])^(a[311] & b[377])^(a[310] & b[378])^(a[309] & b[379])^(a[308] & b[380])^(a[307] & b[381])^(a[306] & b[382])^(a[305] & b[383])^(a[304] & b[384])^(a[303] & b[385])^(a[302] & b[386])^(a[301] & b[387])^(a[300] & b[388])^(a[299] & b[389])^(a[298] & b[390])^(a[297] & b[391])^(a[296] & b[392])^(a[295] & b[393])^(a[294] & b[394])^(a[293] & b[395])^(a[292] & b[396])^(a[291] & b[397])^(a[290] & b[398])^(a[289] & b[399])^(a[288] & b[400])^(a[287] & b[401])^(a[286] & b[402])^(a[285] & b[403])^(a[284] & b[404])^(a[283] & b[405])^(a[282] & b[406])^(a[281] & b[407])^(a[280] & b[408]);
assign y[689] = (a[408] & b[281])^(a[407] & b[282])^(a[406] & b[283])^(a[405] & b[284])^(a[404] & b[285])^(a[403] & b[286])^(a[402] & b[287])^(a[401] & b[288])^(a[400] & b[289])^(a[399] & b[290])^(a[398] & b[291])^(a[397] & b[292])^(a[396] & b[293])^(a[395] & b[294])^(a[394] & b[295])^(a[393] & b[296])^(a[392] & b[297])^(a[391] & b[298])^(a[390] & b[299])^(a[389] & b[300])^(a[388] & b[301])^(a[387] & b[302])^(a[386] & b[303])^(a[385] & b[304])^(a[384] & b[305])^(a[383] & b[306])^(a[382] & b[307])^(a[381] & b[308])^(a[380] & b[309])^(a[379] & b[310])^(a[378] & b[311])^(a[377] & b[312])^(a[376] & b[313])^(a[375] & b[314])^(a[374] & b[315])^(a[373] & b[316])^(a[372] & b[317])^(a[371] & b[318])^(a[370] & b[319])^(a[369] & b[320])^(a[368] & b[321])^(a[367] & b[322])^(a[366] & b[323])^(a[365] & b[324])^(a[364] & b[325])^(a[363] & b[326])^(a[362] & b[327])^(a[361] & b[328])^(a[360] & b[329])^(a[359] & b[330])^(a[358] & b[331])^(a[357] & b[332])^(a[356] & b[333])^(a[355] & b[334])^(a[354] & b[335])^(a[353] & b[336])^(a[352] & b[337])^(a[351] & b[338])^(a[350] & b[339])^(a[349] & b[340])^(a[348] & b[341])^(a[347] & b[342])^(a[346] & b[343])^(a[345] & b[344])^(a[344] & b[345])^(a[343] & b[346])^(a[342] & b[347])^(a[341] & b[348])^(a[340] & b[349])^(a[339] & b[350])^(a[338] & b[351])^(a[337] & b[352])^(a[336] & b[353])^(a[335] & b[354])^(a[334] & b[355])^(a[333] & b[356])^(a[332] & b[357])^(a[331] & b[358])^(a[330] & b[359])^(a[329] & b[360])^(a[328] & b[361])^(a[327] & b[362])^(a[326] & b[363])^(a[325] & b[364])^(a[324] & b[365])^(a[323] & b[366])^(a[322] & b[367])^(a[321] & b[368])^(a[320] & b[369])^(a[319] & b[370])^(a[318] & b[371])^(a[317] & b[372])^(a[316] & b[373])^(a[315] & b[374])^(a[314] & b[375])^(a[313] & b[376])^(a[312] & b[377])^(a[311] & b[378])^(a[310] & b[379])^(a[309] & b[380])^(a[308] & b[381])^(a[307] & b[382])^(a[306] & b[383])^(a[305] & b[384])^(a[304] & b[385])^(a[303] & b[386])^(a[302] & b[387])^(a[301] & b[388])^(a[300] & b[389])^(a[299] & b[390])^(a[298] & b[391])^(a[297] & b[392])^(a[296] & b[393])^(a[295] & b[394])^(a[294] & b[395])^(a[293] & b[396])^(a[292] & b[397])^(a[291] & b[398])^(a[290] & b[399])^(a[289] & b[400])^(a[288] & b[401])^(a[287] & b[402])^(a[286] & b[403])^(a[285] & b[404])^(a[284] & b[405])^(a[283] & b[406])^(a[282] & b[407])^(a[281] & b[408]);
assign y[690] = (a[408] & b[282])^(a[407] & b[283])^(a[406] & b[284])^(a[405] & b[285])^(a[404] & b[286])^(a[403] & b[287])^(a[402] & b[288])^(a[401] & b[289])^(a[400] & b[290])^(a[399] & b[291])^(a[398] & b[292])^(a[397] & b[293])^(a[396] & b[294])^(a[395] & b[295])^(a[394] & b[296])^(a[393] & b[297])^(a[392] & b[298])^(a[391] & b[299])^(a[390] & b[300])^(a[389] & b[301])^(a[388] & b[302])^(a[387] & b[303])^(a[386] & b[304])^(a[385] & b[305])^(a[384] & b[306])^(a[383] & b[307])^(a[382] & b[308])^(a[381] & b[309])^(a[380] & b[310])^(a[379] & b[311])^(a[378] & b[312])^(a[377] & b[313])^(a[376] & b[314])^(a[375] & b[315])^(a[374] & b[316])^(a[373] & b[317])^(a[372] & b[318])^(a[371] & b[319])^(a[370] & b[320])^(a[369] & b[321])^(a[368] & b[322])^(a[367] & b[323])^(a[366] & b[324])^(a[365] & b[325])^(a[364] & b[326])^(a[363] & b[327])^(a[362] & b[328])^(a[361] & b[329])^(a[360] & b[330])^(a[359] & b[331])^(a[358] & b[332])^(a[357] & b[333])^(a[356] & b[334])^(a[355] & b[335])^(a[354] & b[336])^(a[353] & b[337])^(a[352] & b[338])^(a[351] & b[339])^(a[350] & b[340])^(a[349] & b[341])^(a[348] & b[342])^(a[347] & b[343])^(a[346] & b[344])^(a[345] & b[345])^(a[344] & b[346])^(a[343] & b[347])^(a[342] & b[348])^(a[341] & b[349])^(a[340] & b[350])^(a[339] & b[351])^(a[338] & b[352])^(a[337] & b[353])^(a[336] & b[354])^(a[335] & b[355])^(a[334] & b[356])^(a[333] & b[357])^(a[332] & b[358])^(a[331] & b[359])^(a[330] & b[360])^(a[329] & b[361])^(a[328] & b[362])^(a[327] & b[363])^(a[326] & b[364])^(a[325] & b[365])^(a[324] & b[366])^(a[323] & b[367])^(a[322] & b[368])^(a[321] & b[369])^(a[320] & b[370])^(a[319] & b[371])^(a[318] & b[372])^(a[317] & b[373])^(a[316] & b[374])^(a[315] & b[375])^(a[314] & b[376])^(a[313] & b[377])^(a[312] & b[378])^(a[311] & b[379])^(a[310] & b[380])^(a[309] & b[381])^(a[308] & b[382])^(a[307] & b[383])^(a[306] & b[384])^(a[305] & b[385])^(a[304] & b[386])^(a[303] & b[387])^(a[302] & b[388])^(a[301] & b[389])^(a[300] & b[390])^(a[299] & b[391])^(a[298] & b[392])^(a[297] & b[393])^(a[296] & b[394])^(a[295] & b[395])^(a[294] & b[396])^(a[293] & b[397])^(a[292] & b[398])^(a[291] & b[399])^(a[290] & b[400])^(a[289] & b[401])^(a[288] & b[402])^(a[287] & b[403])^(a[286] & b[404])^(a[285] & b[405])^(a[284] & b[406])^(a[283] & b[407])^(a[282] & b[408]);
assign y[691] = (a[408] & b[283])^(a[407] & b[284])^(a[406] & b[285])^(a[405] & b[286])^(a[404] & b[287])^(a[403] & b[288])^(a[402] & b[289])^(a[401] & b[290])^(a[400] & b[291])^(a[399] & b[292])^(a[398] & b[293])^(a[397] & b[294])^(a[396] & b[295])^(a[395] & b[296])^(a[394] & b[297])^(a[393] & b[298])^(a[392] & b[299])^(a[391] & b[300])^(a[390] & b[301])^(a[389] & b[302])^(a[388] & b[303])^(a[387] & b[304])^(a[386] & b[305])^(a[385] & b[306])^(a[384] & b[307])^(a[383] & b[308])^(a[382] & b[309])^(a[381] & b[310])^(a[380] & b[311])^(a[379] & b[312])^(a[378] & b[313])^(a[377] & b[314])^(a[376] & b[315])^(a[375] & b[316])^(a[374] & b[317])^(a[373] & b[318])^(a[372] & b[319])^(a[371] & b[320])^(a[370] & b[321])^(a[369] & b[322])^(a[368] & b[323])^(a[367] & b[324])^(a[366] & b[325])^(a[365] & b[326])^(a[364] & b[327])^(a[363] & b[328])^(a[362] & b[329])^(a[361] & b[330])^(a[360] & b[331])^(a[359] & b[332])^(a[358] & b[333])^(a[357] & b[334])^(a[356] & b[335])^(a[355] & b[336])^(a[354] & b[337])^(a[353] & b[338])^(a[352] & b[339])^(a[351] & b[340])^(a[350] & b[341])^(a[349] & b[342])^(a[348] & b[343])^(a[347] & b[344])^(a[346] & b[345])^(a[345] & b[346])^(a[344] & b[347])^(a[343] & b[348])^(a[342] & b[349])^(a[341] & b[350])^(a[340] & b[351])^(a[339] & b[352])^(a[338] & b[353])^(a[337] & b[354])^(a[336] & b[355])^(a[335] & b[356])^(a[334] & b[357])^(a[333] & b[358])^(a[332] & b[359])^(a[331] & b[360])^(a[330] & b[361])^(a[329] & b[362])^(a[328] & b[363])^(a[327] & b[364])^(a[326] & b[365])^(a[325] & b[366])^(a[324] & b[367])^(a[323] & b[368])^(a[322] & b[369])^(a[321] & b[370])^(a[320] & b[371])^(a[319] & b[372])^(a[318] & b[373])^(a[317] & b[374])^(a[316] & b[375])^(a[315] & b[376])^(a[314] & b[377])^(a[313] & b[378])^(a[312] & b[379])^(a[311] & b[380])^(a[310] & b[381])^(a[309] & b[382])^(a[308] & b[383])^(a[307] & b[384])^(a[306] & b[385])^(a[305] & b[386])^(a[304] & b[387])^(a[303] & b[388])^(a[302] & b[389])^(a[301] & b[390])^(a[300] & b[391])^(a[299] & b[392])^(a[298] & b[393])^(a[297] & b[394])^(a[296] & b[395])^(a[295] & b[396])^(a[294] & b[397])^(a[293] & b[398])^(a[292] & b[399])^(a[291] & b[400])^(a[290] & b[401])^(a[289] & b[402])^(a[288] & b[403])^(a[287] & b[404])^(a[286] & b[405])^(a[285] & b[406])^(a[284] & b[407])^(a[283] & b[408]);
assign y[692] = (a[408] & b[284])^(a[407] & b[285])^(a[406] & b[286])^(a[405] & b[287])^(a[404] & b[288])^(a[403] & b[289])^(a[402] & b[290])^(a[401] & b[291])^(a[400] & b[292])^(a[399] & b[293])^(a[398] & b[294])^(a[397] & b[295])^(a[396] & b[296])^(a[395] & b[297])^(a[394] & b[298])^(a[393] & b[299])^(a[392] & b[300])^(a[391] & b[301])^(a[390] & b[302])^(a[389] & b[303])^(a[388] & b[304])^(a[387] & b[305])^(a[386] & b[306])^(a[385] & b[307])^(a[384] & b[308])^(a[383] & b[309])^(a[382] & b[310])^(a[381] & b[311])^(a[380] & b[312])^(a[379] & b[313])^(a[378] & b[314])^(a[377] & b[315])^(a[376] & b[316])^(a[375] & b[317])^(a[374] & b[318])^(a[373] & b[319])^(a[372] & b[320])^(a[371] & b[321])^(a[370] & b[322])^(a[369] & b[323])^(a[368] & b[324])^(a[367] & b[325])^(a[366] & b[326])^(a[365] & b[327])^(a[364] & b[328])^(a[363] & b[329])^(a[362] & b[330])^(a[361] & b[331])^(a[360] & b[332])^(a[359] & b[333])^(a[358] & b[334])^(a[357] & b[335])^(a[356] & b[336])^(a[355] & b[337])^(a[354] & b[338])^(a[353] & b[339])^(a[352] & b[340])^(a[351] & b[341])^(a[350] & b[342])^(a[349] & b[343])^(a[348] & b[344])^(a[347] & b[345])^(a[346] & b[346])^(a[345] & b[347])^(a[344] & b[348])^(a[343] & b[349])^(a[342] & b[350])^(a[341] & b[351])^(a[340] & b[352])^(a[339] & b[353])^(a[338] & b[354])^(a[337] & b[355])^(a[336] & b[356])^(a[335] & b[357])^(a[334] & b[358])^(a[333] & b[359])^(a[332] & b[360])^(a[331] & b[361])^(a[330] & b[362])^(a[329] & b[363])^(a[328] & b[364])^(a[327] & b[365])^(a[326] & b[366])^(a[325] & b[367])^(a[324] & b[368])^(a[323] & b[369])^(a[322] & b[370])^(a[321] & b[371])^(a[320] & b[372])^(a[319] & b[373])^(a[318] & b[374])^(a[317] & b[375])^(a[316] & b[376])^(a[315] & b[377])^(a[314] & b[378])^(a[313] & b[379])^(a[312] & b[380])^(a[311] & b[381])^(a[310] & b[382])^(a[309] & b[383])^(a[308] & b[384])^(a[307] & b[385])^(a[306] & b[386])^(a[305] & b[387])^(a[304] & b[388])^(a[303] & b[389])^(a[302] & b[390])^(a[301] & b[391])^(a[300] & b[392])^(a[299] & b[393])^(a[298] & b[394])^(a[297] & b[395])^(a[296] & b[396])^(a[295] & b[397])^(a[294] & b[398])^(a[293] & b[399])^(a[292] & b[400])^(a[291] & b[401])^(a[290] & b[402])^(a[289] & b[403])^(a[288] & b[404])^(a[287] & b[405])^(a[286] & b[406])^(a[285] & b[407])^(a[284] & b[408]);
assign y[693] = (a[408] & b[285])^(a[407] & b[286])^(a[406] & b[287])^(a[405] & b[288])^(a[404] & b[289])^(a[403] & b[290])^(a[402] & b[291])^(a[401] & b[292])^(a[400] & b[293])^(a[399] & b[294])^(a[398] & b[295])^(a[397] & b[296])^(a[396] & b[297])^(a[395] & b[298])^(a[394] & b[299])^(a[393] & b[300])^(a[392] & b[301])^(a[391] & b[302])^(a[390] & b[303])^(a[389] & b[304])^(a[388] & b[305])^(a[387] & b[306])^(a[386] & b[307])^(a[385] & b[308])^(a[384] & b[309])^(a[383] & b[310])^(a[382] & b[311])^(a[381] & b[312])^(a[380] & b[313])^(a[379] & b[314])^(a[378] & b[315])^(a[377] & b[316])^(a[376] & b[317])^(a[375] & b[318])^(a[374] & b[319])^(a[373] & b[320])^(a[372] & b[321])^(a[371] & b[322])^(a[370] & b[323])^(a[369] & b[324])^(a[368] & b[325])^(a[367] & b[326])^(a[366] & b[327])^(a[365] & b[328])^(a[364] & b[329])^(a[363] & b[330])^(a[362] & b[331])^(a[361] & b[332])^(a[360] & b[333])^(a[359] & b[334])^(a[358] & b[335])^(a[357] & b[336])^(a[356] & b[337])^(a[355] & b[338])^(a[354] & b[339])^(a[353] & b[340])^(a[352] & b[341])^(a[351] & b[342])^(a[350] & b[343])^(a[349] & b[344])^(a[348] & b[345])^(a[347] & b[346])^(a[346] & b[347])^(a[345] & b[348])^(a[344] & b[349])^(a[343] & b[350])^(a[342] & b[351])^(a[341] & b[352])^(a[340] & b[353])^(a[339] & b[354])^(a[338] & b[355])^(a[337] & b[356])^(a[336] & b[357])^(a[335] & b[358])^(a[334] & b[359])^(a[333] & b[360])^(a[332] & b[361])^(a[331] & b[362])^(a[330] & b[363])^(a[329] & b[364])^(a[328] & b[365])^(a[327] & b[366])^(a[326] & b[367])^(a[325] & b[368])^(a[324] & b[369])^(a[323] & b[370])^(a[322] & b[371])^(a[321] & b[372])^(a[320] & b[373])^(a[319] & b[374])^(a[318] & b[375])^(a[317] & b[376])^(a[316] & b[377])^(a[315] & b[378])^(a[314] & b[379])^(a[313] & b[380])^(a[312] & b[381])^(a[311] & b[382])^(a[310] & b[383])^(a[309] & b[384])^(a[308] & b[385])^(a[307] & b[386])^(a[306] & b[387])^(a[305] & b[388])^(a[304] & b[389])^(a[303] & b[390])^(a[302] & b[391])^(a[301] & b[392])^(a[300] & b[393])^(a[299] & b[394])^(a[298] & b[395])^(a[297] & b[396])^(a[296] & b[397])^(a[295] & b[398])^(a[294] & b[399])^(a[293] & b[400])^(a[292] & b[401])^(a[291] & b[402])^(a[290] & b[403])^(a[289] & b[404])^(a[288] & b[405])^(a[287] & b[406])^(a[286] & b[407])^(a[285] & b[408]);
assign y[694] = (a[408] & b[286])^(a[407] & b[287])^(a[406] & b[288])^(a[405] & b[289])^(a[404] & b[290])^(a[403] & b[291])^(a[402] & b[292])^(a[401] & b[293])^(a[400] & b[294])^(a[399] & b[295])^(a[398] & b[296])^(a[397] & b[297])^(a[396] & b[298])^(a[395] & b[299])^(a[394] & b[300])^(a[393] & b[301])^(a[392] & b[302])^(a[391] & b[303])^(a[390] & b[304])^(a[389] & b[305])^(a[388] & b[306])^(a[387] & b[307])^(a[386] & b[308])^(a[385] & b[309])^(a[384] & b[310])^(a[383] & b[311])^(a[382] & b[312])^(a[381] & b[313])^(a[380] & b[314])^(a[379] & b[315])^(a[378] & b[316])^(a[377] & b[317])^(a[376] & b[318])^(a[375] & b[319])^(a[374] & b[320])^(a[373] & b[321])^(a[372] & b[322])^(a[371] & b[323])^(a[370] & b[324])^(a[369] & b[325])^(a[368] & b[326])^(a[367] & b[327])^(a[366] & b[328])^(a[365] & b[329])^(a[364] & b[330])^(a[363] & b[331])^(a[362] & b[332])^(a[361] & b[333])^(a[360] & b[334])^(a[359] & b[335])^(a[358] & b[336])^(a[357] & b[337])^(a[356] & b[338])^(a[355] & b[339])^(a[354] & b[340])^(a[353] & b[341])^(a[352] & b[342])^(a[351] & b[343])^(a[350] & b[344])^(a[349] & b[345])^(a[348] & b[346])^(a[347] & b[347])^(a[346] & b[348])^(a[345] & b[349])^(a[344] & b[350])^(a[343] & b[351])^(a[342] & b[352])^(a[341] & b[353])^(a[340] & b[354])^(a[339] & b[355])^(a[338] & b[356])^(a[337] & b[357])^(a[336] & b[358])^(a[335] & b[359])^(a[334] & b[360])^(a[333] & b[361])^(a[332] & b[362])^(a[331] & b[363])^(a[330] & b[364])^(a[329] & b[365])^(a[328] & b[366])^(a[327] & b[367])^(a[326] & b[368])^(a[325] & b[369])^(a[324] & b[370])^(a[323] & b[371])^(a[322] & b[372])^(a[321] & b[373])^(a[320] & b[374])^(a[319] & b[375])^(a[318] & b[376])^(a[317] & b[377])^(a[316] & b[378])^(a[315] & b[379])^(a[314] & b[380])^(a[313] & b[381])^(a[312] & b[382])^(a[311] & b[383])^(a[310] & b[384])^(a[309] & b[385])^(a[308] & b[386])^(a[307] & b[387])^(a[306] & b[388])^(a[305] & b[389])^(a[304] & b[390])^(a[303] & b[391])^(a[302] & b[392])^(a[301] & b[393])^(a[300] & b[394])^(a[299] & b[395])^(a[298] & b[396])^(a[297] & b[397])^(a[296] & b[398])^(a[295] & b[399])^(a[294] & b[400])^(a[293] & b[401])^(a[292] & b[402])^(a[291] & b[403])^(a[290] & b[404])^(a[289] & b[405])^(a[288] & b[406])^(a[287] & b[407])^(a[286] & b[408]);
assign y[695] = (a[408] & b[287])^(a[407] & b[288])^(a[406] & b[289])^(a[405] & b[290])^(a[404] & b[291])^(a[403] & b[292])^(a[402] & b[293])^(a[401] & b[294])^(a[400] & b[295])^(a[399] & b[296])^(a[398] & b[297])^(a[397] & b[298])^(a[396] & b[299])^(a[395] & b[300])^(a[394] & b[301])^(a[393] & b[302])^(a[392] & b[303])^(a[391] & b[304])^(a[390] & b[305])^(a[389] & b[306])^(a[388] & b[307])^(a[387] & b[308])^(a[386] & b[309])^(a[385] & b[310])^(a[384] & b[311])^(a[383] & b[312])^(a[382] & b[313])^(a[381] & b[314])^(a[380] & b[315])^(a[379] & b[316])^(a[378] & b[317])^(a[377] & b[318])^(a[376] & b[319])^(a[375] & b[320])^(a[374] & b[321])^(a[373] & b[322])^(a[372] & b[323])^(a[371] & b[324])^(a[370] & b[325])^(a[369] & b[326])^(a[368] & b[327])^(a[367] & b[328])^(a[366] & b[329])^(a[365] & b[330])^(a[364] & b[331])^(a[363] & b[332])^(a[362] & b[333])^(a[361] & b[334])^(a[360] & b[335])^(a[359] & b[336])^(a[358] & b[337])^(a[357] & b[338])^(a[356] & b[339])^(a[355] & b[340])^(a[354] & b[341])^(a[353] & b[342])^(a[352] & b[343])^(a[351] & b[344])^(a[350] & b[345])^(a[349] & b[346])^(a[348] & b[347])^(a[347] & b[348])^(a[346] & b[349])^(a[345] & b[350])^(a[344] & b[351])^(a[343] & b[352])^(a[342] & b[353])^(a[341] & b[354])^(a[340] & b[355])^(a[339] & b[356])^(a[338] & b[357])^(a[337] & b[358])^(a[336] & b[359])^(a[335] & b[360])^(a[334] & b[361])^(a[333] & b[362])^(a[332] & b[363])^(a[331] & b[364])^(a[330] & b[365])^(a[329] & b[366])^(a[328] & b[367])^(a[327] & b[368])^(a[326] & b[369])^(a[325] & b[370])^(a[324] & b[371])^(a[323] & b[372])^(a[322] & b[373])^(a[321] & b[374])^(a[320] & b[375])^(a[319] & b[376])^(a[318] & b[377])^(a[317] & b[378])^(a[316] & b[379])^(a[315] & b[380])^(a[314] & b[381])^(a[313] & b[382])^(a[312] & b[383])^(a[311] & b[384])^(a[310] & b[385])^(a[309] & b[386])^(a[308] & b[387])^(a[307] & b[388])^(a[306] & b[389])^(a[305] & b[390])^(a[304] & b[391])^(a[303] & b[392])^(a[302] & b[393])^(a[301] & b[394])^(a[300] & b[395])^(a[299] & b[396])^(a[298] & b[397])^(a[297] & b[398])^(a[296] & b[399])^(a[295] & b[400])^(a[294] & b[401])^(a[293] & b[402])^(a[292] & b[403])^(a[291] & b[404])^(a[290] & b[405])^(a[289] & b[406])^(a[288] & b[407])^(a[287] & b[408]);
assign y[696] = (a[408] & b[288])^(a[407] & b[289])^(a[406] & b[290])^(a[405] & b[291])^(a[404] & b[292])^(a[403] & b[293])^(a[402] & b[294])^(a[401] & b[295])^(a[400] & b[296])^(a[399] & b[297])^(a[398] & b[298])^(a[397] & b[299])^(a[396] & b[300])^(a[395] & b[301])^(a[394] & b[302])^(a[393] & b[303])^(a[392] & b[304])^(a[391] & b[305])^(a[390] & b[306])^(a[389] & b[307])^(a[388] & b[308])^(a[387] & b[309])^(a[386] & b[310])^(a[385] & b[311])^(a[384] & b[312])^(a[383] & b[313])^(a[382] & b[314])^(a[381] & b[315])^(a[380] & b[316])^(a[379] & b[317])^(a[378] & b[318])^(a[377] & b[319])^(a[376] & b[320])^(a[375] & b[321])^(a[374] & b[322])^(a[373] & b[323])^(a[372] & b[324])^(a[371] & b[325])^(a[370] & b[326])^(a[369] & b[327])^(a[368] & b[328])^(a[367] & b[329])^(a[366] & b[330])^(a[365] & b[331])^(a[364] & b[332])^(a[363] & b[333])^(a[362] & b[334])^(a[361] & b[335])^(a[360] & b[336])^(a[359] & b[337])^(a[358] & b[338])^(a[357] & b[339])^(a[356] & b[340])^(a[355] & b[341])^(a[354] & b[342])^(a[353] & b[343])^(a[352] & b[344])^(a[351] & b[345])^(a[350] & b[346])^(a[349] & b[347])^(a[348] & b[348])^(a[347] & b[349])^(a[346] & b[350])^(a[345] & b[351])^(a[344] & b[352])^(a[343] & b[353])^(a[342] & b[354])^(a[341] & b[355])^(a[340] & b[356])^(a[339] & b[357])^(a[338] & b[358])^(a[337] & b[359])^(a[336] & b[360])^(a[335] & b[361])^(a[334] & b[362])^(a[333] & b[363])^(a[332] & b[364])^(a[331] & b[365])^(a[330] & b[366])^(a[329] & b[367])^(a[328] & b[368])^(a[327] & b[369])^(a[326] & b[370])^(a[325] & b[371])^(a[324] & b[372])^(a[323] & b[373])^(a[322] & b[374])^(a[321] & b[375])^(a[320] & b[376])^(a[319] & b[377])^(a[318] & b[378])^(a[317] & b[379])^(a[316] & b[380])^(a[315] & b[381])^(a[314] & b[382])^(a[313] & b[383])^(a[312] & b[384])^(a[311] & b[385])^(a[310] & b[386])^(a[309] & b[387])^(a[308] & b[388])^(a[307] & b[389])^(a[306] & b[390])^(a[305] & b[391])^(a[304] & b[392])^(a[303] & b[393])^(a[302] & b[394])^(a[301] & b[395])^(a[300] & b[396])^(a[299] & b[397])^(a[298] & b[398])^(a[297] & b[399])^(a[296] & b[400])^(a[295] & b[401])^(a[294] & b[402])^(a[293] & b[403])^(a[292] & b[404])^(a[291] & b[405])^(a[290] & b[406])^(a[289] & b[407])^(a[288] & b[408]);
assign y[697] = (a[408] & b[289])^(a[407] & b[290])^(a[406] & b[291])^(a[405] & b[292])^(a[404] & b[293])^(a[403] & b[294])^(a[402] & b[295])^(a[401] & b[296])^(a[400] & b[297])^(a[399] & b[298])^(a[398] & b[299])^(a[397] & b[300])^(a[396] & b[301])^(a[395] & b[302])^(a[394] & b[303])^(a[393] & b[304])^(a[392] & b[305])^(a[391] & b[306])^(a[390] & b[307])^(a[389] & b[308])^(a[388] & b[309])^(a[387] & b[310])^(a[386] & b[311])^(a[385] & b[312])^(a[384] & b[313])^(a[383] & b[314])^(a[382] & b[315])^(a[381] & b[316])^(a[380] & b[317])^(a[379] & b[318])^(a[378] & b[319])^(a[377] & b[320])^(a[376] & b[321])^(a[375] & b[322])^(a[374] & b[323])^(a[373] & b[324])^(a[372] & b[325])^(a[371] & b[326])^(a[370] & b[327])^(a[369] & b[328])^(a[368] & b[329])^(a[367] & b[330])^(a[366] & b[331])^(a[365] & b[332])^(a[364] & b[333])^(a[363] & b[334])^(a[362] & b[335])^(a[361] & b[336])^(a[360] & b[337])^(a[359] & b[338])^(a[358] & b[339])^(a[357] & b[340])^(a[356] & b[341])^(a[355] & b[342])^(a[354] & b[343])^(a[353] & b[344])^(a[352] & b[345])^(a[351] & b[346])^(a[350] & b[347])^(a[349] & b[348])^(a[348] & b[349])^(a[347] & b[350])^(a[346] & b[351])^(a[345] & b[352])^(a[344] & b[353])^(a[343] & b[354])^(a[342] & b[355])^(a[341] & b[356])^(a[340] & b[357])^(a[339] & b[358])^(a[338] & b[359])^(a[337] & b[360])^(a[336] & b[361])^(a[335] & b[362])^(a[334] & b[363])^(a[333] & b[364])^(a[332] & b[365])^(a[331] & b[366])^(a[330] & b[367])^(a[329] & b[368])^(a[328] & b[369])^(a[327] & b[370])^(a[326] & b[371])^(a[325] & b[372])^(a[324] & b[373])^(a[323] & b[374])^(a[322] & b[375])^(a[321] & b[376])^(a[320] & b[377])^(a[319] & b[378])^(a[318] & b[379])^(a[317] & b[380])^(a[316] & b[381])^(a[315] & b[382])^(a[314] & b[383])^(a[313] & b[384])^(a[312] & b[385])^(a[311] & b[386])^(a[310] & b[387])^(a[309] & b[388])^(a[308] & b[389])^(a[307] & b[390])^(a[306] & b[391])^(a[305] & b[392])^(a[304] & b[393])^(a[303] & b[394])^(a[302] & b[395])^(a[301] & b[396])^(a[300] & b[397])^(a[299] & b[398])^(a[298] & b[399])^(a[297] & b[400])^(a[296] & b[401])^(a[295] & b[402])^(a[294] & b[403])^(a[293] & b[404])^(a[292] & b[405])^(a[291] & b[406])^(a[290] & b[407])^(a[289] & b[408]);
assign y[698] = (a[408] & b[290])^(a[407] & b[291])^(a[406] & b[292])^(a[405] & b[293])^(a[404] & b[294])^(a[403] & b[295])^(a[402] & b[296])^(a[401] & b[297])^(a[400] & b[298])^(a[399] & b[299])^(a[398] & b[300])^(a[397] & b[301])^(a[396] & b[302])^(a[395] & b[303])^(a[394] & b[304])^(a[393] & b[305])^(a[392] & b[306])^(a[391] & b[307])^(a[390] & b[308])^(a[389] & b[309])^(a[388] & b[310])^(a[387] & b[311])^(a[386] & b[312])^(a[385] & b[313])^(a[384] & b[314])^(a[383] & b[315])^(a[382] & b[316])^(a[381] & b[317])^(a[380] & b[318])^(a[379] & b[319])^(a[378] & b[320])^(a[377] & b[321])^(a[376] & b[322])^(a[375] & b[323])^(a[374] & b[324])^(a[373] & b[325])^(a[372] & b[326])^(a[371] & b[327])^(a[370] & b[328])^(a[369] & b[329])^(a[368] & b[330])^(a[367] & b[331])^(a[366] & b[332])^(a[365] & b[333])^(a[364] & b[334])^(a[363] & b[335])^(a[362] & b[336])^(a[361] & b[337])^(a[360] & b[338])^(a[359] & b[339])^(a[358] & b[340])^(a[357] & b[341])^(a[356] & b[342])^(a[355] & b[343])^(a[354] & b[344])^(a[353] & b[345])^(a[352] & b[346])^(a[351] & b[347])^(a[350] & b[348])^(a[349] & b[349])^(a[348] & b[350])^(a[347] & b[351])^(a[346] & b[352])^(a[345] & b[353])^(a[344] & b[354])^(a[343] & b[355])^(a[342] & b[356])^(a[341] & b[357])^(a[340] & b[358])^(a[339] & b[359])^(a[338] & b[360])^(a[337] & b[361])^(a[336] & b[362])^(a[335] & b[363])^(a[334] & b[364])^(a[333] & b[365])^(a[332] & b[366])^(a[331] & b[367])^(a[330] & b[368])^(a[329] & b[369])^(a[328] & b[370])^(a[327] & b[371])^(a[326] & b[372])^(a[325] & b[373])^(a[324] & b[374])^(a[323] & b[375])^(a[322] & b[376])^(a[321] & b[377])^(a[320] & b[378])^(a[319] & b[379])^(a[318] & b[380])^(a[317] & b[381])^(a[316] & b[382])^(a[315] & b[383])^(a[314] & b[384])^(a[313] & b[385])^(a[312] & b[386])^(a[311] & b[387])^(a[310] & b[388])^(a[309] & b[389])^(a[308] & b[390])^(a[307] & b[391])^(a[306] & b[392])^(a[305] & b[393])^(a[304] & b[394])^(a[303] & b[395])^(a[302] & b[396])^(a[301] & b[397])^(a[300] & b[398])^(a[299] & b[399])^(a[298] & b[400])^(a[297] & b[401])^(a[296] & b[402])^(a[295] & b[403])^(a[294] & b[404])^(a[293] & b[405])^(a[292] & b[406])^(a[291] & b[407])^(a[290] & b[408]);
assign y[699] = (a[408] & b[291])^(a[407] & b[292])^(a[406] & b[293])^(a[405] & b[294])^(a[404] & b[295])^(a[403] & b[296])^(a[402] & b[297])^(a[401] & b[298])^(a[400] & b[299])^(a[399] & b[300])^(a[398] & b[301])^(a[397] & b[302])^(a[396] & b[303])^(a[395] & b[304])^(a[394] & b[305])^(a[393] & b[306])^(a[392] & b[307])^(a[391] & b[308])^(a[390] & b[309])^(a[389] & b[310])^(a[388] & b[311])^(a[387] & b[312])^(a[386] & b[313])^(a[385] & b[314])^(a[384] & b[315])^(a[383] & b[316])^(a[382] & b[317])^(a[381] & b[318])^(a[380] & b[319])^(a[379] & b[320])^(a[378] & b[321])^(a[377] & b[322])^(a[376] & b[323])^(a[375] & b[324])^(a[374] & b[325])^(a[373] & b[326])^(a[372] & b[327])^(a[371] & b[328])^(a[370] & b[329])^(a[369] & b[330])^(a[368] & b[331])^(a[367] & b[332])^(a[366] & b[333])^(a[365] & b[334])^(a[364] & b[335])^(a[363] & b[336])^(a[362] & b[337])^(a[361] & b[338])^(a[360] & b[339])^(a[359] & b[340])^(a[358] & b[341])^(a[357] & b[342])^(a[356] & b[343])^(a[355] & b[344])^(a[354] & b[345])^(a[353] & b[346])^(a[352] & b[347])^(a[351] & b[348])^(a[350] & b[349])^(a[349] & b[350])^(a[348] & b[351])^(a[347] & b[352])^(a[346] & b[353])^(a[345] & b[354])^(a[344] & b[355])^(a[343] & b[356])^(a[342] & b[357])^(a[341] & b[358])^(a[340] & b[359])^(a[339] & b[360])^(a[338] & b[361])^(a[337] & b[362])^(a[336] & b[363])^(a[335] & b[364])^(a[334] & b[365])^(a[333] & b[366])^(a[332] & b[367])^(a[331] & b[368])^(a[330] & b[369])^(a[329] & b[370])^(a[328] & b[371])^(a[327] & b[372])^(a[326] & b[373])^(a[325] & b[374])^(a[324] & b[375])^(a[323] & b[376])^(a[322] & b[377])^(a[321] & b[378])^(a[320] & b[379])^(a[319] & b[380])^(a[318] & b[381])^(a[317] & b[382])^(a[316] & b[383])^(a[315] & b[384])^(a[314] & b[385])^(a[313] & b[386])^(a[312] & b[387])^(a[311] & b[388])^(a[310] & b[389])^(a[309] & b[390])^(a[308] & b[391])^(a[307] & b[392])^(a[306] & b[393])^(a[305] & b[394])^(a[304] & b[395])^(a[303] & b[396])^(a[302] & b[397])^(a[301] & b[398])^(a[300] & b[399])^(a[299] & b[400])^(a[298] & b[401])^(a[297] & b[402])^(a[296] & b[403])^(a[295] & b[404])^(a[294] & b[405])^(a[293] & b[406])^(a[292] & b[407])^(a[291] & b[408]);
assign y[700] = (a[408] & b[292])^(a[407] & b[293])^(a[406] & b[294])^(a[405] & b[295])^(a[404] & b[296])^(a[403] & b[297])^(a[402] & b[298])^(a[401] & b[299])^(a[400] & b[300])^(a[399] & b[301])^(a[398] & b[302])^(a[397] & b[303])^(a[396] & b[304])^(a[395] & b[305])^(a[394] & b[306])^(a[393] & b[307])^(a[392] & b[308])^(a[391] & b[309])^(a[390] & b[310])^(a[389] & b[311])^(a[388] & b[312])^(a[387] & b[313])^(a[386] & b[314])^(a[385] & b[315])^(a[384] & b[316])^(a[383] & b[317])^(a[382] & b[318])^(a[381] & b[319])^(a[380] & b[320])^(a[379] & b[321])^(a[378] & b[322])^(a[377] & b[323])^(a[376] & b[324])^(a[375] & b[325])^(a[374] & b[326])^(a[373] & b[327])^(a[372] & b[328])^(a[371] & b[329])^(a[370] & b[330])^(a[369] & b[331])^(a[368] & b[332])^(a[367] & b[333])^(a[366] & b[334])^(a[365] & b[335])^(a[364] & b[336])^(a[363] & b[337])^(a[362] & b[338])^(a[361] & b[339])^(a[360] & b[340])^(a[359] & b[341])^(a[358] & b[342])^(a[357] & b[343])^(a[356] & b[344])^(a[355] & b[345])^(a[354] & b[346])^(a[353] & b[347])^(a[352] & b[348])^(a[351] & b[349])^(a[350] & b[350])^(a[349] & b[351])^(a[348] & b[352])^(a[347] & b[353])^(a[346] & b[354])^(a[345] & b[355])^(a[344] & b[356])^(a[343] & b[357])^(a[342] & b[358])^(a[341] & b[359])^(a[340] & b[360])^(a[339] & b[361])^(a[338] & b[362])^(a[337] & b[363])^(a[336] & b[364])^(a[335] & b[365])^(a[334] & b[366])^(a[333] & b[367])^(a[332] & b[368])^(a[331] & b[369])^(a[330] & b[370])^(a[329] & b[371])^(a[328] & b[372])^(a[327] & b[373])^(a[326] & b[374])^(a[325] & b[375])^(a[324] & b[376])^(a[323] & b[377])^(a[322] & b[378])^(a[321] & b[379])^(a[320] & b[380])^(a[319] & b[381])^(a[318] & b[382])^(a[317] & b[383])^(a[316] & b[384])^(a[315] & b[385])^(a[314] & b[386])^(a[313] & b[387])^(a[312] & b[388])^(a[311] & b[389])^(a[310] & b[390])^(a[309] & b[391])^(a[308] & b[392])^(a[307] & b[393])^(a[306] & b[394])^(a[305] & b[395])^(a[304] & b[396])^(a[303] & b[397])^(a[302] & b[398])^(a[301] & b[399])^(a[300] & b[400])^(a[299] & b[401])^(a[298] & b[402])^(a[297] & b[403])^(a[296] & b[404])^(a[295] & b[405])^(a[294] & b[406])^(a[293] & b[407])^(a[292] & b[408]);
assign y[701] = (a[408] & b[293])^(a[407] & b[294])^(a[406] & b[295])^(a[405] & b[296])^(a[404] & b[297])^(a[403] & b[298])^(a[402] & b[299])^(a[401] & b[300])^(a[400] & b[301])^(a[399] & b[302])^(a[398] & b[303])^(a[397] & b[304])^(a[396] & b[305])^(a[395] & b[306])^(a[394] & b[307])^(a[393] & b[308])^(a[392] & b[309])^(a[391] & b[310])^(a[390] & b[311])^(a[389] & b[312])^(a[388] & b[313])^(a[387] & b[314])^(a[386] & b[315])^(a[385] & b[316])^(a[384] & b[317])^(a[383] & b[318])^(a[382] & b[319])^(a[381] & b[320])^(a[380] & b[321])^(a[379] & b[322])^(a[378] & b[323])^(a[377] & b[324])^(a[376] & b[325])^(a[375] & b[326])^(a[374] & b[327])^(a[373] & b[328])^(a[372] & b[329])^(a[371] & b[330])^(a[370] & b[331])^(a[369] & b[332])^(a[368] & b[333])^(a[367] & b[334])^(a[366] & b[335])^(a[365] & b[336])^(a[364] & b[337])^(a[363] & b[338])^(a[362] & b[339])^(a[361] & b[340])^(a[360] & b[341])^(a[359] & b[342])^(a[358] & b[343])^(a[357] & b[344])^(a[356] & b[345])^(a[355] & b[346])^(a[354] & b[347])^(a[353] & b[348])^(a[352] & b[349])^(a[351] & b[350])^(a[350] & b[351])^(a[349] & b[352])^(a[348] & b[353])^(a[347] & b[354])^(a[346] & b[355])^(a[345] & b[356])^(a[344] & b[357])^(a[343] & b[358])^(a[342] & b[359])^(a[341] & b[360])^(a[340] & b[361])^(a[339] & b[362])^(a[338] & b[363])^(a[337] & b[364])^(a[336] & b[365])^(a[335] & b[366])^(a[334] & b[367])^(a[333] & b[368])^(a[332] & b[369])^(a[331] & b[370])^(a[330] & b[371])^(a[329] & b[372])^(a[328] & b[373])^(a[327] & b[374])^(a[326] & b[375])^(a[325] & b[376])^(a[324] & b[377])^(a[323] & b[378])^(a[322] & b[379])^(a[321] & b[380])^(a[320] & b[381])^(a[319] & b[382])^(a[318] & b[383])^(a[317] & b[384])^(a[316] & b[385])^(a[315] & b[386])^(a[314] & b[387])^(a[313] & b[388])^(a[312] & b[389])^(a[311] & b[390])^(a[310] & b[391])^(a[309] & b[392])^(a[308] & b[393])^(a[307] & b[394])^(a[306] & b[395])^(a[305] & b[396])^(a[304] & b[397])^(a[303] & b[398])^(a[302] & b[399])^(a[301] & b[400])^(a[300] & b[401])^(a[299] & b[402])^(a[298] & b[403])^(a[297] & b[404])^(a[296] & b[405])^(a[295] & b[406])^(a[294] & b[407])^(a[293] & b[408]);
assign y[702] = (a[408] & b[294])^(a[407] & b[295])^(a[406] & b[296])^(a[405] & b[297])^(a[404] & b[298])^(a[403] & b[299])^(a[402] & b[300])^(a[401] & b[301])^(a[400] & b[302])^(a[399] & b[303])^(a[398] & b[304])^(a[397] & b[305])^(a[396] & b[306])^(a[395] & b[307])^(a[394] & b[308])^(a[393] & b[309])^(a[392] & b[310])^(a[391] & b[311])^(a[390] & b[312])^(a[389] & b[313])^(a[388] & b[314])^(a[387] & b[315])^(a[386] & b[316])^(a[385] & b[317])^(a[384] & b[318])^(a[383] & b[319])^(a[382] & b[320])^(a[381] & b[321])^(a[380] & b[322])^(a[379] & b[323])^(a[378] & b[324])^(a[377] & b[325])^(a[376] & b[326])^(a[375] & b[327])^(a[374] & b[328])^(a[373] & b[329])^(a[372] & b[330])^(a[371] & b[331])^(a[370] & b[332])^(a[369] & b[333])^(a[368] & b[334])^(a[367] & b[335])^(a[366] & b[336])^(a[365] & b[337])^(a[364] & b[338])^(a[363] & b[339])^(a[362] & b[340])^(a[361] & b[341])^(a[360] & b[342])^(a[359] & b[343])^(a[358] & b[344])^(a[357] & b[345])^(a[356] & b[346])^(a[355] & b[347])^(a[354] & b[348])^(a[353] & b[349])^(a[352] & b[350])^(a[351] & b[351])^(a[350] & b[352])^(a[349] & b[353])^(a[348] & b[354])^(a[347] & b[355])^(a[346] & b[356])^(a[345] & b[357])^(a[344] & b[358])^(a[343] & b[359])^(a[342] & b[360])^(a[341] & b[361])^(a[340] & b[362])^(a[339] & b[363])^(a[338] & b[364])^(a[337] & b[365])^(a[336] & b[366])^(a[335] & b[367])^(a[334] & b[368])^(a[333] & b[369])^(a[332] & b[370])^(a[331] & b[371])^(a[330] & b[372])^(a[329] & b[373])^(a[328] & b[374])^(a[327] & b[375])^(a[326] & b[376])^(a[325] & b[377])^(a[324] & b[378])^(a[323] & b[379])^(a[322] & b[380])^(a[321] & b[381])^(a[320] & b[382])^(a[319] & b[383])^(a[318] & b[384])^(a[317] & b[385])^(a[316] & b[386])^(a[315] & b[387])^(a[314] & b[388])^(a[313] & b[389])^(a[312] & b[390])^(a[311] & b[391])^(a[310] & b[392])^(a[309] & b[393])^(a[308] & b[394])^(a[307] & b[395])^(a[306] & b[396])^(a[305] & b[397])^(a[304] & b[398])^(a[303] & b[399])^(a[302] & b[400])^(a[301] & b[401])^(a[300] & b[402])^(a[299] & b[403])^(a[298] & b[404])^(a[297] & b[405])^(a[296] & b[406])^(a[295] & b[407])^(a[294] & b[408]);
assign y[703] = (a[408] & b[295])^(a[407] & b[296])^(a[406] & b[297])^(a[405] & b[298])^(a[404] & b[299])^(a[403] & b[300])^(a[402] & b[301])^(a[401] & b[302])^(a[400] & b[303])^(a[399] & b[304])^(a[398] & b[305])^(a[397] & b[306])^(a[396] & b[307])^(a[395] & b[308])^(a[394] & b[309])^(a[393] & b[310])^(a[392] & b[311])^(a[391] & b[312])^(a[390] & b[313])^(a[389] & b[314])^(a[388] & b[315])^(a[387] & b[316])^(a[386] & b[317])^(a[385] & b[318])^(a[384] & b[319])^(a[383] & b[320])^(a[382] & b[321])^(a[381] & b[322])^(a[380] & b[323])^(a[379] & b[324])^(a[378] & b[325])^(a[377] & b[326])^(a[376] & b[327])^(a[375] & b[328])^(a[374] & b[329])^(a[373] & b[330])^(a[372] & b[331])^(a[371] & b[332])^(a[370] & b[333])^(a[369] & b[334])^(a[368] & b[335])^(a[367] & b[336])^(a[366] & b[337])^(a[365] & b[338])^(a[364] & b[339])^(a[363] & b[340])^(a[362] & b[341])^(a[361] & b[342])^(a[360] & b[343])^(a[359] & b[344])^(a[358] & b[345])^(a[357] & b[346])^(a[356] & b[347])^(a[355] & b[348])^(a[354] & b[349])^(a[353] & b[350])^(a[352] & b[351])^(a[351] & b[352])^(a[350] & b[353])^(a[349] & b[354])^(a[348] & b[355])^(a[347] & b[356])^(a[346] & b[357])^(a[345] & b[358])^(a[344] & b[359])^(a[343] & b[360])^(a[342] & b[361])^(a[341] & b[362])^(a[340] & b[363])^(a[339] & b[364])^(a[338] & b[365])^(a[337] & b[366])^(a[336] & b[367])^(a[335] & b[368])^(a[334] & b[369])^(a[333] & b[370])^(a[332] & b[371])^(a[331] & b[372])^(a[330] & b[373])^(a[329] & b[374])^(a[328] & b[375])^(a[327] & b[376])^(a[326] & b[377])^(a[325] & b[378])^(a[324] & b[379])^(a[323] & b[380])^(a[322] & b[381])^(a[321] & b[382])^(a[320] & b[383])^(a[319] & b[384])^(a[318] & b[385])^(a[317] & b[386])^(a[316] & b[387])^(a[315] & b[388])^(a[314] & b[389])^(a[313] & b[390])^(a[312] & b[391])^(a[311] & b[392])^(a[310] & b[393])^(a[309] & b[394])^(a[308] & b[395])^(a[307] & b[396])^(a[306] & b[397])^(a[305] & b[398])^(a[304] & b[399])^(a[303] & b[400])^(a[302] & b[401])^(a[301] & b[402])^(a[300] & b[403])^(a[299] & b[404])^(a[298] & b[405])^(a[297] & b[406])^(a[296] & b[407])^(a[295] & b[408]);
assign y[704] = (a[408] & b[296])^(a[407] & b[297])^(a[406] & b[298])^(a[405] & b[299])^(a[404] & b[300])^(a[403] & b[301])^(a[402] & b[302])^(a[401] & b[303])^(a[400] & b[304])^(a[399] & b[305])^(a[398] & b[306])^(a[397] & b[307])^(a[396] & b[308])^(a[395] & b[309])^(a[394] & b[310])^(a[393] & b[311])^(a[392] & b[312])^(a[391] & b[313])^(a[390] & b[314])^(a[389] & b[315])^(a[388] & b[316])^(a[387] & b[317])^(a[386] & b[318])^(a[385] & b[319])^(a[384] & b[320])^(a[383] & b[321])^(a[382] & b[322])^(a[381] & b[323])^(a[380] & b[324])^(a[379] & b[325])^(a[378] & b[326])^(a[377] & b[327])^(a[376] & b[328])^(a[375] & b[329])^(a[374] & b[330])^(a[373] & b[331])^(a[372] & b[332])^(a[371] & b[333])^(a[370] & b[334])^(a[369] & b[335])^(a[368] & b[336])^(a[367] & b[337])^(a[366] & b[338])^(a[365] & b[339])^(a[364] & b[340])^(a[363] & b[341])^(a[362] & b[342])^(a[361] & b[343])^(a[360] & b[344])^(a[359] & b[345])^(a[358] & b[346])^(a[357] & b[347])^(a[356] & b[348])^(a[355] & b[349])^(a[354] & b[350])^(a[353] & b[351])^(a[352] & b[352])^(a[351] & b[353])^(a[350] & b[354])^(a[349] & b[355])^(a[348] & b[356])^(a[347] & b[357])^(a[346] & b[358])^(a[345] & b[359])^(a[344] & b[360])^(a[343] & b[361])^(a[342] & b[362])^(a[341] & b[363])^(a[340] & b[364])^(a[339] & b[365])^(a[338] & b[366])^(a[337] & b[367])^(a[336] & b[368])^(a[335] & b[369])^(a[334] & b[370])^(a[333] & b[371])^(a[332] & b[372])^(a[331] & b[373])^(a[330] & b[374])^(a[329] & b[375])^(a[328] & b[376])^(a[327] & b[377])^(a[326] & b[378])^(a[325] & b[379])^(a[324] & b[380])^(a[323] & b[381])^(a[322] & b[382])^(a[321] & b[383])^(a[320] & b[384])^(a[319] & b[385])^(a[318] & b[386])^(a[317] & b[387])^(a[316] & b[388])^(a[315] & b[389])^(a[314] & b[390])^(a[313] & b[391])^(a[312] & b[392])^(a[311] & b[393])^(a[310] & b[394])^(a[309] & b[395])^(a[308] & b[396])^(a[307] & b[397])^(a[306] & b[398])^(a[305] & b[399])^(a[304] & b[400])^(a[303] & b[401])^(a[302] & b[402])^(a[301] & b[403])^(a[300] & b[404])^(a[299] & b[405])^(a[298] & b[406])^(a[297] & b[407])^(a[296] & b[408]);
assign y[705] = (a[408] & b[297])^(a[407] & b[298])^(a[406] & b[299])^(a[405] & b[300])^(a[404] & b[301])^(a[403] & b[302])^(a[402] & b[303])^(a[401] & b[304])^(a[400] & b[305])^(a[399] & b[306])^(a[398] & b[307])^(a[397] & b[308])^(a[396] & b[309])^(a[395] & b[310])^(a[394] & b[311])^(a[393] & b[312])^(a[392] & b[313])^(a[391] & b[314])^(a[390] & b[315])^(a[389] & b[316])^(a[388] & b[317])^(a[387] & b[318])^(a[386] & b[319])^(a[385] & b[320])^(a[384] & b[321])^(a[383] & b[322])^(a[382] & b[323])^(a[381] & b[324])^(a[380] & b[325])^(a[379] & b[326])^(a[378] & b[327])^(a[377] & b[328])^(a[376] & b[329])^(a[375] & b[330])^(a[374] & b[331])^(a[373] & b[332])^(a[372] & b[333])^(a[371] & b[334])^(a[370] & b[335])^(a[369] & b[336])^(a[368] & b[337])^(a[367] & b[338])^(a[366] & b[339])^(a[365] & b[340])^(a[364] & b[341])^(a[363] & b[342])^(a[362] & b[343])^(a[361] & b[344])^(a[360] & b[345])^(a[359] & b[346])^(a[358] & b[347])^(a[357] & b[348])^(a[356] & b[349])^(a[355] & b[350])^(a[354] & b[351])^(a[353] & b[352])^(a[352] & b[353])^(a[351] & b[354])^(a[350] & b[355])^(a[349] & b[356])^(a[348] & b[357])^(a[347] & b[358])^(a[346] & b[359])^(a[345] & b[360])^(a[344] & b[361])^(a[343] & b[362])^(a[342] & b[363])^(a[341] & b[364])^(a[340] & b[365])^(a[339] & b[366])^(a[338] & b[367])^(a[337] & b[368])^(a[336] & b[369])^(a[335] & b[370])^(a[334] & b[371])^(a[333] & b[372])^(a[332] & b[373])^(a[331] & b[374])^(a[330] & b[375])^(a[329] & b[376])^(a[328] & b[377])^(a[327] & b[378])^(a[326] & b[379])^(a[325] & b[380])^(a[324] & b[381])^(a[323] & b[382])^(a[322] & b[383])^(a[321] & b[384])^(a[320] & b[385])^(a[319] & b[386])^(a[318] & b[387])^(a[317] & b[388])^(a[316] & b[389])^(a[315] & b[390])^(a[314] & b[391])^(a[313] & b[392])^(a[312] & b[393])^(a[311] & b[394])^(a[310] & b[395])^(a[309] & b[396])^(a[308] & b[397])^(a[307] & b[398])^(a[306] & b[399])^(a[305] & b[400])^(a[304] & b[401])^(a[303] & b[402])^(a[302] & b[403])^(a[301] & b[404])^(a[300] & b[405])^(a[299] & b[406])^(a[298] & b[407])^(a[297] & b[408]);
assign y[706] = (a[408] & b[298])^(a[407] & b[299])^(a[406] & b[300])^(a[405] & b[301])^(a[404] & b[302])^(a[403] & b[303])^(a[402] & b[304])^(a[401] & b[305])^(a[400] & b[306])^(a[399] & b[307])^(a[398] & b[308])^(a[397] & b[309])^(a[396] & b[310])^(a[395] & b[311])^(a[394] & b[312])^(a[393] & b[313])^(a[392] & b[314])^(a[391] & b[315])^(a[390] & b[316])^(a[389] & b[317])^(a[388] & b[318])^(a[387] & b[319])^(a[386] & b[320])^(a[385] & b[321])^(a[384] & b[322])^(a[383] & b[323])^(a[382] & b[324])^(a[381] & b[325])^(a[380] & b[326])^(a[379] & b[327])^(a[378] & b[328])^(a[377] & b[329])^(a[376] & b[330])^(a[375] & b[331])^(a[374] & b[332])^(a[373] & b[333])^(a[372] & b[334])^(a[371] & b[335])^(a[370] & b[336])^(a[369] & b[337])^(a[368] & b[338])^(a[367] & b[339])^(a[366] & b[340])^(a[365] & b[341])^(a[364] & b[342])^(a[363] & b[343])^(a[362] & b[344])^(a[361] & b[345])^(a[360] & b[346])^(a[359] & b[347])^(a[358] & b[348])^(a[357] & b[349])^(a[356] & b[350])^(a[355] & b[351])^(a[354] & b[352])^(a[353] & b[353])^(a[352] & b[354])^(a[351] & b[355])^(a[350] & b[356])^(a[349] & b[357])^(a[348] & b[358])^(a[347] & b[359])^(a[346] & b[360])^(a[345] & b[361])^(a[344] & b[362])^(a[343] & b[363])^(a[342] & b[364])^(a[341] & b[365])^(a[340] & b[366])^(a[339] & b[367])^(a[338] & b[368])^(a[337] & b[369])^(a[336] & b[370])^(a[335] & b[371])^(a[334] & b[372])^(a[333] & b[373])^(a[332] & b[374])^(a[331] & b[375])^(a[330] & b[376])^(a[329] & b[377])^(a[328] & b[378])^(a[327] & b[379])^(a[326] & b[380])^(a[325] & b[381])^(a[324] & b[382])^(a[323] & b[383])^(a[322] & b[384])^(a[321] & b[385])^(a[320] & b[386])^(a[319] & b[387])^(a[318] & b[388])^(a[317] & b[389])^(a[316] & b[390])^(a[315] & b[391])^(a[314] & b[392])^(a[313] & b[393])^(a[312] & b[394])^(a[311] & b[395])^(a[310] & b[396])^(a[309] & b[397])^(a[308] & b[398])^(a[307] & b[399])^(a[306] & b[400])^(a[305] & b[401])^(a[304] & b[402])^(a[303] & b[403])^(a[302] & b[404])^(a[301] & b[405])^(a[300] & b[406])^(a[299] & b[407])^(a[298] & b[408]);
assign y[707] = (a[408] & b[299])^(a[407] & b[300])^(a[406] & b[301])^(a[405] & b[302])^(a[404] & b[303])^(a[403] & b[304])^(a[402] & b[305])^(a[401] & b[306])^(a[400] & b[307])^(a[399] & b[308])^(a[398] & b[309])^(a[397] & b[310])^(a[396] & b[311])^(a[395] & b[312])^(a[394] & b[313])^(a[393] & b[314])^(a[392] & b[315])^(a[391] & b[316])^(a[390] & b[317])^(a[389] & b[318])^(a[388] & b[319])^(a[387] & b[320])^(a[386] & b[321])^(a[385] & b[322])^(a[384] & b[323])^(a[383] & b[324])^(a[382] & b[325])^(a[381] & b[326])^(a[380] & b[327])^(a[379] & b[328])^(a[378] & b[329])^(a[377] & b[330])^(a[376] & b[331])^(a[375] & b[332])^(a[374] & b[333])^(a[373] & b[334])^(a[372] & b[335])^(a[371] & b[336])^(a[370] & b[337])^(a[369] & b[338])^(a[368] & b[339])^(a[367] & b[340])^(a[366] & b[341])^(a[365] & b[342])^(a[364] & b[343])^(a[363] & b[344])^(a[362] & b[345])^(a[361] & b[346])^(a[360] & b[347])^(a[359] & b[348])^(a[358] & b[349])^(a[357] & b[350])^(a[356] & b[351])^(a[355] & b[352])^(a[354] & b[353])^(a[353] & b[354])^(a[352] & b[355])^(a[351] & b[356])^(a[350] & b[357])^(a[349] & b[358])^(a[348] & b[359])^(a[347] & b[360])^(a[346] & b[361])^(a[345] & b[362])^(a[344] & b[363])^(a[343] & b[364])^(a[342] & b[365])^(a[341] & b[366])^(a[340] & b[367])^(a[339] & b[368])^(a[338] & b[369])^(a[337] & b[370])^(a[336] & b[371])^(a[335] & b[372])^(a[334] & b[373])^(a[333] & b[374])^(a[332] & b[375])^(a[331] & b[376])^(a[330] & b[377])^(a[329] & b[378])^(a[328] & b[379])^(a[327] & b[380])^(a[326] & b[381])^(a[325] & b[382])^(a[324] & b[383])^(a[323] & b[384])^(a[322] & b[385])^(a[321] & b[386])^(a[320] & b[387])^(a[319] & b[388])^(a[318] & b[389])^(a[317] & b[390])^(a[316] & b[391])^(a[315] & b[392])^(a[314] & b[393])^(a[313] & b[394])^(a[312] & b[395])^(a[311] & b[396])^(a[310] & b[397])^(a[309] & b[398])^(a[308] & b[399])^(a[307] & b[400])^(a[306] & b[401])^(a[305] & b[402])^(a[304] & b[403])^(a[303] & b[404])^(a[302] & b[405])^(a[301] & b[406])^(a[300] & b[407])^(a[299] & b[408]);
assign y[708] = (a[408] & b[300])^(a[407] & b[301])^(a[406] & b[302])^(a[405] & b[303])^(a[404] & b[304])^(a[403] & b[305])^(a[402] & b[306])^(a[401] & b[307])^(a[400] & b[308])^(a[399] & b[309])^(a[398] & b[310])^(a[397] & b[311])^(a[396] & b[312])^(a[395] & b[313])^(a[394] & b[314])^(a[393] & b[315])^(a[392] & b[316])^(a[391] & b[317])^(a[390] & b[318])^(a[389] & b[319])^(a[388] & b[320])^(a[387] & b[321])^(a[386] & b[322])^(a[385] & b[323])^(a[384] & b[324])^(a[383] & b[325])^(a[382] & b[326])^(a[381] & b[327])^(a[380] & b[328])^(a[379] & b[329])^(a[378] & b[330])^(a[377] & b[331])^(a[376] & b[332])^(a[375] & b[333])^(a[374] & b[334])^(a[373] & b[335])^(a[372] & b[336])^(a[371] & b[337])^(a[370] & b[338])^(a[369] & b[339])^(a[368] & b[340])^(a[367] & b[341])^(a[366] & b[342])^(a[365] & b[343])^(a[364] & b[344])^(a[363] & b[345])^(a[362] & b[346])^(a[361] & b[347])^(a[360] & b[348])^(a[359] & b[349])^(a[358] & b[350])^(a[357] & b[351])^(a[356] & b[352])^(a[355] & b[353])^(a[354] & b[354])^(a[353] & b[355])^(a[352] & b[356])^(a[351] & b[357])^(a[350] & b[358])^(a[349] & b[359])^(a[348] & b[360])^(a[347] & b[361])^(a[346] & b[362])^(a[345] & b[363])^(a[344] & b[364])^(a[343] & b[365])^(a[342] & b[366])^(a[341] & b[367])^(a[340] & b[368])^(a[339] & b[369])^(a[338] & b[370])^(a[337] & b[371])^(a[336] & b[372])^(a[335] & b[373])^(a[334] & b[374])^(a[333] & b[375])^(a[332] & b[376])^(a[331] & b[377])^(a[330] & b[378])^(a[329] & b[379])^(a[328] & b[380])^(a[327] & b[381])^(a[326] & b[382])^(a[325] & b[383])^(a[324] & b[384])^(a[323] & b[385])^(a[322] & b[386])^(a[321] & b[387])^(a[320] & b[388])^(a[319] & b[389])^(a[318] & b[390])^(a[317] & b[391])^(a[316] & b[392])^(a[315] & b[393])^(a[314] & b[394])^(a[313] & b[395])^(a[312] & b[396])^(a[311] & b[397])^(a[310] & b[398])^(a[309] & b[399])^(a[308] & b[400])^(a[307] & b[401])^(a[306] & b[402])^(a[305] & b[403])^(a[304] & b[404])^(a[303] & b[405])^(a[302] & b[406])^(a[301] & b[407])^(a[300] & b[408]);
assign y[709] = (a[408] & b[301])^(a[407] & b[302])^(a[406] & b[303])^(a[405] & b[304])^(a[404] & b[305])^(a[403] & b[306])^(a[402] & b[307])^(a[401] & b[308])^(a[400] & b[309])^(a[399] & b[310])^(a[398] & b[311])^(a[397] & b[312])^(a[396] & b[313])^(a[395] & b[314])^(a[394] & b[315])^(a[393] & b[316])^(a[392] & b[317])^(a[391] & b[318])^(a[390] & b[319])^(a[389] & b[320])^(a[388] & b[321])^(a[387] & b[322])^(a[386] & b[323])^(a[385] & b[324])^(a[384] & b[325])^(a[383] & b[326])^(a[382] & b[327])^(a[381] & b[328])^(a[380] & b[329])^(a[379] & b[330])^(a[378] & b[331])^(a[377] & b[332])^(a[376] & b[333])^(a[375] & b[334])^(a[374] & b[335])^(a[373] & b[336])^(a[372] & b[337])^(a[371] & b[338])^(a[370] & b[339])^(a[369] & b[340])^(a[368] & b[341])^(a[367] & b[342])^(a[366] & b[343])^(a[365] & b[344])^(a[364] & b[345])^(a[363] & b[346])^(a[362] & b[347])^(a[361] & b[348])^(a[360] & b[349])^(a[359] & b[350])^(a[358] & b[351])^(a[357] & b[352])^(a[356] & b[353])^(a[355] & b[354])^(a[354] & b[355])^(a[353] & b[356])^(a[352] & b[357])^(a[351] & b[358])^(a[350] & b[359])^(a[349] & b[360])^(a[348] & b[361])^(a[347] & b[362])^(a[346] & b[363])^(a[345] & b[364])^(a[344] & b[365])^(a[343] & b[366])^(a[342] & b[367])^(a[341] & b[368])^(a[340] & b[369])^(a[339] & b[370])^(a[338] & b[371])^(a[337] & b[372])^(a[336] & b[373])^(a[335] & b[374])^(a[334] & b[375])^(a[333] & b[376])^(a[332] & b[377])^(a[331] & b[378])^(a[330] & b[379])^(a[329] & b[380])^(a[328] & b[381])^(a[327] & b[382])^(a[326] & b[383])^(a[325] & b[384])^(a[324] & b[385])^(a[323] & b[386])^(a[322] & b[387])^(a[321] & b[388])^(a[320] & b[389])^(a[319] & b[390])^(a[318] & b[391])^(a[317] & b[392])^(a[316] & b[393])^(a[315] & b[394])^(a[314] & b[395])^(a[313] & b[396])^(a[312] & b[397])^(a[311] & b[398])^(a[310] & b[399])^(a[309] & b[400])^(a[308] & b[401])^(a[307] & b[402])^(a[306] & b[403])^(a[305] & b[404])^(a[304] & b[405])^(a[303] & b[406])^(a[302] & b[407])^(a[301] & b[408]);
assign y[710] = (a[408] & b[302])^(a[407] & b[303])^(a[406] & b[304])^(a[405] & b[305])^(a[404] & b[306])^(a[403] & b[307])^(a[402] & b[308])^(a[401] & b[309])^(a[400] & b[310])^(a[399] & b[311])^(a[398] & b[312])^(a[397] & b[313])^(a[396] & b[314])^(a[395] & b[315])^(a[394] & b[316])^(a[393] & b[317])^(a[392] & b[318])^(a[391] & b[319])^(a[390] & b[320])^(a[389] & b[321])^(a[388] & b[322])^(a[387] & b[323])^(a[386] & b[324])^(a[385] & b[325])^(a[384] & b[326])^(a[383] & b[327])^(a[382] & b[328])^(a[381] & b[329])^(a[380] & b[330])^(a[379] & b[331])^(a[378] & b[332])^(a[377] & b[333])^(a[376] & b[334])^(a[375] & b[335])^(a[374] & b[336])^(a[373] & b[337])^(a[372] & b[338])^(a[371] & b[339])^(a[370] & b[340])^(a[369] & b[341])^(a[368] & b[342])^(a[367] & b[343])^(a[366] & b[344])^(a[365] & b[345])^(a[364] & b[346])^(a[363] & b[347])^(a[362] & b[348])^(a[361] & b[349])^(a[360] & b[350])^(a[359] & b[351])^(a[358] & b[352])^(a[357] & b[353])^(a[356] & b[354])^(a[355] & b[355])^(a[354] & b[356])^(a[353] & b[357])^(a[352] & b[358])^(a[351] & b[359])^(a[350] & b[360])^(a[349] & b[361])^(a[348] & b[362])^(a[347] & b[363])^(a[346] & b[364])^(a[345] & b[365])^(a[344] & b[366])^(a[343] & b[367])^(a[342] & b[368])^(a[341] & b[369])^(a[340] & b[370])^(a[339] & b[371])^(a[338] & b[372])^(a[337] & b[373])^(a[336] & b[374])^(a[335] & b[375])^(a[334] & b[376])^(a[333] & b[377])^(a[332] & b[378])^(a[331] & b[379])^(a[330] & b[380])^(a[329] & b[381])^(a[328] & b[382])^(a[327] & b[383])^(a[326] & b[384])^(a[325] & b[385])^(a[324] & b[386])^(a[323] & b[387])^(a[322] & b[388])^(a[321] & b[389])^(a[320] & b[390])^(a[319] & b[391])^(a[318] & b[392])^(a[317] & b[393])^(a[316] & b[394])^(a[315] & b[395])^(a[314] & b[396])^(a[313] & b[397])^(a[312] & b[398])^(a[311] & b[399])^(a[310] & b[400])^(a[309] & b[401])^(a[308] & b[402])^(a[307] & b[403])^(a[306] & b[404])^(a[305] & b[405])^(a[304] & b[406])^(a[303] & b[407])^(a[302] & b[408]);
assign y[711] = (a[408] & b[303])^(a[407] & b[304])^(a[406] & b[305])^(a[405] & b[306])^(a[404] & b[307])^(a[403] & b[308])^(a[402] & b[309])^(a[401] & b[310])^(a[400] & b[311])^(a[399] & b[312])^(a[398] & b[313])^(a[397] & b[314])^(a[396] & b[315])^(a[395] & b[316])^(a[394] & b[317])^(a[393] & b[318])^(a[392] & b[319])^(a[391] & b[320])^(a[390] & b[321])^(a[389] & b[322])^(a[388] & b[323])^(a[387] & b[324])^(a[386] & b[325])^(a[385] & b[326])^(a[384] & b[327])^(a[383] & b[328])^(a[382] & b[329])^(a[381] & b[330])^(a[380] & b[331])^(a[379] & b[332])^(a[378] & b[333])^(a[377] & b[334])^(a[376] & b[335])^(a[375] & b[336])^(a[374] & b[337])^(a[373] & b[338])^(a[372] & b[339])^(a[371] & b[340])^(a[370] & b[341])^(a[369] & b[342])^(a[368] & b[343])^(a[367] & b[344])^(a[366] & b[345])^(a[365] & b[346])^(a[364] & b[347])^(a[363] & b[348])^(a[362] & b[349])^(a[361] & b[350])^(a[360] & b[351])^(a[359] & b[352])^(a[358] & b[353])^(a[357] & b[354])^(a[356] & b[355])^(a[355] & b[356])^(a[354] & b[357])^(a[353] & b[358])^(a[352] & b[359])^(a[351] & b[360])^(a[350] & b[361])^(a[349] & b[362])^(a[348] & b[363])^(a[347] & b[364])^(a[346] & b[365])^(a[345] & b[366])^(a[344] & b[367])^(a[343] & b[368])^(a[342] & b[369])^(a[341] & b[370])^(a[340] & b[371])^(a[339] & b[372])^(a[338] & b[373])^(a[337] & b[374])^(a[336] & b[375])^(a[335] & b[376])^(a[334] & b[377])^(a[333] & b[378])^(a[332] & b[379])^(a[331] & b[380])^(a[330] & b[381])^(a[329] & b[382])^(a[328] & b[383])^(a[327] & b[384])^(a[326] & b[385])^(a[325] & b[386])^(a[324] & b[387])^(a[323] & b[388])^(a[322] & b[389])^(a[321] & b[390])^(a[320] & b[391])^(a[319] & b[392])^(a[318] & b[393])^(a[317] & b[394])^(a[316] & b[395])^(a[315] & b[396])^(a[314] & b[397])^(a[313] & b[398])^(a[312] & b[399])^(a[311] & b[400])^(a[310] & b[401])^(a[309] & b[402])^(a[308] & b[403])^(a[307] & b[404])^(a[306] & b[405])^(a[305] & b[406])^(a[304] & b[407])^(a[303] & b[408]);
assign y[712] = (a[408] & b[304])^(a[407] & b[305])^(a[406] & b[306])^(a[405] & b[307])^(a[404] & b[308])^(a[403] & b[309])^(a[402] & b[310])^(a[401] & b[311])^(a[400] & b[312])^(a[399] & b[313])^(a[398] & b[314])^(a[397] & b[315])^(a[396] & b[316])^(a[395] & b[317])^(a[394] & b[318])^(a[393] & b[319])^(a[392] & b[320])^(a[391] & b[321])^(a[390] & b[322])^(a[389] & b[323])^(a[388] & b[324])^(a[387] & b[325])^(a[386] & b[326])^(a[385] & b[327])^(a[384] & b[328])^(a[383] & b[329])^(a[382] & b[330])^(a[381] & b[331])^(a[380] & b[332])^(a[379] & b[333])^(a[378] & b[334])^(a[377] & b[335])^(a[376] & b[336])^(a[375] & b[337])^(a[374] & b[338])^(a[373] & b[339])^(a[372] & b[340])^(a[371] & b[341])^(a[370] & b[342])^(a[369] & b[343])^(a[368] & b[344])^(a[367] & b[345])^(a[366] & b[346])^(a[365] & b[347])^(a[364] & b[348])^(a[363] & b[349])^(a[362] & b[350])^(a[361] & b[351])^(a[360] & b[352])^(a[359] & b[353])^(a[358] & b[354])^(a[357] & b[355])^(a[356] & b[356])^(a[355] & b[357])^(a[354] & b[358])^(a[353] & b[359])^(a[352] & b[360])^(a[351] & b[361])^(a[350] & b[362])^(a[349] & b[363])^(a[348] & b[364])^(a[347] & b[365])^(a[346] & b[366])^(a[345] & b[367])^(a[344] & b[368])^(a[343] & b[369])^(a[342] & b[370])^(a[341] & b[371])^(a[340] & b[372])^(a[339] & b[373])^(a[338] & b[374])^(a[337] & b[375])^(a[336] & b[376])^(a[335] & b[377])^(a[334] & b[378])^(a[333] & b[379])^(a[332] & b[380])^(a[331] & b[381])^(a[330] & b[382])^(a[329] & b[383])^(a[328] & b[384])^(a[327] & b[385])^(a[326] & b[386])^(a[325] & b[387])^(a[324] & b[388])^(a[323] & b[389])^(a[322] & b[390])^(a[321] & b[391])^(a[320] & b[392])^(a[319] & b[393])^(a[318] & b[394])^(a[317] & b[395])^(a[316] & b[396])^(a[315] & b[397])^(a[314] & b[398])^(a[313] & b[399])^(a[312] & b[400])^(a[311] & b[401])^(a[310] & b[402])^(a[309] & b[403])^(a[308] & b[404])^(a[307] & b[405])^(a[306] & b[406])^(a[305] & b[407])^(a[304] & b[408]);
assign y[713] = (a[408] & b[305])^(a[407] & b[306])^(a[406] & b[307])^(a[405] & b[308])^(a[404] & b[309])^(a[403] & b[310])^(a[402] & b[311])^(a[401] & b[312])^(a[400] & b[313])^(a[399] & b[314])^(a[398] & b[315])^(a[397] & b[316])^(a[396] & b[317])^(a[395] & b[318])^(a[394] & b[319])^(a[393] & b[320])^(a[392] & b[321])^(a[391] & b[322])^(a[390] & b[323])^(a[389] & b[324])^(a[388] & b[325])^(a[387] & b[326])^(a[386] & b[327])^(a[385] & b[328])^(a[384] & b[329])^(a[383] & b[330])^(a[382] & b[331])^(a[381] & b[332])^(a[380] & b[333])^(a[379] & b[334])^(a[378] & b[335])^(a[377] & b[336])^(a[376] & b[337])^(a[375] & b[338])^(a[374] & b[339])^(a[373] & b[340])^(a[372] & b[341])^(a[371] & b[342])^(a[370] & b[343])^(a[369] & b[344])^(a[368] & b[345])^(a[367] & b[346])^(a[366] & b[347])^(a[365] & b[348])^(a[364] & b[349])^(a[363] & b[350])^(a[362] & b[351])^(a[361] & b[352])^(a[360] & b[353])^(a[359] & b[354])^(a[358] & b[355])^(a[357] & b[356])^(a[356] & b[357])^(a[355] & b[358])^(a[354] & b[359])^(a[353] & b[360])^(a[352] & b[361])^(a[351] & b[362])^(a[350] & b[363])^(a[349] & b[364])^(a[348] & b[365])^(a[347] & b[366])^(a[346] & b[367])^(a[345] & b[368])^(a[344] & b[369])^(a[343] & b[370])^(a[342] & b[371])^(a[341] & b[372])^(a[340] & b[373])^(a[339] & b[374])^(a[338] & b[375])^(a[337] & b[376])^(a[336] & b[377])^(a[335] & b[378])^(a[334] & b[379])^(a[333] & b[380])^(a[332] & b[381])^(a[331] & b[382])^(a[330] & b[383])^(a[329] & b[384])^(a[328] & b[385])^(a[327] & b[386])^(a[326] & b[387])^(a[325] & b[388])^(a[324] & b[389])^(a[323] & b[390])^(a[322] & b[391])^(a[321] & b[392])^(a[320] & b[393])^(a[319] & b[394])^(a[318] & b[395])^(a[317] & b[396])^(a[316] & b[397])^(a[315] & b[398])^(a[314] & b[399])^(a[313] & b[400])^(a[312] & b[401])^(a[311] & b[402])^(a[310] & b[403])^(a[309] & b[404])^(a[308] & b[405])^(a[307] & b[406])^(a[306] & b[407])^(a[305] & b[408]);
assign y[714] = (a[408] & b[306])^(a[407] & b[307])^(a[406] & b[308])^(a[405] & b[309])^(a[404] & b[310])^(a[403] & b[311])^(a[402] & b[312])^(a[401] & b[313])^(a[400] & b[314])^(a[399] & b[315])^(a[398] & b[316])^(a[397] & b[317])^(a[396] & b[318])^(a[395] & b[319])^(a[394] & b[320])^(a[393] & b[321])^(a[392] & b[322])^(a[391] & b[323])^(a[390] & b[324])^(a[389] & b[325])^(a[388] & b[326])^(a[387] & b[327])^(a[386] & b[328])^(a[385] & b[329])^(a[384] & b[330])^(a[383] & b[331])^(a[382] & b[332])^(a[381] & b[333])^(a[380] & b[334])^(a[379] & b[335])^(a[378] & b[336])^(a[377] & b[337])^(a[376] & b[338])^(a[375] & b[339])^(a[374] & b[340])^(a[373] & b[341])^(a[372] & b[342])^(a[371] & b[343])^(a[370] & b[344])^(a[369] & b[345])^(a[368] & b[346])^(a[367] & b[347])^(a[366] & b[348])^(a[365] & b[349])^(a[364] & b[350])^(a[363] & b[351])^(a[362] & b[352])^(a[361] & b[353])^(a[360] & b[354])^(a[359] & b[355])^(a[358] & b[356])^(a[357] & b[357])^(a[356] & b[358])^(a[355] & b[359])^(a[354] & b[360])^(a[353] & b[361])^(a[352] & b[362])^(a[351] & b[363])^(a[350] & b[364])^(a[349] & b[365])^(a[348] & b[366])^(a[347] & b[367])^(a[346] & b[368])^(a[345] & b[369])^(a[344] & b[370])^(a[343] & b[371])^(a[342] & b[372])^(a[341] & b[373])^(a[340] & b[374])^(a[339] & b[375])^(a[338] & b[376])^(a[337] & b[377])^(a[336] & b[378])^(a[335] & b[379])^(a[334] & b[380])^(a[333] & b[381])^(a[332] & b[382])^(a[331] & b[383])^(a[330] & b[384])^(a[329] & b[385])^(a[328] & b[386])^(a[327] & b[387])^(a[326] & b[388])^(a[325] & b[389])^(a[324] & b[390])^(a[323] & b[391])^(a[322] & b[392])^(a[321] & b[393])^(a[320] & b[394])^(a[319] & b[395])^(a[318] & b[396])^(a[317] & b[397])^(a[316] & b[398])^(a[315] & b[399])^(a[314] & b[400])^(a[313] & b[401])^(a[312] & b[402])^(a[311] & b[403])^(a[310] & b[404])^(a[309] & b[405])^(a[308] & b[406])^(a[307] & b[407])^(a[306] & b[408]);
assign y[715] = (a[408] & b[307])^(a[407] & b[308])^(a[406] & b[309])^(a[405] & b[310])^(a[404] & b[311])^(a[403] & b[312])^(a[402] & b[313])^(a[401] & b[314])^(a[400] & b[315])^(a[399] & b[316])^(a[398] & b[317])^(a[397] & b[318])^(a[396] & b[319])^(a[395] & b[320])^(a[394] & b[321])^(a[393] & b[322])^(a[392] & b[323])^(a[391] & b[324])^(a[390] & b[325])^(a[389] & b[326])^(a[388] & b[327])^(a[387] & b[328])^(a[386] & b[329])^(a[385] & b[330])^(a[384] & b[331])^(a[383] & b[332])^(a[382] & b[333])^(a[381] & b[334])^(a[380] & b[335])^(a[379] & b[336])^(a[378] & b[337])^(a[377] & b[338])^(a[376] & b[339])^(a[375] & b[340])^(a[374] & b[341])^(a[373] & b[342])^(a[372] & b[343])^(a[371] & b[344])^(a[370] & b[345])^(a[369] & b[346])^(a[368] & b[347])^(a[367] & b[348])^(a[366] & b[349])^(a[365] & b[350])^(a[364] & b[351])^(a[363] & b[352])^(a[362] & b[353])^(a[361] & b[354])^(a[360] & b[355])^(a[359] & b[356])^(a[358] & b[357])^(a[357] & b[358])^(a[356] & b[359])^(a[355] & b[360])^(a[354] & b[361])^(a[353] & b[362])^(a[352] & b[363])^(a[351] & b[364])^(a[350] & b[365])^(a[349] & b[366])^(a[348] & b[367])^(a[347] & b[368])^(a[346] & b[369])^(a[345] & b[370])^(a[344] & b[371])^(a[343] & b[372])^(a[342] & b[373])^(a[341] & b[374])^(a[340] & b[375])^(a[339] & b[376])^(a[338] & b[377])^(a[337] & b[378])^(a[336] & b[379])^(a[335] & b[380])^(a[334] & b[381])^(a[333] & b[382])^(a[332] & b[383])^(a[331] & b[384])^(a[330] & b[385])^(a[329] & b[386])^(a[328] & b[387])^(a[327] & b[388])^(a[326] & b[389])^(a[325] & b[390])^(a[324] & b[391])^(a[323] & b[392])^(a[322] & b[393])^(a[321] & b[394])^(a[320] & b[395])^(a[319] & b[396])^(a[318] & b[397])^(a[317] & b[398])^(a[316] & b[399])^(a[315] & b[400])^(a[314] & b[401])^(a[313] & b[402])^(a[312] & b[403])^(a[311] & b[404])^(a[310] & b[405])^(a[309] & b[406])^(a[308] & b[407])^(a[307] & b[408]);
assign y[716] = (a[408] & b[308])^(a[407] & b[309])^(a[406] & b[310])^(a[405] & b[311])^(a[404] & b[312])^(a[403] & b[313])^(a[402] & b[314])^(a[401] & b[315])^(a[400] & b[316])^(a[399] & b[317])^(a[398] & b[318])^(a[397] & b[319])^(a[396] & b[320])^(a[395] & b[321])^(a[394] & b[322])^(a[393] & b[323])^(a[392] & b[324])^(a[391] & b[325])^(a[390] & b[326])^(a[389] & b[327])^(a[388] & b[328])^(a[387] & b[329])^(a[386] & b[330])^(a[385] & b[331])^(a[384] & b[332])^(a[383] & b[333])^(a[382] & b[334])^(a[381] & b[335])^(a[380] & b[336])^(a[379] & b[337])^(a[378] & b[338])^(a[377] & b[339])^(a[376] & b[340])^(a[375] & b[341])^(a[374] & b[342])^(a[373] & b[343])^(a[372] & b[344])^(a[371] & b[345])^(a[370] & b[346])^(a[369] & b[347])^(a[368] & b[348])^(a[367] & b[349])^(a[366] & b[350])^(a[365] & b[351])^(a[364] & b[352])^(a[363] & b[353])^(a[362] & b[354])^(a[361] & b[355])^(a[360] & b[356])^(a[359] & b[357])^(a[358] & b[358])^(a[357] & b[359])^(a[356] & b[360])^(a[355] & b[361])^(a[354] & b[362])^(a[353] & b[363])^(a[352] & b[364])^(a[351] & b[365])^(a[350] & b[366])^(a[349] & b[367])^(a[348] & b[368])^(a[347] & b[369])^(a[346] & b[370])^(a[345] & b[371])^(a[344] & b[372])^(a[343] & b[373])^(a[342] & b[374])^(a[341] & b[375])^(a[340] & b[376])^(a[339] & b[377])^(a[338] & b[378])^(a[337] & b[379])^(a[336] & b[380])^(a[335] & b[381])^(a[334] & b[382])^(a[333] & b[383])^(a[332] & b[384])^(a[331] & b[385])^(a[330] & b[386])^(a[329] & b[387])^(a[328] & b[388])^(a[327] & b[389])^(a[326] & b[390])^(a[325] & b[391])^(a[324] & b[392])^(a[323] & b[393])^(a[322] & b[394])^(a[321] & b[395])^(a[320] & b[396])^(a[319] & b[397])^(a[318] & b[398])^(a[317] & b[399])^(a[316] & b[400])^(a[315] & b[401])^(a[314] & b[402])^(a[313] & b[403])^(a[312] & b[404])^(a[311] & b[405])^(a[310] & b[406])^(a[309] & b[407])^(a[308] & b[408]);
assign y[717] = (a[408] & b[309])^(a[407] & b[310])^(a[406] & b[311])^(a[405] & b[312])^(a[404] & b[313])^(a[403] & b[314])^(a[402] & b[315])^(a[401] & b[316])^(a[400] & b[317])^(a[399] & b[318])^(a[398] & b[319])^(a[397] & b[320])^(a[396] & b[321])^(a[395] & b[322])^(a[394] & b[323])^(a[393] & b[324])^(a[392] & b[325])^(a[391] & b[326])^(a[390] & b[327])^(a[389] & b[328])^(a[388] & b[329])^(a[387] & b[330])^(a[386] & b[331])^(a[385] & b[332])^(a[384] & b[333])^(a[383] & b[334])^(a[382] & b[335])^(a[381] & b[336])^(a[380] & b[337])^(a[379] & b[338])^(a[378] & b[339])^(a[377] & b[340])^(a[376] & b[341])^(a[375] & b[342])^(a[374] & b[343])^(a[373] & b[344])^(a[372] & b[345])^(a[371] & b[346])^(a[370] & b[347])^(a[369] & b[348])^(a[368] & b[349])^(a[367] & b[350])^(a[366] & b[351])^(a[365] & b[352])^(a[364] & b[353])^(a[363] & b[354])^(a[362] & b[355])^(a[361] & b[356])^(a[360] & b[357])^(a[359] & b[358])^(a[358] & b[359])^(a[357] & b[360])^(a[356] & b[361])^(a[355] & b[362])^(a[354] & b[363])^(a[353] & b[364])^(a[352] & b[365])^(a[351] & b[366])^(a[350] & b[367])^(a[349] & b[368])^(a[348] & b[369])^(a[347] & b[370])^(a[346] & b[371])^(a[345] & b[372])^(a[344] & b[373])^(a[343] & b[374])^(a[342] & b[375])^(a[341] & b[376])^(a[340] & b[377])^(a[339] & b[378])^(a[338] & b[379])^(a[337] & b[380])^(a[336] & b[381])^(a[335] & b[382])^(a[334] & b[383])^(a[333] & b[384])^(a[332] & b[385])^(a[331] & b[386])^(a[330] & b[387])^(a[329] & b[388])^(a[328] & b[389])^(a[327] & b[390])^(a[326] & b[391])^(a[325] & b[392])^(a[324] & b[393])^(a[323] & b[394])^(a[322] & b[395])^(a[321] & b[396])^(a[320] & b[397])^(a[319] & b[398])^(a[318] & b[399])^(a[317] & b[400])^(a[316] & b[401])^(a[315] & b[402])^(a[314] & b[403])^(a[313] & b[404])^(a[312] & b[405])^(a[311] & b[406])^(a[310] & b[407])^(a[309] & b[408]);
assign y[718] = (a[408] & b[310])^(a[407] & b[311])^(a[406] & b[312])^(a[405] & b[313])^(a[404] & b[314])^(a[403] & b[315])^(a[402] & b[316])^(a[401] & b[317])^(a[400] & b[318])^(a[399] & b[319])^(a[398] & b[320])^(a[397] & b[321])^(a[396] & b[322])^(a[395] & b[323])^(a[394] & b[324])^(a[393] & b[325])^(a[392] & b[326])^(a[391] & b[327])^(a[390] & b[328])^(a[389] & b[329])^(a[388] & b[330])^(a[387] & b[331])^(a[386] & b[332])^(a[385] & b[333])^(a[384] & b[334])^(a[383] & b[335])^(a[382] & b[336])^(a[381] & b[337])^(a[380] & b[338])^(a[379] & b[339])^(a[378] & b[340])^(a[377] & b[341])^(a[376] & b[342])^(a[375] & b[343])^(a[374] & b[344])^(a[373] & b[345])^(a[372] & b[346])^(a[371] & b[347])^(a[370] & b[348])^(a[369] & b[349])^(a[368] & b[350])^(a[367] & b[351])^(a[366] & b[352])^(a[365] & b[353])^(a[364] & b[354])^(a[363] & b[355])^(a[362] & b[356])^(a[361] & b[357])^(a[360] & b[358])^(a[359] & b[359])^(a[358] & b[360])^(a[357] & b[361])^(a[356] & b[362])^(a[355] & b[363])^(a[354] & b[364])^(a[353] & b[365])^(a[352] & b[366])^(a[351] & b[367])^(a[350] & b[368])^(a[349] & b[369])^(a[348] & b[370])^(a[347] & b[371])^(a[346] & b[372])^(a[345] & b[373])^(a[344] & b[374])^(a[343] & b[375])^(a[342] & b[376])^(a[341] & b[377])^(a[340] & b[378])^(a[339] & b[379])^(a[338] & b[380])^(a[337] & b[381])^(a[336] & b[382])^(a[335] & b[383])^(a[334] & b[384])^(a[333] & b[385])^(a[332] & b[386])^(a[331] & b[387])^(a[330] & b[388])^(a[329] & b[389])^(a[328] & b[390])^(a[327] & b[391])^(a[326] & b[392])^(a[325] & b[393])^(a[324] & b[394])^(a[323] & b[395])^(a[322] & b[396])^(a[321] & b[397])^(a[320] & b[398])^(a[319] & b[399])^(a[318] & b[400])^(a[317] & b[401])^(a[316] & b[402])^(a[315] & b[403])^(a[314] & b[404])^(a[313] & b[405])^(a[312] & b[406])^(a[311] & b[407])^(a[310] & b[408]);
assign y[719] = (a[408] & b[311])^(a[407] & b[312])^(a[406] & b[313])^(a[405] & b[314])^(a[404] & b[315])^(a[403] & b[316])^(a[402] & b[317])^(a[401] & b[318])^(a[400] & b[319])^(a[399] & b[320])^(a[398] & b[321])^(a[397] & b[322])^(a[396] & b[323])^(a[395] & b[324])^(a[394] & b[325])^(a[393] & b[326])^(a[392] & b[327])^(a[391] & b[328])^(a[390] & b[329])^(a[389] & b[330])^(a[388] & b[331])^(a[387] & b[332])^(a[386] & b[333])^(a[385] & b[334])^(a[384] & b[335])^(a[383] & b[336])^(a[382] & b[337])^(a[381] & b[338])^(a[380] & b[339])^(a[379] & b[340])^(a[378] & b[341])^(a[377] & b[342])^(a[376] & b[343])^(a[375] & b[344])^(a[374] & b[345])^(a[373] & b[346])^(a[372] & b[347])^(a[371] & b[348])^(a[370] & b[349])^(a[369] & b[350])^(a[368] & b[351])^(a[367] & b[352])^(a[366] & b[353])^(a[365] & b[354])^(a[364] & b[355])^(a[363] & b[356])^(a[362] & b[357])^(a[361] & b[358])^(a[360] & b[359])^(a[359] & b[360])^(a[358] & b[361])^(a[357] & b[362])^(a[356] & b[363])^(a[355] & b[364])^(a[354] & b[365])^(a[353] & b[366])^(a[352] & b[367])^(a[351] & b[368])^(a[350] & b[369])^(a[349] & b[370])^(a[348] & b[371])^(a[347] & b[372])^(a[346] & b[373])^(a[345] & b[374])^(a[344] & b[375])^(a[343] & b[376])^(a[342] & b[377])^(a[341] & b[378])^(a[340] & b[379])^(a[339] & b[380])^(a[338] & b[381])^(a[337] & b[382])^(a[336] & b[383])^(a[335] & b[384])^(a[334] & b[385])^(a[333] & b[386])^(a[332] & b[387])^(a[331] & b[388])^(a[330] & b[389])^(a[329] & b[390])^(a[328] & b[391])^(a[327] & b[392])^(a[326] & b[393])^(a[325] & b[394])^(a[324] & b[395])^(a[323] & b[396])^(a[322] & b[397])^(a[321] & b[398])^(a[320] & b[399])^(a[319] & b[400])^(a[318] & b[401])^(a[317] & b[402])^(a[316] & b[403])^(a[315] & b[404])^(a[314] & b[405])^(a[313] & b[406])^(a[312] & b[407])^(a[311] & b[408]);
assign y[720] = (a[408] & b[312])^(a[407] & b[313])^(a[406] & b[314])^(a[405] & b[315])^(a[404] & b[316])^(a[403] & b[317])^(a[402] & b[318])^(a[401] & b[319])^(a[400] & b[320])^(a[399] & b[321])^(a[398] & b[322])^(a[397] & b[323])^(a[396] & b[324])^(a[395] & b[325])^(a[394] & b[326])^(a[393] & b[327])^(a[392] & b[328])^(a[391] & b[329])^(a[390] & b[330])^(a[389] & b[331])^(a[388] & b[332])^(a[387] & b[333])^(a[386] & b[334])^(a[385] & b[335])^(a[384] & b[336])^(a[383] & b[337])^(a[382] & b[338])^(a[381] & b[339])^(a[380] & b[340])^(a[379] & b[341])^(a[378] & b[342])^(a[377] & b[343])^(a[376] & b[344])^(a[375] & b[345])^(a[374] & b[346])^(a[373] & b[347])^(a[372] & b[348])^(a[371] & b[349])^(a[370] & b[350])^(a[369] & b[351])^(a[368] & b[352])^(a[367] & b[353])^(a[366] & b[354])^(a[365] & b[355])^(a[364] & b[356])^(a[363] & b[357])^(a[362] & b[358])^(a[361] & b[359])^(a[360] & b[360])^(a[359] & b[361])^(a[358] & b[362])^(a[357] & b[363])^(a[356] & b[364])^(a[355] & b[365])^(a[354] & b[366])^(a[353] & b[367])^(a[352] & b[368])^(a[351] & b[369])^(a[350] & b[370])^(a[349] & b[371])^(a[348] & b[372])^(a[347] & b[373])^(a[346] & b[374])^(a[345] & b[375])^(a[344] & b[376])^(a[343] & b[377])^(a[342] & b[378])^(a[341] & b[379])^(a[340] & b[380])^(a[339] & b[381])^(a[338] & b[382])^(a[337] & b[383])^(a[336] & b[384])^(a[335] & b[385])^(a[334] & b[386])^(a[333] & b[387])^(a[332] & b[388])^(a[331] & b[389])^(a[330] & b[390])^(a[329] & b[391])^(a[328] & b[392])^(a[327] & b[393])^(a[326] & b[394])^(a[325] & b[395])^(a[324] & b[396])^(a[323] & b[397])^(a[322] & b[398])^(a[321] & b[399])^(a[320] & b[400])^(a[319] & b[401])^(a[318] & b[402])^(a[317] & b[403])^(a[316] & b[404])^(a[315] & b[405])^(a[314] & b[406])^(a[313] & b[407])^(a[312] & b[408]);
assign y[721] = (a[408] & b[313])^(a[407] & b[314])^(a[406] & b[315])^(a[405] & b[316])^(a[404] & b[317])^(a[403] & b[318])^(a[402] & b[319])^(a[401] & b[320])^(a[400] & b[321])^(a[399] & b[322])^(a[398] & b[323])^(a[397] & b[324])^(a[396] & b[325])^(a[395] & b[326])^(a[394] & b[327])^(a[393] & b[328])^(a[392] & b[329])^(a[391] & b[330])^(a[390] & b[331])^(a[389] & b[332])^(a[388] & b[333])^(a[387] & b[334])^(a[386] & b[335])^(a[385] & b[336])^(a[384] & b[337])^(a[383] & b[338])^(a[382] & b[339])^(a[381] & b[340])^(a[380] & b[341])^(a[379] & b[342])^(a[378] & b[343])^(a[377] & b[344])^(a[376] & b[345])^(a[375] & b[346])^(a[374] & b[347])^(a[373] & b[348])^(a[372] & b[349])^(a[371] & b[350])^(a[370] & b[351])^(a[369] & b[352])^(a[368] & b[353])^(a[367] & b[354])^(a[366] & b[355])^(a[365] & b[356])^(a[364] & b[357])^(a[363] & b[358])^(a[362] & b[359])^(a[361] & b[360])^(a[360] & b[361])^(a[359] & b[362])^(a[358] & b[363])^(a[357] & b[364])^(a[356] & b[365])^(a[355] & b[366])^(a[354] & b[367])^(a[353] & b[368])^(a[352] & b[369])^(a[351] & b[370])^(a[350] & b[371])^(a[349] & b[372])^(a[348] & b[373])^(a[347] & b[374])^(a[346] & b[375])^(a[345] & b[376])^(a[344] & b[377])^(a[343] & b[378])^(a[342] & b[379])^(a[341] & b[380])^(a[340] & b[381])^(a[339] & b[382])^(a[338] & b[383])^(a[337] & b[384])^(a[336] & b[385])^(a[335] & b[386])^(a[334] & b[387])^(a[333] & b[388])^(a[332] & b[389])^(a[331] & b[390])^(a[330] & b[391])^(a[329] & b[392])^(a[328] & b[393])^(a[327] & b[394])^(a[326] & b[395])^(a[325] & b[396])^(a[324] & b[397])^(a[323] & b[398])^(a[322] & b[399])^(a[321] & b[400])^(a[320] & b[401])^(a[319] & b[402])^(a[318] & b[403])^(a[317] & b[404])^(a[316] & b[405])^(a[315] & b[406])^(a[314] & b[407])^(a[313] & b[408]);
assign y[722] = (a[408] & b[314])^(a[407] & b[315])^(a[406] & b[316])^(a[405] & b[317])^(a[404] & b[318])^(a[403] & b[319])^(a[402] & b[320])^(a[401] & b[321])^(a[400] & b[322])^(a[399] & b[323])^(a[398] & b[324])^(a[397] & b[325])^(a[396] & b[326])^(a[395] & b[327])^(a[394] & b[328])^(a[393] & b[329])^(a[392] & b[330])^(a[391] & b[331])^(a[390] & b[332])^(a[389] & b[333])^(a[388] & b[334])^(a[387] & b[335])^(a[386] & b[336])^(a[385] & b[337])^(a[384] & b[338])^(a[383] & b[339])^(a[382] & b[340])^(a[381] & b[341])^(a[380] & b[342])^(a[379] & b[343])^(a[378] & b[344])^(a[377] & b[345])^(a[376] & b[346])^(a[375] & b[347])^(a[374] & b[348])^(a[373] & b[349])^(a[372] & b[350])^(a[371] & b[351])^(a[370] & b[352])^(a[369] & b[353])^(a[368] & b[354])^(a[367] & b[355])^(a[366] & b[356])^(a[365] & b[357])^(a[364] & b[358])^(a[363] & b[359])^(a[362] & b[360])^(a[361] & b[361])^(a[360] & b[362])^(a[359] & b[363])^(a[358] & b[364])^(a[357] & b[365])^(a[356] & b[366])^(a[355] & b[367])^(a[354] & b[368])^(a[353] & b[369])^(a[352] & b[370])^(a[351] & b[371])^(a[350] & b[372])^(a[349] & b[373])^(a[348] & b[374])^(a[347] & b[375])^(a[346] & b[376])^(a[345] & b[377])^(a[344] & b[378])^(a[343] & b[379])^(a[342] & b[380])^(a[341] & b[381])^(a[340] & b[382])^(a[339] & b[383])^(a[338] & b[384])^(a[337] & b[385])^(a[336] & b[386])^(a[335] & b[387])^(a[334] & b[388])^(a[333] & b[389])^(a[332] & b[390])^(a[331] & b[391])^(a[330] & b[392])^(a[329] & b[393])^(a[328] & b[394])^(a[327] & b[395])^(a[326] & b[396])^(a[325] & b[397])^(a[324] & b[398])^(a[323] & b[399])^(a[322] & b[400])^(a[321] & b[401])^(a[320] & b[402])^(a[319] & b[403])^(a[318] & b[404])^(a[317] & b[405])^(a[316] & b[406])^(a[315] & b[407])^(a[314] & b[408]);
assign y[723] = (a[408] & b[315])^(a[407] & b[316])^(a[406] & b[317])^(a[405] & b[318])^(a[404] & b[319])^(a[403] & b[320])^(a[402] & b[321])^(a[401] & b[322])^(a[400] & b[323])^(a[399] & b[324])^(a[398] & b[325])^(a[397] & b[326])^(a[396] & b[327])^(a[395] & b[328])^(a[394] & b[329])^(a[393] & b[330])^(a[392] & b[331])^(a[391] & b[332])^(a[390] & b[333])^(a[389] & b[334])^(a[388] & b[335])^(a[387] & b[336])^(a[386] & b[337])^(a[385] & b[338])^(a[384] & b[339])^(a[383] & b[340])^(a[382] & b[341])^(a[381] & b[342])^(a[380] & b[343])^(a[379] & b[344])^(a[378] & b[345])^(a[377] & b[346])^(a[376] & b[347])^(a[375] & b[348])^(a[374] & b[349])^(a[373] & b[350])^(a[372] & b[351])^(a[371] & b[352])^(a[370] & b[353])^(a[369] & b[354])^(a[368] & b[355])^(a[367] & b[356])^(a[366] & b[357])^(a[365] & b[358])^(a[364] & b[359])^(a[363] & b[360])^(a[362] & b[361])^(a[361] & b[362])^(a[360] & b[363])^(a[359] & b[364])^(a[358] & b[365])^(a[357] & b[366])^(a[356] & b[367])^(a[355] & b[368])^(a[354] & b[369])^(a[353] & b[370])^(a[352] & b[371])^(a[351] & b[372])^(a[350] & b[373])^(a[349] & b[374])^(a[348] & b[375])^(a[347] & b[376])^(a[346] & b[377])^(a[345] & b[378])^(a[344] & b[379])^(a[343] & b[380])^(a[342] & b[381])^(a[341] & b[382])^(a[340] & b[383])^(a[339] & b[384])^(a[338] & b[385])^(a[337] & b[386])^(a[336] & b[387])^(a[335] & b[388])^(a[334] & b[389])^(a[333] & b[390])^(a[332] & b[391])^(a[331] & b[392])^(a[330] & b[393])^(a[329] & b[394])^(a[328] & b[395])^(a[327] & b[396])^(a[326] & b[397])^(a[325] & b[398])^(a[324] & b[399])^(a[323] & b[400])^(a[322] & b[401])^(a[321] & b[402])^(a[320] & b[403])^(a[319] & b[404])^(a[318] & b[405])^(a[317] & b[406])^(a[316] & b[407])^(a[315] & b[408]);
assign y[724] = (a[408] & b[316])^(a[407] & b[317])^(a[406] & b[318])^(a[405] & b[319])^(a[404] & b[320])^(a[403] & b[321])^(a[402] & b[322])^(a[401] & b[323])^(a[400] & b[324])^(a[399] & b[325])^(a[398] & b[326])^(a[397] & b[327])^(a[396] & b[328])^(a[395] & b[329])^(a[394] & b[330])^(a[393] & b[331])^(a[392] & b[332])^(a[391] & b[333])^(a[390] & b[334])^(a[389] & b[335])^(a[388] & b[336])^(a[387] & b[337])^(a[386] & b[338])^(a[385] & b[339])^(a[384] & b[340])^(a[383] & b[341])^(a[382] & b[342])^(a[381] & b[343])^(a[380] & b[344])^(a[379] & b[345])^(a[378] & b[346])^(a[377] & b[347])^(a[376] & b[348])^(a[375] & b[349])^(a[374] & b[350])^(a[373] & b[351])^(a[372] & b[352])^(a[371] & b[353])^(a[370] & b[354])^(a[369] & b[355])^(a[368] & b[356])^(a[367] & b[357])^(a[366] & b[358])^(a[365] & b[359])^(a[364] & b[360])^(a[363] & b[361])^(a[362] & b[362])^(a[361] & b[363])^(a[360] & b[364])^(a[359] & b[365])^(a[358] & b[366])^(a[357] & b[367])^(a[356] & b[368])^(a[355] & b[369])^(a[354] & b[370])^(a[353] & b[371])^(a[352] & b[372])^(a[351] & b[373])^(a[350] & b[374])^(a[349] & b[375])^(a[348] & b[376])^(a[347] & b[377])^(a[346] & b[378])^(a[345] & b[379])^(a[344] & b[380])^(a[343] & b[381])^(a[342] & b[382])^(a[341] & b[383])^(a[340] & b[384])^(a[339] & b[385])^(a[338] & b[386])^(a[337] & b[387])^(a[336] & b[388])^(a[335] & b[389])^(a[334] & b[390])^(a[333] & b[391])^(a[332] & b[392])^(a[331] & b[393])^(a[330] & b[394])^(a[329] & b[395])^(a[328] & b[396])^(a[327] & b[397])^(a[326] & b[398])^(a[325] & b[399])^(a[324] & b[400])^(a[323] & b[401])^(a[322] & b[402])^(a[321] & b[403])^(a[320] & b[404])^(a[319] & b[405])^(a[318] & b[406])^(a[317] & b[407])^(a[316] & b[408]);
assign y[725] = (a[408] & b[317])^(a[407] & b[318])^(a[406] & b[319])^(a[405] & b[320])^(a[404] & b[321])^(a[403] & b[322])^(a[402] & b[323])^(a[401] & b[324])^(a[400] & b[325])^(a[399] & b[326])^(a[398] & b[327])^(a[397] & b[328])^(a[396] & b[329])^(a[395] & b[330])^(a[394] & b[331])^(a[393] & b[332])^(a[392] & b[333])^(a[391] & b[334])^(a[390] & b[335])^(a[389] & b[336])^(a[388] & b[337])^(a[387] & b[338])^(a[386] & b[339])^(a[385] & b[340])^(a[384] & b[341])^(a[383] & b[342])^(a[382] & b[343])^(a[381] & b[344])^(a[380] & b[345])^(a[379] & b[346])^(a[378] & b[347])^(a[377] & b[348])^(a[376] & b[349])^(a[375] & b[350])^(a[374] & b[351])^(a[373] & b[352])^(a[372] & b[353])^(a[371] & b[354])^(a[370] & b[355])^(a[369] & b[356])^(a[368] & b[357])^(a[367] & b[358])^(a[366] & b[359])^(a[365] & b[360])^(a[364] & b[361])^(a[363] & b[362])^(a[362] & b[363])^(a[361] & b[364])^(a[360] & b[365])^(a[359] & b[366])^(a[358] & b[367])^(a[357] & b[368])^(a[356] & b[369])^(a[355] & b[370])^(a[354] & b[371])^(a[353] & b[372])^(a[352] & b[373])^(a[351] & b[374])^(a[350] & b[375])^(a[349] & b[376])^(a[348] & b[377])^(a[347] & b[378])^(a[346] & b[379])^(a[345] & b[380])^(a[344] & b[381])^(a[343] & b[382])^(a[342] & b[383])^(a[341] & b[384])^(a[340] & b[385])^(a[339] & b[386])^(a[338] & b[387])^(a[337] & b[388])^(a[336] & b[389])^(a[335] & b[390])^(a[334] & b[391])^(a[333] & b[392])^(a[332] & b[393])^(a[331] & b[394])^(a[330] & b[395])^(a[329] & b[396])^(a[328] & b[397])^(a[327] & b[398])^(a[326] & b[399])^(a[325] & b[400])^(a[324] & b[401])^(a[323] & b[402])^(a[322] & b[403])^(a[321] & b[404])^(a[320] & b[405])^(a[319] & b[406])^(a[318] & b[407])^(a[317] & b[408]);
assign y[726] = (a[408] & b[318])^(a[407] & b[319])^(a[406] & b[320])^(a[405] & b[321])^(a[404] & b[322])^(a[403] & b[323])^(a[402] & b[324])^(a[401] & b[325])^(a[400] & b[326])^(a[399] & b[327])^(a[398] & b[328])^(a[397] & b[329])^(a[396] & b[330])^(a[395] & b[331])^(a[394] & b[332])^(a[393] & b[333])^(a[392] & b[334])^(a[391] & b[335])^(a[390] & b[336])^(a[389] & b[337])^(a[388] & b[338])^(a[387] & b[339])^(a[386] & b[340])^(a[385] & b[341])^(a[384] & b[342])^(a[383] & b[343])^(a[382] & b[344])^(a[381] & b[345])^(a[380] & b[346])^(a[379] & b[347])^(a[378] & b[348])^(a[377] & b[349])^(a[376] & b[350])^(a[375] & b[351])^(a[374] & b[352])^(a[373] & b[353])^(a[372] & b[354])^(a[371] & b[355])^(a[370] & b[356])^(a[369] & b[357])^(a[368] & b[358])^(a[367] & b[359])^(a[366] & b[360])^(a[365] & b[361])^(a[364] & b[362])^(a[363] & b[363])^(a[362] & b[364])^(a[361] & b[365])^(a[360] & b[366])^(a[359] & b[367])^(a[358] & b[368])^(a[357] & b[369])^(a[356] & b[370])^(a[355] & b[371])^(a[354] & b[372])^(a[353] & b[373])^(a[352] & b[374])^(a[351] & b[375])^(a[350] & b[376])^(a[349] & b[377])^(a[348] & b[378])^(a[347] & b[379])^(a[346] & b[380])^(a[345] & b[381])^(a[344] & b[382])^(a[343] & b[383])^(a[342] & b[384])^(a[341] & b[385])^(a[340] & b[386])^(a[339] & b[387])^(a[338] & b[388])^(a[337] & b[389])^(a[336] & b[390])^(a[335] & b[391])^(a[334] & b[392])^(a[333] & b[393])^(a[332] & b[394])^(a[331] & b[395])^(a[330] & b[396])^(a[329] & b[397])^(a[328] & b[398])^(a[327] & b[399])^(a[326] & b[400])^(a[325] & b[401])^(a[324] & b[402])^(a[323] & b[403])^(a[322] & b[404])^(a[321] & b[405])^(a[320] & b[406])^(a[319] & b[407])^(a[318] & b[408]);
assign y[727] = (a[408] & b[319])^(a[407] & b[320])^(a[406] & b[321])^(a[405] & b[322])^(a[404] & b[323])^(a[403] & b[324])^(a[402] & b[325])^(a[401] & b[326])^(a[400] & b[327])^(a[399] & b[328])^(a[398] & b[329])^(a[397] & b[330])^(a[396] & b[331])^(a[395] & b[332])^(a[394] & b[333])^(a[393] & b[334])^(a[392] & b[335])^(a[391] & b[336])^(a[390] & b[337])^(a[389] & b[338])^(a[388] & b[339])^(a[387] & b[340])^(a[386] & b[341])^(a[385] & b[342])^(a[384] & b[343])^(a[383] & b[344])^(a[382] & b[345])^(a[381] & b[346])^(a[380] & b[347])^(a[379] & b[348])^(a[378] & b[349])^(a[377] & b[350])^(a[376] & b[351])^(a[375] & b[352])^(a[374] & b[353])^(a[373] & b[354])^(a[372] & b[355])^(a[371] & b[356])^(a[370] & b[357])^(a[369] & b[358])^(a[368] & b[359])^(a[367] & b[360])^(a[366] & b[361])^(a[365] & b[362])^(a[364] & b[363])^(a[363] & b[364])^(a[362] & b[365])^(a[361] & b[366])^(a[360] & b[367])^(a[359] & b[368])^(a[358] & b[369])^(a[357] & b[370])^(a[356] & b[371])^(a[355] & b[372])^(a[354] & b[373])^(a[353] & b[374])^(a[352] & b[375])^(a[351] & b[376])^(a[350] & b[377])^(a[349] & b[378])^(a[348] & b[379])^(a[347] & b[380])^(a[346] & b[381])^(a[345] & b[382])^(a[344] & b[383])^(a[343] & b[384])^(a[342] & b[385])^(a[341] & b[386])^(a[340] & b[387])^(a[339] & b[388])^(a[338] & b[389])^(a[337] & b[390])^(a[336] & b[391])^(a[335] & b[392])^(a[334] & b[393])^(a[333] & b[394])^(a[332] & b[395])^(a[331] & b[396])^(a[330] & b[397])^(a[329] & b[398])^(a[328] & b[399])^(a[327] & b[400])^(a[326] & b[401])^(a[325] & b[402])^(a[324] & b[403])^(a[323] & b[404])^(a[322] & b[405])^(a[321] & b[406])^(a[320] & b[407])^(a[319] & b[408]);
assign y[728] = (a[408] & b[320])^(a[407] & b[321])^(a[406] & b[322])^(a[405] & b[323])^(a[404] & b[324])^(a[403] & b[325])^(a[402] & b[326])^(a[401] & b[327])^(a[400] & b[328])^(a[399] & b[329])^(a[398] & b[330])^(a[397] & b[331])^(a[396] & b[332])^(a[395] & b[333])^(a[394] & b[334])^(a[393] & b[335])^(a[392] & b[336])^(a[391] & b[337])^(a[390] & b[338])^(a[389] & b[339])^(a[388] & b[340])^(a[387] & b[341])^(a[386] & b[342])^(a[385] & b[343])^(a[384] & b[344])^(a[383] & b[345])^(a[382] & b[346])^(a[381] & b[347])^(a[380] & b[348])^(a[379] & b[349])^(a[378] & b[350])^(a[377] & b[351])^(a[376] & b[352])^(a[375] & b[353])^(a[374] & b[354])^(a[373] & b[355])^(a[372] & b[356])^(a[371] & b[357])^(a[370] & b[358])^(a[369] & b[359])^(a[368] & b[360])^(a[367] & b[361])^(a[366] & b[362])^(a[365] & b[363])^(a[364] & b[364])^(a[363] & b[365])^(a[362] & b[366])^(a[361] & b[367])^(a[360] & b[368])^(a[359] & b[369])^(a[358] & b[370])^(a[357] & b[371])^(a[356] & b[372])^(a[355] & b[373])^(a[354] & b[374])^(a[353] & b[375])^(a[352] & b[376])^(a[351] & b[377])^(a[350] & b[378])^(a[349] & b[379])^(a[348] & b[380])^(a[347] & b[381])^(a[346] & b[382])^(a[345] & b[383])^(a[344] & b[384])^(a[343] & b[385])^(a[342] & b[386])^(a[341] & b[387])^(a[340] & b[388])^(a[339] & b[389])^(a[338] & b[390])^(a[337] & b[391])^(a[336] & b[392])^(a[335] & b[393])^(a[334] & b[394])^(a[333] & b[395])^(a[332] & b[396])^(a[331] & b[397])^(a[330] & b[398])^(a[329] & b[399])^(a[328] & b[400])^(a[327] & b[401])^(a[326] & b[402])^(a[325] & b[403])^(a[324] & b[404])^(a[323] & b[405])^(a[322] & b[406])^(a[321] & b[407])^(a[320] & b[408]);
assign y[729] = (a[408] & b[321])^(a[407] & b[322])^(a[406] & b[323])^(a[405] & b[324])^(a[404] & b[325])^(a[403] & b[326])^(a[402] & b[327])^(a[401] & b[328])^(a[400] & b[329])^(a[399] & b[330])^(a[398] & b[331])^(a[397] & b[332])^(a[396] & b[333])^(a[395] & b[334])^(a[394] & b[335])^(a[393] & b[336])^(a[392] & b[337])^(a[391] & b[338])^(a[390] & b[339])^(a[389] & b[340])^(a[388] & b[341])^(a[387] & b[342])^(a[386] & b[343])^(a[385] & b[344])^(a[384] & b[345])^(a[383] & b[346])^(a[382] & b[347])^(a[381] & b[348])^(a[380] & b[349])^(a[379] & b[350])^(a[378] & b[351])^(a[377] & b[352])^(a[376] & b[353])^(a[375] & b[354])^(a[374] & b[355])^(a[373] & b[356])^(a[372] & b[357])^(a[371] & b[358])^(a[370] & b[359])^(a[369] & b[360])^(a[368] & b[361])^(a[367] & b[362])^(a[366] & b[363])^(a[365] & b[364])^(a[364] & b[365])^(a[363] & b[366])^(a[362] & b[367])^(a[361] & b[368])^(a[360] & b[369])^(a[359] & b[370])^(a[358] & b[371])^(a[357] & b[372])^(a[356] & b[373])^(a[355] & b[374])^(a[354] & b[375])^(a[353] & b[376])^(a[352] & b[377])^(a[351] & b[378])^(a[350] & b[379])^(a[349] & b[380])^(a[348] & b[381])^(a[347] & b[382])^(a[346] & b[383])^(a[345] & b[384])^(a[344] & b[385])^(a[343] & b[386])^(a[342] & b[387])^(a[341] & b[388])^(a[340] & b[389])^(a[339] & b[390])^(a[338] & b[391])^(a[337] & b[392])^(a[336] & b[393])^(a[335] & b[394])^(a[334] & b[395])^(a[333] & b[396])^(a[332] & b[397])^(a[331] & b[398])^(a[330] & b[399])^(a[329] & b[400])^(a[328] & b[401])^(a[327] & b[402])^(a[326] & b[403])^(a[325] & b[404])^(a[324] & b[405])^(a[323] & b[406])^(a[322] & b[407])^(a[321] & b[408]);
assign y[730] = (a[408] & b[322])^(a[407] & b[323])^(a[406] & b[324])^(a[405] & b[325])^(a[404] & b[326])^(a[403] & b[327])^(a[402] & b[328])^(a[401] & b[329])^(a[400] & b[330])^(a[399] & b[331])^(a[398] & b[332])^(a[397] & b[333])^(a[396] & b[334])^(a[395] & b[335])^(a[394] & b[336])^(a[393] & b[337])^(a[392] & b[338])^(a[391] & b[339])^(a[390] & b[340])^(a[389] & b[341])^(a[388] & b[342])^(a[387] & b[343])^(a[386] & b[344])^(a[385] & b[345])^(a[384] & b[346])^(a[383] & b[347])^(a[382] & b[348])^(a[381] & b[349])^(a[380] & b[350])^(a[379] & b[351])^(a[378] & b[352])^(a[377] & b[353])^(a[376] & b[354])^(a[375] & b[355])^(a[374] & b[356])^(a[373] & b[357])^(a[372] & b[358])^(a[371] & b[359])^(a[370] & b[360])^(a[369] & b[361])^(a[368] & b[362])^(a[367] & b[363])^(a[366] & b[364])^(a[365] & b[365])^(a[364] & b[366])^(a[363] & b[367])^(a[362] & b[368])^(a[361] & b[369])^(a[360] & b[370])^(a[359] & b[371])^(a[358] & b[372])^(a[357] & b[373])^(a[356] & b[374])^(a[355] & b[375])^(a[354] & b[376])^(a[353] & b[377])^(a[352] & b[378])^(a[351] & b[379])^(a[350] & b[380])^(a[349] & b[381])^(a[348] & b[382])^(a[347] & b[383])^(a[346] & b[384])^(a[345] & b[385])^(a[344] & b[386])^(a[343] & b[387])^(a[342] & b[388])^(a[341] & b[389])^(a[340] & b[390])^(a[339] & b[391])^(a[338] & b[392])^(a[337] & b[393])^(a[336] & b[394])^(a[335] & b[395])^(a[334] & b[396])^(a[333] & b[397])^(a[332] & b[398])^(a[331] & b[399])^(a[330] & b[400])^(a[329] & b[401])^(a[328] & b[402])^(a[327] & b[403])^(a[326] & b[404])^(a[325] & b[405])^(a[324] & b[406])^(a[323] & b[407])^(a[322] & b[408]);
assign y[731] = (a[408] & b[323])^(a[407] & b[324])^(a[406] & b[325])^(a[405] & b[326])^(a[404] & b[327])^(a[403] & b[328])^(a[402] & b[329])^(a[401] & b[330])^(a[400] & b[331])^(a[399] & b[332])^(a[398] & b[333])^(a[397] & b[334])^(a[396] & b[335])^(a[395] & b[336])^(a[394] & b[337])^(a[393] & b[338])^(a[392] & b[339])^(a[391] & b[340])^(a[390] & b[341])^(a[389] & b[342])^(a[388] & b[343])^(a[387] & b[344])^(a[386] & b[345])^(a[385] & b[346])^(a[384] & b[347])^(a[383] & b[348])^(a[382] & b[349])^(a[381] & b[350])^(a[380] & b[351])^(a[379] & b[352])^(a[378] & b[353])^(a[377] & b[354])^(a[376] & b[355])^(a[375] & b[356])^(a[374] & b[357])^(a[373] & b[358])^(a[372] & b[359])^(a[371] & b[360])^(a[370] & b[361])^(a[369] & b[362])^(a[368] & b[363])^(a[367] & b[364])^(a[366] & b[365])^(a[365] & b[366])^(a[364] & b[367])^(a[363] & b[368])^(a[362] & b[369])^(a[361] & b[370])^(a[360] & b[371])^(a[359] & b[372])^(a[358] & b[373])^(a[357] & b[374])^(a[356] & b[375])^(a[355] & b[376])^(a[354] & b[377])^(a[353] & b[378])^(a[352] & b[379])^(a[351] & b[380])^(a[350] & b[381])^(a[349] & b[382])^(a[348] & b[383])^(a[347] & b[384])^(a[346] & b[385])^(a[345] & b[386])^(a[344] & b[387])^(a[343] & b[388])^(a[342] & b[389])^(a[341] & b[390])^(a[340] & b[391])^(a[339] & b[392])^(a[338] & b[393])^(a[337] & b[394])^(a[336] & b[395])^(a[335] & b[396])^(a[334] & b[397])^(a[333] & b[398])^(a[332] & b[399])^(a[331] & b[400])^(a[330] & b[401])^(a[329] & b[402])^(a[328] & b[403])^(a[327] & b[404])^(a[326] & b[405])^(a[325] & b[406])^(a[324] & b[407])^(a[323] & b[408]);
assign y[732] = (a[408] & b[324])^(a[407] & b[325])^(a[406] & b[326])^(a[405] & b[327])^(a[404] & b[328])^(a[403] & b[329])^(a[402] & b[330])^(a[401] & b[331])^(a[400] & b[332])^(a[399] & b[333])^(a[398] & b[334])^(a[397] & b[335])^(a[396] & b[336])^(a[395] & b[337])^(a[394] & b[338])^(a[393] & b[339])^(a[392] & b[340])^(a[391] & b[341])^(a[390] & b[342])^(a[389] & b[343])^(a[388] & b[344])^(a[387] & b[345])^(a[386] & b[346])^(a[385] & b[347])^(a[384] & b[348])^(a[383] & b[349])^(a[382] & b[350])^(a[381] & b[351])^(a[380] & b[352])^(a[379] & b[353])^(a[378] & b[354])^(a[377] & b[355])^(a[376] & b[356])^(a[375] & b[357])^(a[374] & b[358])^(a[373] & b[359])^(a[372] & b[360])^(a[371] & b[361])^(a[370] & b[362])^(a[369] & b[363])^(a[368] & b[364])^(a[367] & b[365])^(a[366] & b[366])^(a[365] & b[367])^(a[364] & b[368])^(a[363] & b[369])^(a[362] & b[370])^(a[361] & b[371])^(a[360] & b[372])^(a[359] & b[373])^(a[358] & b[374])^(a[357] & b[375])^(a[356] & b[376])^(a[355] & b[377])^(a[354] & b[378])^(a[353] & b[379])^(a[352] & b[380])^(a[351] & b[381])^(a[350] & b[382])^(a[349] & b[383])^(a[348] & b[384])^(a[347] & b[385])^(a[346] & b[386])^(a[345] & b[387])^(a[344] & b[388])^(a[343] & b[389])^(a[342] & b[390])^(a[341] & b[391])^(a[340] & b[392])^(a[339] & b[393])^(a[338] & b[394])^(a[337] & b[395])^(a[336] & b[396])^(a[335] & b[397])^(a[334] & b[398])^(a[333] & b[399])^(a[332] & b[400])^(a[331] & b[401])^(a[330] & b[402])^(a[329] & b[403])^(a[328] & b[404])^(a[327] & b[405])^(a[326] & b[406])^(a[325] & b[407])^(a[324] & b[408]);
assign y[733] = (a[408] & b[325])^(a[407] & b[326])^(a[406] & b[327])^(a[405] & b[328])^(a[404] & b[329])^(a[403] & b[330])^(a[402] & b[331])^(a[401] & b[332])^(a[400] & b[333])^(a[399] & b[334])^(a[398] & b[335])^(a[397] & b[336])^(a[396] & b[337])^(a[395] & b[338])^(a[394] & b[339])^(a[393] & b[340])^(a[392] & b[341])^(a[391] & b[342])^(a[390] & b[343])^(a[389] & b[344])^(a[388] & b[345])^(a[387] & b[346])^(a[386] & b[347])^(a[385] & b[348])^(a[384] & b[349])^(a[383] & b[350])^(a[382] & b[351])^(a[381] & b[352])^(a[380] & b[353])^(a[379] & b[354])^(a[378] & b[355])^(a[377] & b[356])^(a[376] & b[357])^(a[375] & b[358])^(a[374] & b[359])^(a[373] & b[360])^(a[372] & b[361])^(a[371] & b[362])^(a[370] & b[363])^(a[369] & b[364])^(a[368] & b[365])^(a[367] & b[366])^(a[366] & b[367])^(a[365] & b[368])^(a[364] & b[369])^(a[363] & b[370])^(a[362] & b[371])^(a[361] & b[372])^(a[360] & b[373])^(a[359] & b[374])^(a[358] & b[375])^(a[357] & b[376])^(a[356] & b[377])^(a[355] & b[378])^(a[354] & b[379])^(a[353] & b[380])^(a[352] & b[381])^(a[351] & b[382])^(a[350] & b[383])^(a[349] & b[384])^(a[348] & b[385])^(a[347] & b[386])^(a[346] & b[387])^(a[345] & b[388])^(a[344] & b[389])^(a[343] & b[390])^(a[342] & b[391])^(a[341] & b[392])^(a[340] & b[393])^(a[339] & b[394])^(a[338] & b[395])^(a[337] & b[396])^(a[336] & b[397])^(a[335] & b[398])^(a[334] & b[399])^(a[333] & b[400])^(a[332] & b[401])^(a[331] & b[402])^(a[330] & b[403])^(a[329] & b[404])^(a[328] & b[405])^(a[327] & b[406])^(a[326] & b[407])^(a[325] & b[408]);
assign y[734] = (a[408] & b[326])^(a[407] & b[327])^(a[406] & b[328])^(a[405] & b[329])^(a[404] & b[330])^(a[403] & b[331])^(a[402] & b[332])^(a[401] & b[333])^(a[400] & b[334])^(a[399] & b[335])^(a[398] & b[336])^(a[397] & b[337])^(a[396] & b[338])^(a[395] & b[339])^(a[394] & b[340])^(a[393] & b[341])^(a[392] & b[342])^(a[391] & b[343])^(a[390] & b[344])^(a[389] & b[345])^(a[388] & b[346])^(a[387] & b[347])^(a[386] & b[348])^(a[385] & b[349])^(a[384] & b[350])^(a[383] & b[351])^(a[382] & b[352])^(a[381] & b[353])^(a[380] & b[354])^(a[379] & b[355])^(a[378] & b[356])^(a[377] & b[357])^(a[376] & b[358])^(a[375] & b[359])^(a[374] & b[360])^(a[373] & b[361])^(a[372] & b[362])^(a[371] & b[363])^(a[370] & b[364])^(a[369] & b[365])^(a[368] & b[366])^(a[367] & b[367])^(a[366] & b[368])^(a[365] & b[369])^(a[364] & b[370])^(a[363] & b[371])^(a[362] & b[372])^(a[361] & b[373])^(a[360] & b[374])^(a[359] & b[375])^(a[358] & b[376])^(a[357] & b[377])^(a[356] & b[378])^(a[355] & b[379])^(a[354] & b[380])^(a[353] & b[381])^(a[352] & b[382])^(a[351] & b[383])^(a[350] & b[384])^(a[349] & b[385])^(a[348] & b[386])^(a[347] & b[387])^(a[346] & b[388])^(a[345] & b[389])^(a[344] & b[390])^(a[343] & b[391])^(a[342] & b[392])^(a[341] & b[393])^(a[340] & b[394])^(a[339] & b[395])^(a[338] & b[396])^(a[337] & b[397])^(a[336] & b[398])^(a[335] & b[399])^(a[334] & b[400])^(a[333] & b[401])^(a[332] & b[402])^(a[331] & b[403])^(a[330] & b[404])^(a[329] & b[405])^(a[328] & b[406])^(a[327] & b[407])^(a[326] & b[408]);
assign y[735] = (a[408] & b[327])^(a[407] & b[328])^(a[406] & b[329])^(a[405] & b[330])^(a[404] & b[331])^(a[403] & b[332])^(a[402] & b[333])^(a[401] & b[334])^(a[400] & b[335])^(a[399] & b[336])^(a[398] & b[337])^(a[397] & b[338])^(a[396] & b[339])^(a[395] & b[340])^(a[394] & b[341])^(a[393] & b[342])^(a[392] & b[343])^(a[391] & b[344])^(a[390] & b[345])^(a[389] & b[346])^(a[388] & b[347])^(a[387] & b[348])^(a[386] & b[349])^(a[385] & b[350])^(a[384] & b[351])^(a[383] & b[352])^(a[382] & b[353])^(a[381] & b[354])^(a[380] & b[355])^(a[379] & b[356])^(a[378] & b[357])^(a[377] & b[358])^(a[376] & b[359])^(a[375] & b[360])^(a[374] & b[361])^(a[373] & b[362])^(a[372] & b[363])^(a[371] & b[364])^(a[370] & b[365])^(a[369] & b[366])^(a[368] & b[367])^(a[367] & b[368])^(a[366] & b[369])^(a[365] & b[370])^(a[364] & b[371])^(a[363] & b[372])^(a[362] & b[373])^(a[361] & b[374])^(a[360] & b[375])^(a[359] & b[376])^(a[358] & b[377])^(a[357] & b[378])^(a[356] & b[379])^(a[355] & b[380])^(a[354] & b[381])^(a[353] & b[382])^(a[352] & b[383])^(a[351] & b[384])^(a[350] & b[385])^(a[349] & b[386])^(a[348] & b[387])^(a[347] & b[388])^(a[346] & b[389])^(a[345] & b[390])^(a[344] & b[391])^(a[343] & b[392])^(a[342] & b[393])^(a[341] & b[394])^(a[340] & b[395])^(a[339] & b[396])^(a[338] & b[397])^(a[337] & b[398])^(a[336] & b[399])^(a[335] & b[400])^(a[334] & b[401])^(a[333] & b[402])^(a[332] & b[403])^(a[331] & b[404])^(a[330] & b[405])^(a[329] & b[406])^(a[328] & b[407])^(a[327] & b[408]);
assign y[736] = (a[408] & b[328])^(a[407] & b[329])^(a[406] & b[330])^(a[405] & b[331])^(a[404] & b[332])^(a[403] & b[333])^(a[402] & b[334])^(a[401] & b[335])^(a[400] & b[336])^(a[399] & b[337])^(a[398] & b[338])^(a[397] & b[339])^(a[396] & b[340])^(a[395] & b[341])^(a[394] & b[342])^(a[393] & b[343])^(a[392] & b[344])^(a[391] & b[345])^(a[390] & b[346])^(a[389] & b[347])^(a[388] & b[348])^(a[387] & b[349])^(a[386] & b[350])^(a[385] & b[351])^(a[384] & b[352])^(a[383] & b[353])^(a[382] & b[354])^(a[381] & b[355])^(a[380] & b[356])^(a[379] & b[357])^(a[378] & b[358])^(a[377] & b[359])^(a[376] & b[360])^(a[375] & b[361])^(a[374] & b[362])^(a[373] & b[363])^(a[372] & b[364])^(a[371] & b[365])^(a[370] & b[366])^(a[369] & b[367])^(a[368] & b[368])^(a[367] & b[369])^(a[366] & b[370])^(a[365] & b[371])^(a[364] & b[372])^(a[363] & b[373])^(a[362] & b[374])^(a[361] & b[375])^(a[360] & b[376])^(a[359] & b[377])^(a[358] & b[378])^(a[357] & b[379])^(a[356] & b[380])^(a[355] & b[381])^(a[354] & b[382])^(a[353] & b[383])^(a[352] & b[384])^(a[351] & b[385])^(a[350] & b[386])^(a[349] & b[387])^(a[348] & b[388])^(a[347] & b[389])^(a[346] & b[390])^(a[345] & b[391])^(a[344] & b[392])^(a[343] & b[393])^(a[342] & b[394])^(a[341] & b[395])^(a[340] & b[396])^(a[339] & b[397])^(a[338] & b[398])^(a[337] & b[399])^(a[336] & b[400])^(a[335] & b[401])^(a[334] & b[402])^(a[333] & b[403])^(a[332] & b[404])^(a[331] & b[405])^(a[330] & b[406])^(a[329] & b[407])^(a[328] & b[408]);
assign y[737] = (a[408] & b[329])^(a[407] & b[330])^(a[406] & b[331])^(a[405] & b[332])^(a[404] & b[333])^(a[403] & b[334])^(a[402] & b[335])^(a[401] & b[336])^(a[400] & b[337])^(a[399] & b[338])^(a[398] & b[339])^(a[397] & b[340])^(a[396] & b[341])^(a[395] & b[342])^(a[394] & b[343])^(a[393] & b[344])^(a[392] & b[345])^(a[391] & b[346])^(a[390] & b[347])^(a[389] & b[348])^(a[388] & b[349])^(a[387] & b[350])^(a[386] & b[351])^(a[385] & b[352])^(a[384] & b[353])^(a[383] & b[354])^(a[382] & b[355])^(a[381] & b[356])^(a[380] & b[357])^(a[379] & b[358])^(a[378] & b[359])^(a[377] & b[360])^(a[376] & b[361])^(a[375] & b[362])^(a[374] & b[363])^(a[373] & b[364])^(a[372] & b[365])^(a[371] & b[366])^(a[370] & b[367])^(a[369] & b[368])^(a[368] & b[369])^(a[367] & b[370])^(a[366] & b[371])^(a[365] & b[372])^(a[364] & b[373])^(a[363] & b[374])^(a[362] & b[375])^(a[361] & b[376])^(a[360] & b[377])^(a[359] & b[378])^(a[358] & b[379])^(a[357] & b[380])^(a[356] & b[381])^(a[355] & b[382])^(a[354] & b[383])^(a[353] & b[384])^(a[352] & b[385])^(a[351] & b[386])^(a[350] & b[387])^(a[349] & b[388])^(a[348] & b[389])^(a[347] & b[390])^(a[346] & b[391])^(a[345] & b[392])^(a[344] & b[393])^(a[343] & b[394])^(a[342] & b[395])^(a[341] & b[396])^(a[340] & b[397])^(a[339] & b[398])^(a[338] & b[399])^(a[337] & b[400])^(a[336] & b[401])^(a[335] & b[402])^(a[334] & b[403])^(a[333] & b[404])^(a[332] & b[405])^(a[331] & b[406])^(a[330] & b[407])^(a[329] & b[408]);
assign y[738] = (a[408] & b[330])^(a[407] & b[331])^(a[406] & b[332])^(a[405] & b[333])^(a[404] & b[334])^(a[403] & b[335])^(a[402] & b[336])^(a[401] & b[337])^(a[400] & b[338])^(a[399] & b[339])^(a[398] & b[340])^(a[397] & b[341])^(a[396] & b[342])^(a[395] & b[343])^(a[394] & b[344])^(a[393] & b[345])^(a[392] & b[346])^(a[391] & b[347])^(a[390] & b[348])^(a[389] & b[349])^(a[388] & b[350])^(a[387] & b[351])^(a[386] & b[352])^(a[385] & b[353])^(a[384] & b[354])^(a[383] & b[355])^(a[382] & b[356])^(a[381] & b[357])^(a[380] & b[358])^(a[379] & b[359])^(a[378] & b[360])^(a[377] & b[361])^(a[376] & b[362])^(a[375] & b[363])^(a[374] & b[364])^(a[373] & b[365])^(a[372] & b[366])^(a[371] & b[367])^(a[370] & b[368])^(a[369] & b[369])^(a[368] & b[370])^(a[367] & b[371])^(a[366] & b[372])^(a[365] & b[373])^(a[364] & b[374])^(a[363] & b[375])^(a[362] & b[376])^(a[361] & b[377])^(a[360] & b[378])^(a[359] & b[379])^(a[358] & b[380])^(a[357] & b[381])^(a[356] & b[382])^(a[355] & b[383])^(a[354] & b[384])^(a[353] & b[385])^(a[352] & b[386])^(a[351] & b[387])^(a[350] & b[388])^(a[349] & b[389])^(a[348] & b[390])^(a[347] & b[391])^(a[346] & b[392])^(a[345] & b[393])^(a[344] & b[394])^(a[343] & b[395])^(a[342] & b[396])^(a[341] & b[397])^(a[340] & b[398])^(a[339] & b[399])^(a[338] & b[400])^(a[337] & b[401])^(a[336] & b[402])^(a[335] & b[403])^(a[334] & b[404])^(a[333] & b[405])^(a[332] & b[406])^(a[331] & b[407])^(a[330] & b[408]);
assign y[739] = (a[408] & b[331])^(a[407] & b[332])^(a[406] & b[333])^(a[405] & b[334])^(a[404] & b[335])^(a[403] & b[336])^(a[402] & b[337])^(a[401] & b[338])^(a[400] & b[339])^(a[399] & b[340])^(a[398] & b[341])^(a[397] & b[342])^(a[396] & b[343])^(a[395] & b[344])^(a[394] & b[345])^(a[393] & b[346])^(a[392] & b[347])^(a[391] & b[348])^(a[390] & b[349])^(a[389] & b[350])^(a[388] & b[351])^(a[387] & b[352])^(a[386] & b[353])^(a[385] & b[354])^(a[384] & b[355])^(a[383] & b[356])^(a[382] & b[357])^(a[381] & b[358])^(a[380] & b[359])^(a[379] & b[360])^(a[378] & b[361])^(a[377] & b[362])^(a[376] & b[363])^(a[375] & b[364])^(a[374] & b[365])^(a[373] & b[366])^(a[372] & b[367])^(a[371] & b[368])^(a[370] & b[369])^(a[369] & b[370])^(a[368] & b[371])^(a[367] & b[372])^(a[366] & b[373])^(a[365] & b[374])^(a[364] & b[375])^(a[363] & b[376])^(a[362] & b[377])^(a[361] & b[378])^(a[360] & b[379])^(a[359] & b[380])^(a[358] & b[381])^(a[357] & b[382])^(a[356] & b[383])^(a[355] & b[384])^(a[354] & b[385])^(a[353] & b[386])^(a[352] & b[387])^(a[351] & b[388])^(a[350] & b[389])^(a[349] & b[390])^(a[348] & b[391])^(a[347] & b[392])^(a[346] & b[393])^(a[345] & b[394])^(a[344] & b[395])^(a[343] & b[396])^(a[342] & b[397])^(a[341] & b[398])^(a[340] & b[399])^(a[339] & b[400])^(a[338] & b[401])^(a[337] & b[402])^(a[336] & b[403])^(a[335] & b[404])^(a[334] & b[405])^(a[333] & b[406])^(a[332] & b[407])^(a[331] & b[408]);
assign y[740] = (a[408] & b[332])^(a[407] & b[333])^(a[406] & b[334])^(a[405] & b[335])^(a[404] & b[336])^(a[403] & b[337])^(a[402] & b[338])^(a[401] & b[339])^(a[400] & b[340])^(a[399] & b[341])^(a[398] & b[342])^(a[397] & b[343])^(a[396] & b[344])^(a[395] & b[345])^(a[394] & b[346])^(a[393] & b[347])^(a[392] & b[348])^(a[391] & b[349])^(a[390] & b[350])^(a[389] & b[351])^(a[388] & b[352])^(a[387] & b[353])^(a[386] & b[354])^(a[385] & b[355])^(a[384] & b[356])^(a[383] & b[357])^(a[382] & b[358])^(a[381] & b[359])^(a[380] & b[360])^(a[379] & b[361])^(a[378] & b[362])^(a[377] & b[363])^(a[376] & b[364])^(a[375] & b[365])^(a[374] & b[366])^(a[373] & b[367])^(a[372] & b[368])^(a[371] & b[369])^(a[370] & b[370])^(a[369] & b[371])^(a[368] & b[372])^(a[367] & b[373])^(a[366] & b[374])^(a[365] & b[375])^(a[364] & b[376])^(a[363] & b[377])^(a[362] & b[378])^(a[361] & b[379])^(a[360] & b[380])^(a[359] & b[381])^(a[358] & b[382])^(a[357] & b[383])^(a[356] & b[384])^(a[355] & b[385])^(a[354] & b[386])^(a[353] & b[387])^(a[352] & b[388])^(a[351] & b[389])^(a[350] & b[390])^(a[349] & b[391])^(a[348] & b[392])^(a[347] & b[393])^(a[346] & b[394])^(a[345] & b[395])^(a[344] & b[396])^(a[343] & b[397])^(a[342] & b[398])^(a[341] & b[399])^(a[340] & b[400])^(a[339] & b[401])^(a[338] & b[402])^(a[337] & b[403])^(a[336] & b[404])^(a[335] & b[405])^(a[334] & b[406])^(a[333] & b[407])^(a[332] & b[408]);
assign y[741] = (a[408] & b[333])^(a[407] & b[334])^(a[406] & b[335])^(a[405] & b[336])^(a[404] & b[337])^(a[403] & b[338])^(a[402] & b[339])^(a[401] & b[340])^(a[400] & b[341])^(a[399] & b[342])^(a[398] & b[343])^(a[397] & b[344])^(a[396] & b[345])^(a[395] & b[346])^(a[394] & b[347])^(a[393] & b[348])^(a[392] & b[349])^(a[391] & b[350])^(a[390] & b[351])^(a[389] & b[352])^(a[388] & b[353])^(a[387] & b[354])^(a[386] & b[355])^(a[385] & b[356])^(a[384] & b[357])^(a[383] & b[358])^(a[382] & b[359])^(a[381] & b[360])^(a[380] & b[361])^(a[379] & b[362])^(a[378] & b[363])^(a[377] & b[364])^(a[376] & b[365])^(a[375] & b[366])^(a[374] & b[367])^(a[373] & b[368])^(a[372] & b[369])^(a[371] & b[370])^(a[370] & b[371])^(a[369] & b[372])^(a[368] & b[373])^(a[367] & b[374])^(a[366] & b[375])^(a[365] & b[376])^(a[364] & b[377])^(a[363] & b[378])^(a[362] & b[379])^(a[361] & b[380])^(a[360] & b[381])^(a[359] & b[382])^(a[358] & b[383])^(a[357] & b[384])^(a[356] & b[385])^(a[355] & b[386])^(a[354] & b[387])^(a[353] & b[388])^(a[352] & b[389])^(a[351] & b[390])^(a[350] & b[391])^(a[349] & b[392])^(a[348] & b[393])^(a[347] & b[394])^(a[346] & b[395])^(a[345] & b[396])^(a[344] & b[397])^(a[343] & b[398])^(a[342] & b[399])^(a[341] & b[400])^(a[340] & b[401])^(a[339] & b[402])^(a[338] & b[403])^(a[337] & b[404])^(a[336] & b[405])^(a[335] & b[406])^(a[334] & b[407])^(a[333] & b[408]);
assign y[742] = (a[408] & b[334])^(a[407] & b[335])^(a[406] & b[336])^(a[405] & b[337])^(a[404] & b[338])^(a[403] & b[339])^(a[402] & b[340])^(a[401] & b[341])^(a[400] & b[342])^(a[399] & b[343])^(a[398] & b[344])^(a[397] & b[345])^(a[396] & b[346])^(a[395] & b[347])^(a[394] & b[348])^(a[393] & b[349])^(a[392] & b[350])^(a[391] & b[351])^(a[390] & b[352])^(a[389] & b[353])^(a[388] & b[354])^(a[387] & b[355])^(a[386] & b[356])^(a[385] & b[357])^(a[384] & b[358])^(a[383] & b[359])^(a[382] & b[360])^(a[381] & b[361])^(a[380] & b[362])^(a[379] & b[363])^(a[378] & b[364])^(a[377] & b[365])^(a[376] & b[366])^(a[375] & b[367])^(a[374] & b[368])^(a[373] & b[369])^(a[372] & b[370])^(a[371] & b[371])^(a[370] & b[372])^(a[369] & b[373])^(a[368] & b[374])^(a[367] & b[375])^(a[366] & b[376])^(a[365] & b[377])^(a[364] & b[378])^(a[363] & b[379])^(a[362] & b[380])^(a[361] & b[381])^(a[360] & b[382])^(a[359] & b[383])^(a[358] & b[384])^(a[357] & b[385])^(a[356] & b[386])^(a[355] & b[387])^(a[354] & b[388])^(a[353] & b[389])^(a[352] & b[390])^(a[351] & b[391])^(a[350] & b[392])^(a[349] & b[393])^(a[348] & b[394])^(a[347] & b[395])^(a[346] & b[396])^(a[345] & b[397])^(a[344] & b[398])^(a[343] & b[399])^(a[342] & b[400])^(a[341] & b[401])^(a[340] & b[402])^(a[339] & b[403])^(a[338] & b[404])^(a[337] & b[405])^(a[336] & b[406])^(a[335] & b[407])^(a[334] & b[408]);
assign y[743] = (a[408] & b[335])^(a[407] & b[336])^(a[406] & b[337])^(a[405] & b[338])^(a[404] & b[339])^(a[403] & b[340])^(a[402] & b[341])^(a[401] & b[342])^(a[400] & b[343])^(a[399] & b[344])^(a[398] & b[345])^(a[397] & b[346])^(a[396] & b[347])^(a[395] & b[348])^(a[394] & b[349])^(a[393] & b[350])^(a[392] & b[351])^(a[391] & b[352])^(a[390] & b[353])^(a[389] & b[354])^(a[388] & b[355])^(a[387] & b[356])^(a[386] & b[357])^(a[385] & b[358])^(a[384] & b[359])^(a[383] & b[360])^(a[382] & b[361])^(a[381] & b[362])^(a[380] & b[363])^(a[379] & b[364])^(a[378] & b[365])^(a[377] & b[366])^(a[376] & b[367])^(a[375] & b[368])^(a[374] & b[369])^(a[373] & b[370])^(a[372] & b[371])^(a[371] & b[372])^(a[370] & b[373])^(a[369] & b[374])^(a[368] & b[375])^(a[367] & b[376])^(a[366] & b[377])^(a[365] & b[378])^(a[364] & b[379])^(a[363] & b[380])^(a[362] & b[381])^(a[361] & b[382])^(a[360] & b[383])^(a[359] & b[384])^(a[358] & b[385])^(a[357] & b[386])^(a[356] & b[387])^(a[355] & b[388])^(a[354] & b[389])^(a[353] & b[390])^(a[352] & b[391])^(a[351] & b[392])^(a[350] & b[393])^(a[349] & b[394])^(a[348] & b[395])^(a[347] & b[396])^(a[346] & b[397])^(a[345] & b[398])^(a[344] & b[399])^(a[343] & b[400])^(a[342] & b[401])^(a[341] & b[402])^(a[340] & b[403])^(a[339] & b[404])^(a[338] & b[405])^(a[337] & b[406])^(a[336] & b[407])^(a[335] & b[408]);
assign y[744] = (a[408] & b[336])^(a[407] & b[337])^(a[406] & b[338])^(a[405] & b[339])^(a[404] & b[340])^(a[403] & b[341])^(a[402] & b[342])^(a[401] & b[343])^(a[400] & b[344])^(a[399] & b[345])^(a[398] & b[346])^(a[397] & b[347])^(a[396] & b[348])^(a[395] & b[349])^(a[394] & b[350])^(a[393] & b[351])^(a[392] & b[352])^(a[391] & b[353])^(a[390] & b[354])^(a[389] & b[355])^(a[388] & b[356])^(a[387] & b[357])^(a[386] & b[358])^(a[385] & b[359])^(a[384] & b[360])^(a[383] & b[361])^(a[382] & b[362])^(a[381] & b[363])^(a[380] & b[364])^(a[379] & b[365])^(a[378] & b[366])^(a[377] & b[367])^(a[376] & b[368])^(a[375] & b[369])^(a[374] & b[370])^(a[373] & b[371])^(a[372] & b[372])^(a[371] & b[373])^(a[370] & b[374])^(a[369] & b[375])^(a[368] & b[376])^(a[367] & b[377])^(a[366] & b[378])^(a[365] & b[379])^(a[364] & b[380])^(a[363] & b[381])^(a[362] & b[382])^(a[361] & b[383])^(a[360] & b[384])^(a[359] & b[385])^(a[358] & b[386])^(a[357] & b[387])^(a[356] & b[388])^(a[355] & b[389])^(a[354] & b[390])^(a[353] & b[391])^(a[352] & b[392])^(a[351] & b[393])^(a[350] & b[394])^(a[349] & b[395])^(a[348] & b[396])^(a[347] & b[397])^(a[346] & b[398])^(a[345] & b[399])^(a[344] & b[400])^(a[343] & b[401])^(a[342] & b[402])^(a[341] & b[403])^(a[340] & b[404])^(a[339] & b[405])^(a[338] & b[406])^(a[337] & b[407])^(a[336] & b[408]);
assign y[745] = (a[408] & b[337])^(a[407] & b[338])^(a[406] & b[339])^(a[405] & b[340])^(a[404] & b[341])^(a[403] & b[342])^(a[402] & b[343])^(a[401] & b[344])^(a[400] & b[345])^(a[399] & b[346])^(a[398] & b[347])^(a[397] & b[348])^(a[396] & b[349])^(a[395] & b[350])^(a[394] & b[351])^(a[393] & b[352])^(a[392] & b[353])^(a[391] & b[354])^(a[390] & b[355])^(a[389] & b[356])^(a[388] & b[357])^(a[387] & b[358])^(a[386] & b[359])^(a[385] & b[360])^(a[384] & b[361])^(a[383] & b[362])^(a[382] & b[363])^(a[381] & b[364])^(a[380] & b[365])^(a[379] & b[366])^(a[378] & b[367])^(a[377] & b[368])^(a[376] & b[369])^(a[375] & b[370])^(a[374] & b[371])^(a[373] & b[372])^(a[372] & b[373])^(a[371] & b[374])^(a[370] & b[375])^(a[369] & b[376])^(a[368] & b[377])^(a[367] & b[378])^(a[366] & b[379])^(a[365] & b[380])^(a[364] & b[381])^(a[363] & b[382])^(a[362] & b[383])^(a[361] & b[384])^(a[360] & b[385])^(a[359] & b[386])^(a[358] & b[387])^(a[357] & b[388])^(a[356] & b[389])^(a[355] & b[390])^(a[354] & b[391])^(a[353] & b[392])^(a[352] & b[393])^(a[351] & b[394])^(a[350] & b[395])^(a[349] & b[396])^(a[348] & b[397])^(a[347] & b[398])^(a[346] & b[399])^(a[345] & b[400])^(a[344] & b[401])^(a[343] & b[402])^(a[342] & b[403])^(a[341] & b[404])^(a[340] & b[405])^(a[339] & b[406])^(a[338] & b[407])^(a[337] & b[408]);
assign y[746] = (a[408] & b[338])^(a[407] & b[339])^(a[406] & b[340])^(a[405] & b[341])^(a[404] & b[342])^(a[403] & b[343])^(a[402] & b[344])^(a[401] & b[345])^(a[400] & b[346])^(a[399] & b[347])^(a[398] & b[348])^(a[397] & b[349])^(a[396] & b[350])^(a[395] & b[351])^(a[394] & b[352])^(a[393] & b[353])^(a[392] & b[354])^(a[391] & b[355])^(a[390] & b[356])^(a[389] & b[357])^(a[388] & b[358])^(a[387] & b[359])^(a[386] & b[360])^(a[385] & b[361])^(a[384] & b[362])^(a[383] & b[363])^(a[382] & b[364])^(a[381] & b[365])^(a[380] & b[366])^(a[379] & b[367])^(a[378] & b[368])^(a[377] & b[369])^(a[376] & b[370])^(a[375] & b[371])^(a[374] & b[372])^(a[373] & b[373])^(a[372] & b[374])^(a[371] & b[375])^(a[370] & b[376])^(a[369] & b[377])^(a[368] & b[378])^(a[367] & b[379])^(a[366] & b[380])^(a[365] & b[381])^(a[364] & b[382])^(a[363] & b[383])^(a[362] & b[384])^(a[361] & b[385])^(a[360] & b[386])^(a[359] & b[387])^(a[358] & b[388])^(a[357] & b[389])^(a[356] & b[390])^(a[355] & b[391])^(a[354] & b[392])^(a[353] & b[393])^(a[352] & b[394])^(a[351] & b[395])^(a[350] & b[396])^(a[349] & b[397])^(a[348] & b[398])^(a[347] & b[399])^(a[346] & b[400])^(a[345] & b[401])^(a[344] & b[402])^(a[343] & b[403])^(a[342] & b[404])^(a[341] & b[405])^(a[340] & b[406])^(a[339] & b[407])^(a[338] & b[408]);
assign y[747] = (a[408] & b[339])^(a[407] & b[340])^(a[406] & b[341])^(a[405] & b[342])^(a[404] & b[343])^(a[403] & b[344])^(a[402] & b[345])^(a[401] & b[346])^(a[400] & b[347])^(a[399] & b[348])^(a[398] & b[349])^(a[397] & b[350])^(a[396] & b[351])^(a[395] & b[352])^(a[394] & b[353])^(a[393] & b[354])^(a[392] & b[355])^(a[391] & b[356])^(a[390] & b[357])^(a[389] & b[358])^(a[388] & b[359])^(a[387] & b[360])^(a[386] & b[361])^(a[385] & b[362])^(a[384] & b[363])^(a[383] & b[364])^(a[382] & b[365])^(a[381] & b[366])^(a[380] & b[367])^(a[379] & b[368])^(a[378] & b[369])^(a[377] & b[370])^(a[376] & b[371])^(a[375] & b[372])^(a[374] & b[373])^(a[373] & b[374])^(a[372] & b[375])^(a[371] & b[376])^(a[370] & b[377])^(a[369] & b[378])^(a[368] & b[379])^(a[367] & b[380])^(a[366] & b[381])^(a[365] & b[382])^(a[364] & b[383])^(a[363] & b[384])^(a[362] & b[385])^(a[361] & b[386])^(a[360] & b[387])^(a[359] & b[388])^(a[358] & b[389])^(a[357] & b[390])^(a[356] & b[391])^(a[355] & b[392])^(a[354] & b[393])^(a[353] & b[394])^(a[352] & b[395])^(a[351] & b[396])^(a[350] & b[397])^(a[349] & b[398])^(a[348] & b[399])^(a[347] & b[400])^(a[346] & b[401])^(a[345] & b[402])^(a[344] & b[403])^(a[343] & b[404])^(a[342] & b[405])^(a[341] & b[406])^(a[340] & b[407])^(a[339] & b[408]);
assign y[748] = (a[408] & b[340])^(a[407] & b[341])^(a[406] & b[342])^(a[405] & b[343])^(a[404] & b[344])^(a[403] & b[345])^(a[402] & b[346])^(a[401] & b[347])^(a[400] & b[348])^(a[399] & b[349])^(a[398] & b[350])^(a[397] & b[351])^(a[396] & b[352])^(a[395] & b[353])^(a[394] & b[354])^(a[393] & b[355])^(a[392] & b[356])^(a[391] & b[357])^(a[390] & b[358])^(a[389] & b[359])^(a[388] & b[360])^(a[387] & b[361])^(a[386] & b[362])^(a[385] & b[363])^(a[384] & b[364])^(a[383] & b[365])^(a[382] & b[366])^(a[381] & b[367])^(a[380] & b[368])^(a[379] & b[369])^(a[378] & b[370])^(a[377] & b[371])^(a[376] & b[372])^(a[375] & b[373])^(a[374] & b[374])^(a[373] & b[375])^(a[372] & b[376])^(a[371] & b[377])^(a[370] & b[378])^(a[369] & b[379])^(a[368] & b[380])^(a[367] & b[381])^(a[366] & b[382])^(a[365] & b[383])^(a[364] & b[384])^(a[363] & b[385])^(a[362] & b[386])^(a[361] & b[387])^(a[360] & b[388])^(a[359] & b[389])^(a[358] & b[390])^(a[357] & b[391])^(a[356] & b[392])^(a[355] & b[393])^(a[354] & b[394])^(a[353] & b[395])^(a[352] & b[396])^(a[351] & b[397])^(a[350] & b[398])^(a[349] & b[399])^(a[348] & b[400])^(a[347] & b[401])^(a[346] & b[402])^(a[345] & b[403])^(a[344] & b[404])^(a[343] & b[405])^(a[342] & b[406])^(a[341] & b[407])^(a[340] & b[408]);
assign y[749] = (a[408] & b[341])^(a[407] & b[342])^(a[406] & b[343])^(a[405] & b[344])^(a[404] & b[345])^(a[403] & b[346])^(a[402] & b[347])^(a[401] & b[348])^(a[400] & b[349])^(a[399] & b[350])^(a[398] & b[351])^(a[397] & b[352])^(a[396] & b[353])^(a[395] & b[354])^(a[394] & b[355])^(a[393] & b[356])^(a[392] & b[357])^(a[391] & b[358])^(a[390] & b[359])^(a[389] & b[360])^(a[388] & b[361])^(a[387] & b[362])^(a[386] & b[363])^(a[385] & b[364])^(a[384] & b[365])^(a[383] & b[366])^(a[382] & b[367])^(a[381] & b[368])^(a[380] & b[369])^(a[379] & b[370])^(a[378] & b[371])^(a[377] & b[372])^(a[376] & b[373])^(a[375] & b[374])^(a[374] & b[375])^(a[373] & b[376])^(a[372] & b[377])^(a[371] & b[378])^(a[370] & b[379])^(a[369] & b[380])^(a[368] & b[381])^(a[367] & b[382])^(a[366] & b[383])^(a[365] & b[384])^(a[364] & b[385])^(a[363] & b[386])^(a[362] & b[387])^(a[361] & b[388])^(a[360] & b[389])^(a[359] & b[390])^(a[358] & b[391])^(a[357] & b[392])^(a[356] & b[393])^(a[355] & b[394])^(a[354] & b[395])^(a[353] & b[396])^(a[352] & b[397])^(a[351] & b[398])^(a[350] & b[399])^(a[349] & b[400])^(a[348] & b[401])^(a[347] & b[402])^(a[346] & b[403])^(a[345] & b[404])^(a[344] & b[405])^(a[343] & b[406])^(a[342] & b[407])^(a[341] & b[408]);
assign y[750] = (a[408] & b[342])^(a[407] & b[343])^(a[406] & b[344])^(a[405] & b[345])^(a[404] & b[346])^(a[403] & b[347])^(a[402] & b[348])^(a[401] & b[349])^(a[400] & b[350])^(a[399] & b[351])^(a[398] & b[352])^(a[397] & b[353])^(a[396] & b[354])^(a[395] & b[355])^(a[394] & b[356])^(a[393] & b[357])^(a[392] & b[358])^(a[391] & b[359])^(a[390] & b[360])^(a[389] & b[361])^(a[388] & b[362])^(a[387] & b[363])^(a[386] & b[364])^(a[385] & b[365])^(a[384] & b[366])^(a[383] & b[367])^(a[382] & b[368])^(a[381] & b[369])^(a[380] & b[370])^(a[379] & b[371])^(a[378] & b[372])^(a[377] & b[373])^(a[376] & b[374])^(a[375] & b[375])^(a[374] & b[376])^(a[373] & b[377])^(a[372] & b[378])^(a[371] & b[379])^(a[370] & b[380])^(a[369] & b[381])^(a[368] & b[382])^(a[367] & b[383])^(a[366] & b[384])^(a[365] & b[385])^(a[364] & b[386])^(a[363] & b[387])^(a[362] & b[388])^(a[361] & b[389])^(a[360] & b[390])^(a[359] & b[391])^(a[358] & b[392])^(a[357] & b[393])^(a[356] & b[394])^(a[355] & b[395])^(a[354] & b[396])^(a[353] & b[397])^(a[352] & b[398])^(a[351] & b[399])^(a[350] & b[400])^(a[349] & b[401])^(a[348] & b[402])^(a[347] & b[403])^(a[346] & b[404])^(a[345] & b[405])^(a[344] & b[406])^(a[343] & b[407])^(a[342] & b[408]);
assign y[751] = (a[408] & b[343])^(a[407] & b[344])^(a[406] & b[345])^(a[405] & b[346])^(a[404] & b[347])^(a[403] & b[348])^(a[402] & b[349])^(a[401] & b[350])^(a[400] & b[351])^(a[399] & b[352])^(a[398] & b[353])^(a[397] & b[354])^(a[396] & b[355])^(a[395] & b[356])^(a[394] & b[357])^(a[393] & b[358])^(a[392] & b[359])^(a[391] & b[360])^(a[390] & b[361])^(a[389] & b[362])^(a[388] & b[363])^(a[387] & b[364])^(a[386] & b[365])^(a[385] & b[366])^(a[384] & b[367])^(a[383] & b[368])^(a[382] & b[369])^(a[381] & b[370])^(a[380] & b[371])^(a[379] & b[372])^(a[378] & b[373])^(a[377] & b[374])^(a[376] & b[375])^(a[375] & b[376])^(a[374] & b[377])^(a[373] & b[378])^(a[372] & b[379])^(a[371] & b[380])^(a[370] & b[381])^(a[369] & b[382])^(a[368] & b[383])^(a[367] & b[384])^(a[366] & b[385])^(a[365] & b[386])^(a[364] & b[387])^(a[363] & b[388])^(a[362] & b[389])^(a[361] & b[390])^(a[360] & b[391])^(a[359] & b[392])^(a[358] & b[393])^(a[357] & b[394])^(a[356] & b[395])^(a[355] & b[396])^(a[354] & b[397])^(a[353] & b[398])^(a[352] & b[399])^(a[351] & b[400])^(a[350] & b[401])^(a[349] & b[402])^(a[348] & b[403])^(a[347] & b[404])^(a[346] & b[405])^(a[345] & b[406])^(a[344] & b[407])^(a[343] & b[408]);
assign y[752] = (a[408] & b[344])^(a[407] & b[345])^(a[406] & b[346])^(a[405] & b[347])^(a[404] & b[348])^(a[403] & b[349])^(a[402] & b[350])^(a[401] & b[351])^(a[400] & b[352])^(a[399] & b[353])^(a[398] & b[354])^(a[397] & b[355])^(a[396] & b[356])^(a[395] & b[357])^(a[394] & b[358])^(a[393] & b[359])^(a[392] & b[360])^(a[391] & b[361])^(a[390] & b[362])^(a[389] & b[363])^(a[388] & b[364])^(a[387] & b[365])^(a[386] & b[366])^(a[385] & b[367])^(a[384] & b[368])^(a[383] & b[369])^(a[382] & b[370])^(a[381] & b[371])^(a[380] & b[372])^(a[379] & b[373])^(a[378] & b[374])^(a[377] & b[375])^(a[376] & b[376])^(a[375] & b[377])^(a[374] & b[378])^(a[373] & b[379])^(a[372] & b[380])^(a[371] & b[381])^(a[370] & b[382])^(a[369] & b[383])^(a[368] & b[384])^(a[367] & b[385])^(a[366] & b[386])^(a[365] & b[387])^(a[364] & b[388])^(a[363] & b[389])^(a[362] & b[390])^(a[361] & b[391])^(a[360] & b[392])^(a[359] & b[393])^(a[358] & b[394])^(a[357] & b[395])^(a[356] & b[396])^(a[355] & b[397])^(a[354] & b[398])^(a[353] & b[399])^(a[352] & b[400])^(a[351] & b[401])^(a[350] & b[402])^(a[349] & b[403])^(a[348] & b[404])^(a[347] & b[405])^(a[346] & b[406])^(a[345] & b[407])^(a[344] & b[408]);
assign y[753] = (a[408] & b[345])^(a[407] & b[346])^(a[406] & b[347])^(a[405] & b[348])^(a[404] & b[349])^(a[403] & b[350])^(a[402] & b[351])^(a[401] & b[352])^(a[400] & b[353])^(a[399] & b[354])^(a[398] & b[355])^(a[397] & b[356])^(a[396] & b[357])^(a[395] & b[358])^(a[394] & b[359])^(a[393] & b[360])^(a[392] & b[361])^(a[391] & b[362])^(a[390] & b[363])^(a[389] & b[364])^(a[388] & b[365])^(a[387] & b[366])^(a[386] & b[367])^(a[385] & b[368])^(a[384] & b[369])^(a[383] & b[370])^(a[382] & b[371])^(a[381] & b[372])^(a[380] & b[373])^(a[379] & b[374])^(a[378] & b[375])^(a[377] & b[376])^(a[376] & b[377])^(a[375] & b[378])^(a[374] & b[379])^(a[373] & b[380])^(a[372] & b[381])^(a[371] & b[382])^(a[370] & b[383])^(a[369] & b[384])^(a[368] & b[385])^(a[367] & b[386])^(a[366] & b[387])^(a[365] & b[388])^(a[364] & b[389])^(a[363] & b[390])^(a[362] & b[391])^(a[361] & b[392])^(a[360] & b[393])^(a[359] & b[394])^(a[358] & b[395])^(a[357] & b[396])^(a[356] & b[397])^(a[355] & b[398])^(a[354] & b[399])^(a[353] & b[400])^(a[352] & b[401])^(a[351] & b[402])^(a[350] & b[403])^(a[349] & b[404])^(a[348] & b[405])^(a[347] & b[406])^(a[346] & b[407])^(a[345] & b[408]);
assign y[754] = (a[408] & b[346])^(a[407] & b[347])^(a[406] & b[348])^(a[405] & b[349])^(a[404] & b[350])^(a[403] & b[351])^(a[402] & b[352])^(a[401] & b[353])^(a[400] & b[354])^(a[399] & b[355])^(a[398] & b[356])^(a[397] & b[357])^(a[396] & b[358])^(a[395] & b[359])^(a[394] & b[360])^(a[393] & b[361])^(a[392] & b[362])^(a[391] & b[363])^(a[390] & b[364])^(a[389] & b[365])^(a[388] & b[366])^(a[387] & b[367])^(a[386] & b[368])^(a[385] & b[369])^(a[384] & b[370])^(a[383] & b[371])^(a[382] & b[372])^(a[381] & b[373])^(a[380] & b[374])^(a[379] & b[375])^(a[378] & b[376])^(a[377] & b[377])^(a[376] & b[378])^(a[375] & b[379])^(a[374] & b[380])^(a[373] & b[381])^(a[372] & b[382])^(a[371] & b[383])^(a[370] & b[384])^(a[369] & b[385])^(a[368] & b[386])^(a[367] & b[387])^(a[366] & b[388])^(a[365] & b[389])^(a[364] & b[390])^(a[363] & b[391])^(a[362] & b[392])^(a[361] & b[393])^(a[360] & b[394])^(a[359] & b[395])^(a[358] & b[396])^(a[357] & b[397])^(a[356] & b[398])^(a[355] & b[399])^(a[354] & b[400])^(a[353] & b[401])^(a[352] & b[402])^(a[351] & b[403])^(a[350] & b[404])^(a[349] & b[405])^(a[348] & b[406])^(a[347] & b[407])^(a[346] & b[408]);
assign y[755] = (a[408] & b[347])^(a[407] & b[348])^(a[406] & b[349])^(a[405] & b[350])^(a[404] & b[351])^(a[403] & b[352])^(a[402] & b[353])^(a[401] & b[354])^(a[400] & b[355])^(a[399] & b[356])^(a[398] & b[357])^(a[397] & b[358])^(a[396] & b[359])^(a[395] & b[360])^(a[394] & b[361])^(a[393] & b[362])^(a[392] & b[363])^(a[391] & b[364])^(a[390] & b[365])^(a[389] & b[366])^(a[388] & b[367])^(a[387] & b[368])^(a[386] & b[369])^(a[385] & b[370])^(a[384] & b[371])^(a[383] & b[372])^(a[382] & b[373])^(a[381] & b[374])^(a[380] & b[375])^(a[379] & b[376])^(a[378] & b[377])^(a[377] & b[378])^(a[376] & b[379])^(a[375] & b[380])^(a[374] & b[381])^(a[373] & b[382])^(a[372] & b[383])^(a[371] & b[384])^(a[370] & b[385])^(a[369] & b[386])^(a[368] & b[387])^(a[367] & b[388])^(a[366] & b[389])^(a[365] & b[390])^(a[364] & b[391])^(a[363] & b[392])^(a[362] & b[393])^(a[361] & b[394])^(a[360] & b[395])^(a[359] & b[396])^(a[358] & b[397])^(a[357] & b[398])^(a[356] & b[399])^(a[355] & b[400])^(a[354] & b[401])^(a[353] & b[402])^(a[352] & b[403])^(a[351] & b[404])^(a[350] & b[405])^(a[349] & b[406])^(a[348] & b[407])^(a[347] & b[408]);
assign y[756] = (a[408] & b[348])^(a[407] & b[349])^(a[406] & b[350])^(a[405] & b[351])^(a[404] & b[352])^(a[403] & b[353])^(a[402] & b[354])^(a[401] & b[355])^(a[400] & b[356])^(a[399] & b[357])^(a[398] & b[358])^(a[397] & b[359])^(a[396] & b[360])^(a[395] & b[361])^(a[394] & b[362])^(a[393] & b[363])^(a[392] & b[364])^(a[391] & b[365])^(a[390] & b[366])^(a[389] & b[367])^(a[388] & b[368])^(a[387] & b[369])^(a[386] & b[370])^(a[385] & b[371])^(a[384] & b[372])^(a[383] & b[373])^(a[382] & b[374])^(a[381] & b[375])^(a[380] & b[376])^(a[379] & b[377])^(a[378] & b[378])^(a[377] & b[379])^(a[376] & b[380])^(a[375] & b[381])^(a[374] & b[382])^(a[373] & b[383])^(a[372] & b[384])^(a[371] & b[385])^(a[370] & b[386])^(a[369] & b[387])^(a[368] & b[388])^(a[367] & b[389])^(a[366] & b[390])^(a[365] & b[391])^(a[364] & b[392])^(a[363] & b[393])^(a[362] & b[394])^(a[361] & b[395])^(a[360] & b[396])^(a[359] & b[397])^(a[358] & b[398])^(a[357] & b[399])^(a[356] & b[400])^(a[355] & b[401])^(a[354] & b[402])^(a[353] & b[403])^(a[352] & b[404])^(a[351] & b[405])^(a[350] & b[406])^(a[349] & b[407])^(a[348] & b[408]);
assign y[757] = (a[408] & b[349])^(a[407] & b[350])^(a[406] & b[351])^(a[405] & b[352])^(a[404] & b[353])^(a[403] & b[354])^(a[402] & b[355])^(a[401] & b[356])^(a[400] & b[357])^(a[399] & b[358])^(a[398] & b[359])^(a[397] & b[360])^(a[396] & b[361])^(a[395] & b[362])^(a[394] & b[363])^(a[393] & b[364])^(a[392] & b[365])^(a[391] & b[366])^(a[390] & b[367])^(a[389] & b[368])^(a[388] & b[369])^(a[387] & b[370])^(a[386] & b[371])^(a[385] & b[372])^(a[384] & b[373])^(a[383] & b[374])^(a[382] & b[375])^(a[381] & b[376])^(a[380] & b[377])^(a[379] & b[378])^(a[378] & b[379])^(a[377] & b[380])^(a[376] & b[381])^(a[375] & b[382])^(a[374] & b[383])^(a[373] & b[384])^(a[372] & b[385])^(a[371] & b[386])^(a[370] & b[387])^(a[369] & b[388])^(a[368] & b[389])^(a[367] & b[390])^(a[366] & b[391])^(a[365] & b[392])^(a[364] & b[393])^(a[363] & b[394])^(a[362] & b[395])^(a[361] & b[396])^(a[360] & b[397])^(a[359] & b[398])^(a[358] & b[399])^(a[357] & b[400])^(a[356] & b[401])^(a[355] & b[402])^(a[354] & b[403])^(a[353] & b[404])^(a[352] & b[405])^(a[351] & b[406])^(a[350] & b[407])^(a[349] & b[408]);
assign y[758] = (a[408] & b[350])^(a[407] & b[351])^(a[406] & b[352])^(a[405] & b[353])^(a[404] & b[354])^(a[403] & b[355])^(a[402] & b[356])^(a[401] & b[357])^(a[400] & b[358])^(a[399] & b[359])^(a[398] & b[360])^(a[397] & b[361])^(a[396] & b[362])^(a[395] & b[363])^(a[394] & b[364])^(a[393] & b[365])^(a[392] & b[366])^(a[391] & b[367])^(a[390] & b[368])^(a[389] & b[369])^(a[388] & b[370])^(a[387] & b[371])^(a[386] & b[372])^(a[385] & b[373])^(a[384] & b[374])^(a[383] & b[375])^(a[382] & b[376])^(a[381] & b[377])^(a[380] & b[378])^(a[379] & b[379])^(a[378] & b[380])^(a[377] & b[381])^(a[376] & b[382])^(a[375] & b[383])^(a[374] & b[384])^(a[373] & b[385])^(a[372] & b[386])^(a[371] & b[387])^(a[370] & b[388])^(a[369] & b[389])^(a[368] & b[390])^(a[367] & b[391])^(a[366] & b[392])^(a[365] & b[393])^(a[364] & b[394])^(a[363] & b[395])^(a[362] & b[396])^(a[361] & b[397])^(a[360] & b[398])^(a[359] & b[399])^(a[358] & b[400])^(a[357] & b[401])^(a[356] & b[402])^(a[355] & b[403])^(a[354] & b[404])^(a[353] & b[405])^(a[352] & b[406])^(a[351] & b[407])^(a[350] & b[408]);
assign y[759] = (a[408] & b[351])^(a[407] & b[352])^(a[406] & b[353])^(a[405] & b[354])^(a[404] & b[355])^(a[403] & b[356])^(a[402] & b[357])^(a[401] & b[358])^(a[400] & b[359])^(a[399] & b[360])^(a[398] & b[361])^(a[397] & b[362])^(a[396] & b[363])^(a[395] & b[364])^(a[394] & b[365])^(a[393] & b[366])^(a[392] & b[367])^(a[391] & b[368])^(a[390] & b[369])^(a[389] & b[370])^(a[388] & b[371])^(a[387] & b[372])^(a[386] & b[373])^(a[385] & b[374])^(a[384] & b[375])^(a[383] & b[376])^(a[382] & b[377])^(a[381] & b[378])^(a[380] & b[379])^(a[379] & b[380])^(a[378] & b[381])^(a[377] & b[382])^(a[376] & b[383])^(a[375] & b[384])^(a[374] & b[385])^(a[373] & b[386])^(a[372] & b[387])^(a[371] & b[388])^(a[370] & b[389])^(a[369] & b[390])^(a[368] & b[391])^(a[367] & b[392])^(a[366] & b[393])^(a[365] & b[394])^(a[364] & b[395])^(a[363] & b[396])^(a[362] & b[397])^(a[361] & b[398])^(a[360] & b[399])^(a[359] & b[400])^(a[358] & b[401])^(a[357] & b[402])^(a[356] & b[403])^(a[355] & b[404])^(a[354] & b[405])^(a[353] & b[406])^(a[352] & b[407])^(a[351] & b[408]);
assign y[760] = (a[408] & b[352])^(a[407] & b[353])^(a[406] & b[354])^(a[405] & b[355])^(a[404] & b[356])^(a[403] & b[357])^(a[402] & b[358])^(a[401] & b[359])^(a[400] & b[360])^(a[399] & b[361])^(a[398] & b[362])^(a[397] & b[363])^(a[396] & b[364])^(a[395] & b[365])^(a[394] & b[366])^(a[393] & b[367])^(a[392] & b[368])^(a[391] & b[369])^(a[390] & b[370])^(a[389] & b[371])^(a[388] & b[372])^(a[387] & b[373])^(a[386] & b[374])^(a[385] & b[375])^(a[384] & b[376])^(a[383] & b[377])^(a[382] & b[378])^(a[381] & b[379])^(a[380] & b[380])^(a[379] & b[381])^(a[378] & b[382])^(a[377] & b[383])^(a[376] & b[384])^(a[375] & b[385])^(a[374] & b[386])^(a[373] & b[387])^(a[372] & b[388])^(a[371] & b[389])^(a[370] & b[390])^(a[369] & b[391])^(a[368] & b[392])^(a[367] & b[393])^(a[366] & b[394])^(a[365] & b[395])^(a[364] & b[396])^(a[363] & b[397])^(a[362] & b[398])^(a[361] & b[399])^(a[360] & b[400])^(a[359] & b[401])^(a[358] & b[402])^(a[357] & b[403])^(a[356] & b[404])^(a[355] & b[405])^(a[354] & b[406])^(a[353] & b[407])^(a[352] & b[408]);
assign y[761] = (a[408] & b[353])^(a[407] & b[354])^(a[406] & b[355])^(a[405] & b[356])^(a[404] & b[357])^(a[403] & b[358])^(a[402] & b[359])^(a[401] & b[360])^(a[400] & b[361])^(a[399] & b[362])^(a[398] & b[363])^(a[397] & b[364])^(a[396] & b[365])^(a[395] & b[366])^(a[394] & b[367])^(a[393] & b[368])^(a[392] & b[369])^(a[391] & b[370])^(a[390] & b[371])^(a[389] & b[372])^(a[388] & b[373])^(a[387] & b[374])^(a[386] & b[375])^(a[385] & b[376])^(a[384] & b[377])^(a[383] & b[378])^(a[382] & b[379])^(a[381] & b[380])^(a[380] & b[381])^(a[379] & b[382])^(a[378] & b[383])^(a[377] & b[384])^(a[376] & b[385])^(a[375] & b[386])^(a[374] & b[387])^(a[373] & b[388])^(a[372] & b[389])^(a[371] & b[390])^(a[370] & b[391])^(a[369] & b[392])^(a[368] & b[393])^(a[367] & b[394])^(a[366] & b[395])^(a[365] & b[396])^(a[364] & b[397])^(a[363] & b[398])^(a[362] & b[399])^(a[361] & b[400])^(a[360] & b[401])^(a[359] & b[402])^(a[358] & b[403])^(a[357] & b[404])^(a[356] & b[405])^(a[355] & b[406])^(a[354] & b[407])^(a[353] & b[408]);
assign y[762] = (a[408] & b[354])^(a[407] & b[355])^(a[406] & b[356])^(a[405] & b[357])^(a[404] & b[358])^(a[403] & b[359])^(a[402] & b[360])^(a[401] & b[361])^(a[400] & b[362])^(a[399] & b[363])^(a[398] & b[364])^(a[397] & b[365])^(a[396] & b[366])^(a[395] & b[367])^(a[394] & b[368])^(a[393] & b[369])^(a[392] & b[370])^(a[391] & b[371])^(a[390] & b[372])^(a[389] & b[373])^(a[388] & b[374])^(a[387] & b[375])^(a[386] & b[376])^(a[385] & b[377])^(a[384] & b[378])^(a[383] & b[379])^(a[382] & b[380])^(a[381] & b[381])^(a[380] & b[382])^(a[379] & b[383])^(a[378] & b[384])^(a[377] & b[385])^(a[376] & b[386])^(a[375] & b[387])^(a[374] & b[388])^(a[373] & b[389])^(a[372] & b[390])^(a[371] & b[391])^(a[370] & b[392])^(a[369] & b[393])^(a[368] & b[394])^(a[367] & b[395])^(a[366] & b[396])^(a[365] & b[397])^(a[364] & b[398])^(a[363] & b[399])^(a[362] & b[400])^(a[361] & b[401])^(a[360] & b[402])^(a[359] & b[403])^(a[358] & b[404])^(a[357] & b[405])^(a[356] & b[406])^(a[355] & b[407])^(a[354] & b[408]);
assign y[763] = (a[408] & b[355])^(a[407] & b[356])^(a[406] & b[357])^(a[405] & b[358])^(a[404] & b[359])^(a[403] & b[360])^(a[402] & b[361])^(a[401] & b[362])^(a[400] & b[363])^(a[399] & b[364])^(a[398] & b[365])^(a[397] & b[366])^(a[396] & b[367])^(a[395] & b[368])^(a[394] & b[369])^(a[393] & b[370])^(a[392] & b[371])^(a[391] & b[372])^(a[390] & b[373])^(a[389] & b[374])^(a[388] & b[375])^(a[387] & b[376])^(a[386] & b[377])^(a[385] & b[378])^(a[384] & b[379])^(a[383] & b[380])^(a[382] & b[381])^(a[381] & b[382])^(a[380] & b[383])^(a[379] & b[384])^(a[378] & b[385])^(a[377] & b[386])^(a[376] & b[387])^(a[375] & b[388])^(a[374] & b[389])^(a[373] & b[390])^(a[372] & b[391])^(a[371] & b[392])^(a[370] & b[393])^(a[369] & b[394])^(a[368] & b[395])^(a[367] & b[396])^(a[366] & b[397])^(a[365] & b[398])^(a[364] & b[399])^(a[363] & b[400])^(a[362] & b[401])^(a[361] & b[402])^(a[360] & b[403])^(a[359] & b[404])^(a[358] & b[405])^(a[357] & b[406])^(a[356] & b[407])^(a[355] & b[408]);
assign y[764] = (a[408] & b[356])^(a[407] & b[357])^(a[406] & b[358])^(a[405] & b[359])^(a[404] & b[360])^(a[403] & b[361])^(a[402] & b[362])^(a[401] & b[363])^(a[400] & b[364])^(a[399] & b[365])^(a[398] & b[366])^(a[397] & b[367])^(a[396] & b[368])^(a[395] & b[369])^(a[394] & b[370])^(a[393] & b[371])^(a[392] & b[372])^(a[391] & b[373])^(a[390] & b[374])^(a[389] & b[375])^(a[388] & b[376])^(a[387] & b[377])^(a[386] & b[378])^(a[385] & b[379])^(a[384] & b[380])^(a[383] & b[381])^(a[382] & b[382])^(a[381] & b[383])^(a[380] & b[384])^(a[379] & b[385])^(a[378] & b[386])^(a[377] & b[387])^(a[376] & b[388])^(a[375] & b[389])^(a[374] & b[390])^(a[373] & b[391])^(a[372] & b[392])^(a[371] & b[393])^(a[370] & b[394])^(a[369] & b[395])^(a[368] & b[396])^(a[367] & b[397])^(a[366] & b[398])^(a[365] & b[399])^(a[364] & b[400])^(a[363] & b[401])^(a[362] & b[402])^(a[361] & b[403])^(a[360] & b[404])^(a[359] & b[405])^(a[358] & b[406])^(a[357] & b[407])^(a[356] & b[408]);
assign y[765] = (a[408] & b[357])^(a[407] & b[358])^(a[406] & b[359])^(a[405] & b[360])^(a[404] & b[361])^(a[403] & b[362])^(a[402] & b[363])^(a[401] & b[364])^(a[400] & b[365])^(a[399] & b[366])^(a[398] & b[367])^(a[397] & b[368])^(a[396] & b[369])^(a[395] & b[370])^(a[394] & b[371])^(a[393] & b[372])^(a[392] & b[373])^(a[391] & b[374])^(a[390] & b[375])^(a[389] & b[376])^(a[388] & b[377])^(a[387] & b[378])^(a[386] & b[379])^(a[385] & b[380])^(a[384] & b[381])^(a[383] & b[382])^(a[382] & b[383])^(a[381] & b[384])^(a[380] & b[385])^(a[379] & b[386])^(a[378] & b[387])^(a[377] & b[388])^(a[376] & b[389])^(a[375] & b[390])^(a[374] & b[391])^(a[373] & b[392])^(a[372] & b[393])^(a[371] & b[394])^(a[370] & b[395])^(a[369] & b[396])^(a[368] & b[397])^(a[367] & b[398])^(a[366] & b[399])^(a[365] & b[400])^(a[364] & b[401])^(a[363] & b[402])^(a[362] & b[403])^(a[361] & b[404])^(a[360] & b[405])^(a[359] & b[406])^(a[358] & b[407])^(a[357] & b[408]);
assign y[766] = (a[408] & b[358])^(a[407] & b[359])^(a[406] & b[360])^(a[405] & b[361])^(a[404] & b[362])^(a[403] & b[363])^(a[402] & b[364])^(a[401] & b[365])^(a[400] & b[366])^(a[399] & b[367])^(a[398] & b[368])^(a[397] & b[369])^(a[396] & b[370])^(a[395] & b[371])^(a[394] & b[372])^(a[393] & b[373])^(a[392] & b[374])^(a[391] & b[375])^(a[390] & b[376])^(a[389] & b[377])^(a[388] & b[378])^(a[387] & b[379])^(a[386] & b[380])^(a[385] & b[381])^(a[384] & b[382])^(a[383] & b[383])^(a[382] & b[384])^(a[381] & b[385])^(a[380] & b[386])^(a[379] & b[387])^(a[378] & b[388])^(a[377] & b[389])^(a[376] & b[390])^(a[375] & b[391])^(a[374] & b[392])^(a[373] & b[393])^(a[372] & b[394])^(a[371] & b[395])^(a[370] & b[396])^(a[369] & b[397])^(a[368] & b[398])^(a[367] & b[399])^(a[366] & b[400])^(a[365] & b[401])^(a[364] & b[402])^(a[363] & b[403])^(a[362] & b[404])^(a[361] & b[405])^(a[360] & b[406])^(a[359] & b[407])^(a[358] & b[408]);
assign y[767] = (a[408] & b[359])^(a[407] & b[360])^(a[406] & b[361])^(a[405] & b[362])^(a[404] & b[363])^(a[403] & b[364])^(a[402] & b[365])^(a[401] & b[366])^(a[400] & b[367])^(a[399] & b[368])^(a[398] & b[369])^(a[397] & b[370])^(a[396] & b[371])^(a[395] & b[372])^(a[394] & b[373])^(a[393] & b[374])^(a[392] & b[375])^(a[391] & b[376])^(a[390] & b[377])^(a[389] & b[378])^(a[388] & b[379])^(a[387] & b[380])^(a[386] & b[381])^(a[385] & b[382])^(a[384] & b[383])^(a[383] & b[384])^(a[382] & b[385])^(a[381] & b[386])^(a[380] & b[387])^(a[379] & b[388])^(a[378] & b[389])^(a[377] & b[390])^(a[376] & b[391])^(a[375] & b[392])^(a[374] & b[393])^(a[373] & b[394])^(a[372] & b[395])^(a[371] & b[396])^(a[370] & b[397])^(a[369] & b[398])^(a[368] & b[399])^(a[367] & b[400])^(a[366] & b[401])^(a[365] & b[402])^(a[364] & b[403])^(a[363] & b[404])^(a[362] & b[405])^(a[361] & b[406])^(a[360] & b[407])^(a[359] & b[408]);
assign y[768] = (a[408] & b[360])^(a[407] & b[361])^(a[406] & b[362])^(a[405] & b[363])^(a[404] & b[364])^(a[403] & b[365])^(a[402] & b[366])^(a[401] & b[367])^(a[400] & b[368])^(a[399] & b[369])^(a[398] & b[370])^(a[397] & b[371])^(a[396] & b[372])^(a[395] & b[373])^(a[394] & b[374])^(a[393] & b[375])^(a[392] & b[376])^(a[391] & b[377])^(a[390] & b[378])^(a[389] & b[379])^(a[388] & b[380])^(a[387] & b[381])^(a[386] & b[382])^(a[385] & b[383])^(a[384] & b[384])^(a[383] & b[385])^(a[382] & b[386])^(a[381] & b[387])^(a[380] & b[388])^(a[379] & b[389])^(a[378] & b[390])^(a[377] & b[391])^(a[376] & b[392])^(a[375] & b[393])^(a[374] & b[394])^(a[373] & b[395])^(a[372] & b[396])^(a[371] & b[397])^(a[370] & b[398])^(a[369] & b[399])^(a[368] & b[400])^(a[367] & b[401])^(a[366] & b[402])^(a[365] & b[403])^(a[364] & b[404])^(a[363] & b[405])^(a[362] & b[406])^(a[361] & b[407])^(a[360] & b[408]);
assign y[769] = (a[408] & b[361])^(a[407] & b[362])^(a[406] & b[363])^(a[405] & b[364])^(a[404] & b[365])^(a[403] & b[366])^(a[402] & b[367])^(a[401] & b[368])^(a[400] & b[369])^(a[399] & b[370])^(a[398] & b[371])^(a[397] & b[372])^(a[396] & b[373])^(a[395] & b[374])^(a[394] & b[375])^(a[393] & b[376])^(a[392] & b[377])^(a[391] & b[378])^(a[390] & b[379])^(a[389] & b[380])^(a[388] & b[381])^(a[387] & b[382])^(a[386] & b[383])^(a[385] & b[384])^(a[384] & b[385])^(a[383] & b[386])^(a[382] & b[387])^(a[381] & b[388])^(a[380] & b[389])^(a[379] & b[390])^(a[378] & b[391])^(a[377] & b[392])^(a[376] & b[393])^(a[375] & b[394])^(a[374] & b[395])^(a[373] & b[396])^(a[372] & b[397])^(a[371] & b[398])^(a[370] & b[399])^(a[369] & b[400])^(a[368] & b[401])^(a[367] & b[402])^(a[366] & b[403])^(a[365] & b[404])^(a[364] & b[405])^(a[363] & b[406])^(a[362] & b[407])^(a[361] & b[408]);
assign y[770] = (a[408] & b[362])^(a[407] & b[363])^(a[406] & b[364])^(a[405] & b[365])^(a[404] & b[366])^(a[403] & b[367])^(a[402] & b[368])^(a[401] & b[369])^(a[400] & b[370])^(a[399] & b[371])^(a[398] & b[372])^(a[397] & b[373])^(a[396] & b[374])^(a[395] & b[375])^(a[394] & b[376])^(a[393] & b[377])^(a[392] & b[378])^(a[391] & b[379])^(a[390] & b[380])^(a[389] & b[381])^(a[388] & b[382])^(a[387] & b[383])^(a[386] & b[384])^(a[385] & b[385])^(a[384] & b[386])^(a[383] & b[387])^(a[382] & b[388])^(a[381] & b[389])^(a[380] & b[390])^(a[379] & b[391])^(a[378] & b[392])^(a[377] & b[393])^(a[376] & b[394])^(a[375] & b[395])^(a[374] & b[396])^(a[373] & b[397])^(a[372] & b[398])^(a[371] & b[399])^(a[370] & b[400])^(a[369] & b[401])^(a[368] & b[402])^(a[367] & b[403])^(a[366] & b[404])^(a[365] & b[405])^(a[364] & b[406])^(a[363] & b[407])^(a[362] & b[408]);
assign y[771] = (a[408] & b[363])^(a[407] & b[364])^(a[406] & b[365])^(a[405] & b[366])^(a[404] & b[367])^(a[403] & b[368])^(a[402] & b[369])^(a[401] & b[370])^(a[400] & b[371])^(a[399] & b[372])^(a[398] & b[373])^(a[397] & b[374])^(a[396] & b[375])^(a[395] & b[376])^(a[394] & b[377])^(a[393] & b[378])^(a[392] & b[379])^(a[391] & b[380])^(a[390] & b[381])^(a[389] & b[382])^(a[388] & b[383])^(a[387] & b[384])^(a[386] & b[385])^(a[385] & b[386])^(a[384] & b[387])^(a[383] & b[388])^(a[382] & b[389])^(a[381] & b[390])^(a[380] & b[391])^(a[379] & b[392])^(a[378] & b[393])^(a[377] & b[394])^(a[376] & b[395])^(a[375] & b[396])^(a[374] & b[397])^(a[373] & b[398])^(a[372] & b[399])^(a[371] & b[400])^(a[370] & b[401])^(a[369] & b[402])^(a[368] & b[403])^(a[367] & b[404])^(a[366] & b[405])^(a[365] & b[406])^(a[364] & b[407])^(a[363] & b[408]);
assign y[772] = (a[408] & b[364])^(a[407] & b[365])^(a[406] & b[366])^(a[405] & b[367])^(a[404] & b[368])^(a[403] & b[369])^(a[402] & b[370])^(a[401] & b[371])^(a[400] & b[372])^(a[399] & b[373])^(a[398] & b[374])^(a[397] & b[375])^(a[396] & b[376])^(a[395] & b[377])^(a[394] & b[378])^(a[393] & b[379])^(a[392] & b[380])^(a[391] & b[381])^(a[390] & b[382])^(a[389] & b[383])^(a[388] & b[384])^(a[387] & b[385])^(a[386] & b[386])^(a[385] & b[387])^(a[384] & b[388])^(a[383] & b[389])^(a[382] & b[390])^(a[381] & b[391])^(a[380] & b[392])^(a[379] & b[393])^(a[378] & b[394])^(a[377] & b[395])^(a[376] & b[396])^(a[375] & b[397])^(a[374] & b[398])^(a[373] & b[399])^(a[372] & b[400])^(a[371] & b[401])^(a[370] & b[402])^(a[369] & b[403])^(a[368] & b[404])^(a[367] & b[405])^(a[366] & b[406])^(a[365] & b[407])^(a[364] & b[408]);
assign y[773] = (a[408] & b[365])^(a[407] & b[366])^(a[406] & b[367])^(a[405] & b[368])^(a[404] & b[369])^(a[403] & b[370])^(a[402] & b[371])^(a[401] & b[372])^(a[400] & b[373])^(a[399] & b[374])^(a[398] & b[375])^(a[397] & b[376])^(a[396] & b[377])^(a[395] & b[378])^(a[394] & b[379])^(a[393] & b[380])^(a[392] & b[381])^(a[391] & b[382])^(a[390] & b[383])^(a[389] & b[384])^(a[388] & b[385])^(a[387] & b[386])^(a[386] & b[387])^(a[385] & b[388])^(a[384] & b[389])^(a[383] & b[390])^(a[382] & b[391])^(a[381] & b[392])^(a[380] & b[393])^(a[379] & b[394])^(a[378] & b[395])^(a[377] & b[396])^(a[376] & b[397])^(a[375] & b[398])^(a[374] & b[399])^(a[373] & b[400])^(a[372] & b[401])^(a[371] & b[402])^(a[370] & b[403])^(a[369] & b[404])^(a[368] & b[405])^(a[367] & b[406])^(a[366] & b[407])^(a[365] & b[408]);
assign y[774] = (a[408] & b[366])^(a[407] & b[367])^(a[406] & b[368])^(a[405] & b[369])^(a[404] & b[370])^(a[403] & b[371])^(a[402] & b[372])^(a[401] & b[373])^(a[400] & b[374])^(a[399] & b[375])^(a[398] & b[376])^(a[397] & b[377])^(a[396] & b[378])^(a[395] & b[379])^(a[394] & b[380])^(a[393] & b[381])^(a[392] & b[382])^(a[391] & b[383])^(a[390] & b[384])^(a[389] & b[385])^(a[388] & b[386])^(a[387] & b[387])^(a[386] & b[388])^(a[385] & b[389])^(a[384] & b[390])^(a[383] & b[391])^(a[382] & b[392])^(a[381] & b[393])^(a[380] & b[394])^(a[379] & b[395])^(a[378] & b[396])^(a[377] & b[397])^(a[376] & b[398])^(a[375] & b[399])^(a[374] & b[400])^(a[373] & b[401])^(a[372] & b[402])^(a[371] & b[403])^(a[370] & b[404])^(a[369] & b[405])^(a[368] & b[406])^(a[367] & b[407])^(a[366] & b[408]);
assign y[775] = (a[408] & b[367])^(a[407] & b[368])^(a[406] & b[369])^(a[405] & b[370])^(a[404] & b[371])^(a[403] & b[372])^(a[402] & b[373])^(a[401] & b[374])^(a[400] & b[375])^(a[399] & b[376])^(a[398] & b[377])^(a[397] & b[378])^(a[396] & b[379])^(a[395] & b[380])^(a[394] & b[381])^(a[393] & b[382])^(a[392] & b[383])^(a[391] & b[384])^(a[390] & b[385])^(a[389] & b[386])^(a[388] & b[387])^(a[387] & b[388])^(a[386] & b[389])^(a[385] & b[390])^(a[384] & b[391])^(a[383] & b[392])^(a[382] & b[393])^(a[381] & b[394])^(a[380] & b[395])^(a[379] & b[396])^(a[378] & b[397])^(a[377] & b[398])^(a[376] & b[399])^(a[375] & b[400])^(a[374] & b[401])^(a[373] & b[402])^(a[372] & b[403])^(a[371] & b[404])^(a[370] & b[405])^(a[369] & b[406])^(a[368] & b[407])^(a[367] & b[408]);
assign y[776] = (a[408] & b[368])^(a[407] & b[369])^(a[406] & b[370])^(a[405] & b[371])^(a[404] & b[372])^(a[403] & b[373])^(a[402] & b[374])^(a[401] & b[375])^(a[400] & b[376])^(a[399] & b[377])^(a[398] & b[378])^(a[397] & b[379])^(a[396] & b[380])^(a[395] & b[381])^(a[394] & b[382])^(a[393] & b[383])^(a[392] & b[384])^(a[391] & b[385])^(a[390] & b[386])^(a[389] & b[387])^(a[388] & b[388])^(a[387] & b[389])^(a[386] & b[390])^(a[385] & b[391])^(a[384] & b[392])^(a[383] & b[393])^(a[382] & b[394])^(a[381] & b[395])^(a[380] & b[396])^(a[379] & b[397])^(a[378] & b[398])^(a[377] & b[399])^(a[376] & b[400])^(a[375] & b[401])^(a[374] & b[402])^(a[373] & b[403])^(a[372] & b[404])^(a[371] & b[405])^(a[370] & b[406])^(a[369] & b[407])^(a[368] & b[408]);
assign y[777] = (a[408] & b[369])^(a[407] & b[370])^(a[406] & b[371])^(a[405] & b[372])^(a[404] & b[373])^(a[403] & b[374])^(a[402] & b[375])^(a[401] & b[376])^(a[400] & b[377])^(a[399] & b[378])^(a[398] & b[379])^(a[397] & b[380])^(a[396] & b[381])^(a[395] & b[382])^(a[394] & b[383])^(a[393] & b[384])^(a[392] & b[385])^(a[391] & b[386])^(a[390] & b[387])^(a[389] & b[388])^(a[388] & b[389])^(a[387] & b[390])^(a[386] & b[391])^(a[385] & b[392])^(a[384] & b[393])^(a[383] & b[394])^(a[382] & b[395])^(a[381] & b[396])^(a[380] & b[397])^(a[379] & b[398])^(a[378] & b[399])^(a[377] & b[400])^(a[376] & b[401])^(a[375] & b[402])^(a[374] & b[403])^(a[373] & b[404])^(a[372] & b[405])^(a[371] & b[406])^(a[370] & b[407])^(a[369] & b[408]);
assign y[778] = (a[408] & b[370])^(a[407] & b[371])^(a[406] & b[372])^(a[405] & b[373])^(a[404] & b[374])^(a[403] & b[375])^(a[402] & b[376])^(a[401] & b[377])^(a[400] & b[378])^(a[399] & b[379])^(a[398] & b[380])^(a[397] & b[381])^(a[396] & b[382])^(a[395] & b[383])^(a[394] & b[384])^(a[393] & b[385])^(a[392] & b[386])^(a[391] & b[387])^(a[390] & b[388])^(a[389] & b[389])^(a[388] & b[390])^(a[387] & b[391])^(a[386] & b[392])^(a[385] & b[393])^(a[384] & b[394])^(a[383] & b[395])^(a[382] & b[396])^(a[381] & b[397])^(a[380] & b[398])^(a[379] & b[399])^(a[378] & b[400])^(a[377] & b[401])^(a[376] & b[402])^(a[375] & b[403])^(a[374] & b[404])^(a[373] & b[405])^(a[372] & b[406])^(a[371] & b[407])^(a[370] & b[408]);
assign y[779] = (a[408] & b[371])^(a[407] & b[372])^(a[406] & b[373])^(a[405] & b[374])^(a[404] & b[375])^(a[403] & b[376])^(a[402] & b[377])^(a[401] & b[378])^(a[400] & b[379])^(a[399] & b[380])^(a[398] & b[381])^(a[397] & b[382])^(a[396] & b[383])^(a[395] & b[384])^(a[394] & b[385])^(a[393] & b[386])^(a[392] & b[387])^(a[391] & b[388])^(a[390] & b[389])^(a[389] & b[390])^(a[388] & b[391])^(a[387] & b[392])^(a[386] & b[393])^(a[385] & b[394])^(a[384] & b[395])^(a[383] & b[396])^(a[382] & b[397])^(a[381] & b[398])^(a[380] & b[399])^(a[379] & b[400])^(a[378] & b[401])^(a[377] & b[402])^(a[376] & b[403])^(a[375] & b[404])^(a[374] & b[405])^(a[373] & b[406])^(a[372] & b[407])^(a[371] & b[408]);
assign y[780] = (a[408] & b[372])^(a[407] & b[373])^(a[406] & b[374])^(a[405] & b[375])^(a[404] & b[376])^(a[403] & b[377])^(a[402] & b[378])^(a[401] & b[379])^(a[400] & b[380])^(a[399] & b[381])^(a[398] & b[382])^(a[397] & b[383])^(a[396] & b[384])^(a[395] & b[385])^(a[394] & b[386])^(a[393] & b[387])^(a[392] & b[388])^(a[391] & b[389])^(a[390] & b[390])^(a[389] & b[391])^(a[388] & b[392])^(a[387] & b[393])^(a[386] & b[394])^(a[385] & b[395])^(a[384] & b[396])^(a[383] & b[397])^(a[382] & b[398])^(a[381] & b[399])^(a[380] & b[400])^(a[379] & b[401])^(a[378] & b[402])^(a[377] & b[403])^(a[376] & b[404])^(a[375] & b[405])^(a[374] & b[406])^(a[373] & b[407])^(a[372] & b[408]);
assign y[781] = (a[408] & b[373])^(a[407] & b[374])^(a[406] & b[375])^(a[405] & b[376])^(a[404] & b[377])^(a[403] & b[378])^(a[402] & b[379])^(a[401] & b[380])^(a[400] & b[381])^(a[399] & b[382])^(a[398] & b[383])^(a[397] & b[384])^(a[396] & b[385])^(a[395] & b[386])^(a[394] & b[387])^(a[393] & b[388])^(a[392] & b[389])^(a[391] & b[390])^(a[390] & b[391])^(a[389] & b[392])^(a[388] & b[393])^(a[387] & b[394])^(a[386] & b[395])^(a[385] & b[396])^(a[384] & b[397])^(a[383] & b[398])^(a[382] & b[399])^(a[381] & b[400])^(a[380] & b[401])^(a[379] & b[402])^(a[378] & b[403])^(a[377] & b[404])^(a[376] & b[405])^(a[375] & b[406])^(a[374] & b[407])^(a[373] & b[408]);
assign y[782] = (a[408] & b[374])^(a[407] & b[375])^(a[406] & b[376])^(a[405] & b[377])^(a[404] & b[378])^(a[403] & b[379])^(a[402] & b[380])^(a[401] & b[381])^(a[400] & b[382])^(a[399] & b[383])^(a[398] & b[384])^(a[397] & b[385])^(a[396] & b[386])^(a[395] & b[387])^(a[394] & b[388])^(a[393] & b[389])^(a[392] & b[390])^(a[391] & b[391])^(a[390] & b[392])^(a[389] & b[393])^(a[388] & b[394])^(a[387] & b[395])^(a[386] & b[396])^(a[385] & b[397])^(a[384] & b[398])^(a[383] & b[399])^(a[382] & b[400])^(a[381] & b[401])^(a[380] & b[402])^(a[379] & b[403])^(a[378] & b[404])^(a[377] & b[405])^(a[376] & b[406])^(a[375] & b[407])^(a[374] & b[408]);
assign y[783] = (a[408] & b[375])^(a[407] & b[376])^(a[406] & b[377])^(a[405] & b[378])^(a[404] & b[379])^(a[403] & b[380])^(a[402] & b[381])^(a[401] & b[382])^(a[400] & b[383])^(a[399] & b[384])^(a[398] & b[385])^(a[397] & b[386])^(a[396] & b[387])^(a[395] & b[388])^(a[394] & b[389])^(a[393] & b[390])^(a[392] & b[391])^(a[391] & b[392])^(a[390] & b[393])^(a[389] & b[394])^(a[388] & b[395])^(a[387] & b[396])^(a[386] & b[397])^(a[385] & b[398])^(a[384] & b[399])^(a[383] & b[400])^(a[382] & b[401])^(a[381] & b[402])^(a[380] & b[403])^(a[379] & b[404])^(a[378] & b[405])^(a[377] & b[406])^(a[376] & b[407])^(a[375] & b[408]);
assign y[784] = (a[408] & b[376])^(a[407] & b[377])^(a[406] & b[378])^(a[405] & b[379])^(a[404] & b[380])^(a[403] & b[381])^(a[402] & b[382])^(a[401] & b[383])^(a[400] & b[384])^(a[399] & b[385])^(a[398] & b[386])^(a[397] & b[387])^(a[396] & b[388])^(a[395] & b[389])^(a[394] & b[390])^(a[393] & b[391])^(a[392] & b[392])^(a[391] & b[393])^(a[390] & b[394])^(a[389] & b[395])^(a[388] & b[396])^(a[387] & b[397])^(a[386] & b[398])^(a[385] & b[399])^(a[384] & b[400])^(a[383] & b[401])^(a[382] & b[402])^(a[381] & b[403])^(a[380] & b[404])^(a[379] & b[405])^(a[378] & b[406])^(a[377] & b[407])^(a[376] & b[408]);
assign y[785] = (a[408] & b[377])^(a[407] & b[378])^(a[406] & b[379])^(a[405] & b[380])^(a[404] & b[381])^(a[403] & b[382])^(a[402] & b[383])^(a[401] & b[384])^(a[400] & b[385])^(a[399] & b[386])^(a[398] & b[387])^(a[397] & b[388])^(a[396] & b[389])^(a[395] & b[390])^(a[394] & b[391])^(a[393] & b[392])^(a[392] & b[393])^(a[391] & b[394])^(a[390] & b[395])^(a[389] & b[396])^(a[388] & b[397])^(a[387] & b[398])^(a[386] & b[399])^(a[385] & b[400])^(a[384] & b[401])^(a[383] & b[402])^(a[382] & b[403])^(a[381] & b[404])^(a[380] & b[405])^(a[379] & b[406])^(a[378] & b[407])^(a[377] & b[408]);
assign y[786] = (a[408] & b[378])^(a[407] & b[379])^(a[406] & b[380])^(a[405] & b[381])^(a[404] & b[382])^(a[403] & b[383])^(a[402] & b[384])^(a[401] & b[385])^(a[400] & b[386])^(a[399] & b[387])^(a[398] & b[388])^(a[397] & b[389])^(a[396] & b[390])^(a[395] & b[391])^(a[394] & b[392])^(a[393] & b[393])^(a[392] & b[394])^(a[391] & b[395])^(a[390] & b[396])^(a[389] & b[397])^(a[388] & b[398])^(a[387] & b[399])^(a[386] & b[400])^(a[385] & b[401])^(a[384] & b[402])^(a[383] & b[403])^(a[382] & b[404])^(a[381] & b[405])^(a[380] & b[406])^(a[379] & b[407])^(a[378] & b[408]);
assign y[787] = (a[408] & b[379])^(a[407] & b[380])^(a[406] & b[381])^(a[405] & b[382])^(a[404] & b[383])^(a[403] & b[384])^(a[402] & b[385])^(a[401] & b[386])^(a[400] & b[387])^(a[399] & b[388])^(a[398] & b[389])^(a[397] & b[390])^(a[396] & b[391])^(a[395] & b[392])^(a[394] & b[393])^(a[393] & b[394])^(a[392] & b[395])^(a[391] & b[396])^(a[390] & b[397])^(a[389] & b[398])^(a[388] & b[399])^(a[387] & b[400])^(a[386] & b[401])^(a[385] & b[402])^(a[384] & b[403])^(a[383] & b[404])^(a[382] & b[405])^(a[381] & b[406])^(a[380] & b[407])^(a[379] & b[408]);
assign y[788] = (a[408] & b[380])^(a[407] & b[381])^(a[406] & b[382])^(a[405] & b[383])^(a[404] & b[384])^(a[403] & b[385])^(a[402] & b[386])^(a[401] & b[387])^(a[400] & b[388])^(a[399] & b[389])^(a[398] & b[390])^(a[397] & b[391])^(a[396] & b[392])^(a[395] & b[393])^(a[394] & b[394])^(a[393] & b[395])^(a[392] & b[396])^(a[391] & b[397])^(a[390] & b[398])^(a[389] & b[399])^(a[388] & b[400])^(a[387] & b[401])^(a[386] & b[402])^(a[385] & b[403])^(a[384] & b[404])^(a[383] & b[405])^(a[382] & b[406])^(a[381] & b[407])^(a[380] & b[408]);
assign y[789] = (a[408] & b[381])^(a[407] & b[382])^(a[406] & b[383])^(a[405] & b[384])^(a[404] & b[385])^(a[403] & b[386])^(a[402] & b[387])^(a[401] & b[388])^(a[400] & b[389])^(a[399] & b[390])^(a[398] & b[391])^(a[397] & b[392])^(a[396] & b[393])^(a[395] & b[394])^(a[394] & b[395])^(a[393] & b[396])^(a[392] & b[397])^(a[391] & b[398])^(a[390] & b[399])^(a[389] & b[400])^(a[388] & b[401])^(a[387] & b[402])^(a[386] & b[403])^(a[385] & b[404])^(a[384] & b[405])^(a[383] & b[406])^(a[382] & b[407])^(a[381] & b[408]);
assign y[790] = (a[408] & b[382])^(a[407] & b[383])^(a[406] & b[384])^(a[405] & b[385])^(a[404] & b[386])^(a[403] & b[387])^(a[402] & b[388])^(a[401] & b[389])^(a[400] & b[390])^(a[399] & b[391])^(a[398] & b[392])^(a[397] & b[393])^(a[396] & b[394])^(a[395] & b[395])^(a[394] & b[396])^(a[393] & b[397])^(a[392] & b[398])^(a[391] & b[399])^(a[390] & b[400])^(a[389] & b[401])^(a[388] & b[402])^(a[387] & b[403])^(a[386] & b[404])^(a[385] & b[405])^(a[384] & b[406])^(a[383] & b[407])^(a[382] & b[408]);
assign y[791] = (a[408] & b[383])^(a[407] & b[384])^(a[406] & b[385])^(a[405] & b[386])^(a[404] & b[387])^(a[403] & b[388])^(a[402] & b[389])^(a[401] & b[390])^(a[400] & b[391])^(a[399] & b[392])^(a[398] & b[393])^(a[397] & b[394])^(a[396] & b[395])^(a[395] & b[396])^(a[394] & b[397])^(a[393] & b[398])^(a[392] & b[399])^(a[391] & b[400])^(a[390] & b[401])^(a[389] & b[402])^(a[388] & b[403])^(a[387] & b[404])^(a[386] & b[405])^(a[385] & b[406])^(a[384] & b[407])^(a[383] & b[408]);
assign y[792] = (a[408] & b[384])^(a[407] & b[385])^(a[406] & b[386])^(a[405] & b[387])^(a[404] & b[388])^(a[403] & b[389])^(a[402] & b[390])^(a[401] & b[391])^(a[400] & b[392])^(a[399] & b[393])^(a[398] & b[394])^(a[397] & b[395])^(a[396] & b[396])^(a[395] & b[397])^(a[394] & b[398])^(a[393] & b[399])^(a[392] & b[400])^(a[391] & b[401])^(a[390] & b[402])^(a[389] & b[403])^(a[388] & b[404])^(a[387] & b[405])^(a[386] & b[406])^(a[385] & b[407])^(a[384] & b[408]);
assign y[793] = (a[408] & b[385])^(a[407] & b[386])^(a[406] & b[387])^(a[405] & b[388])^(a[404] & b[389])^(a[403] & b[390])^(a[402] & b[391])^(a[401] & b[392])^(a[400] & b[393])^(a[399] & b[394])^(a[398] & b[395])^(a[397] & b[396])^(a[396] & b[397])^(a[395] & b[398])^(a[394] & b[399])^(a[393] & b[400])^(a[392] & b[401])^(a[391] & b[402])^(a[390] & b[403])^(a[389] & b[404])^(a[388] & b[405])^(a[387] & b[406])^(a[386] & b[407])^(a[385] & b[408]);
assign y[794] = (a[408] & b[386])^(a[407] & b[387])^(a[406] & b[388])^(a[405] & b[389])^(a[404] & b[390])^(a[403] & b[391])^(a[402] & b[392])^(a[401] & b[393])^(a[400] & b[394])^(a[399] & b[395])^(a[398] & b[396])^(a[397] & b[397])^(a[396] & b[398])^(a[395] & b[399])^(a[394] & b[400])^(a[393] & b[401])^(a[392] & b[402])^(a[391] & b[403])^(a[390] & b[404])^(a[389] & b[405])^(a[388] & b[406])^(a[387] & b[407])^(a[386] & b[408]);
assign y[795] = (a[408] & b[387])^(a[407] & b[388])^(a[406] & b[389])^(a[405] & b[390])^(a[404] & b[391])^(a[403] & b[392])^(a[402] & b[393])^(a[401] & b[394])^(a[400] & b[395])^(a[399] & b[396])^(a[398] & b[397])^(a[397] & b[398])^(a[396] & b[399])^(a[395] & b[400])^(a[394] & b[401])^(a[393] & b[402])^(a[392] & b[403])^(a[391] & b[404])^(a[390] & b[405])^(a[389] & b[406])^(a[388] & b[407])^(a[387] & b[408]);
assign y[796] = (a[408] & b[388])^(a[407] & b[389])^(a[406] & b[390])^(a[405] & b[391])^(a[404] & b[392])^(a[403] & b[393])^(a[402] & b[394])^(a[401] & b[395])^(a[400] & b[396])^(a[399] & b[397])^(a[398] & b[398])^(a[397] & b[399])^(a[396] & b[400])^(a[395] & b[401])^(a[394] & b[402])^(a[393] & b[403])^(a[392] & b[404])^(a[391] & b[405])^(a[390] & b[406])^(a[389] & b[407])^(a[388] & b[408]);
assign y[797] = (a[408] & b[389])^(a[407] & b[390])^(a[406] & b[391])^(a[405] & b[392])^(a[404] & b[393])^(a[403] & b[394])^(a[402] & b[395])^(a[401] & b[396])^(a[400] & b[397])^(a[399] & b[398])^(a[398] & b[399])^(a[397] & b[400])^(a[396] & b[401])^(a[395] & b[402])^(a[394] & b[403])^(a[393] & b[404])^(a[392] & b[405])^(a[391] & b[406])^(a[390] & b[407])^(a[389] & b[408]);
assign y[798] = (a[408] & b[390])^(a[407] & b[391])^(a[406] & b[392])^(a[405] & b[393])^(a[404] & b[394])^(a[403] & b[395])^(a[402] & b[396])^(a[401] & b[397])^(a[400] & b[398])^(a[399] & b[399])^(a[398] & b[400])^(a[397] & b[401])^(a[396] & b[402])^(a[395] & b[403])^(a[394] & b[404])^(a[393] & b[405])^(a[392] & b[406])^(a[391] & b[407])^(a[390] & b[408]);
assign y[799] = (a[408] & b[391])^(a[407] & b[392])^(a[406] & b[393])^(a[405] & b[394])^(a[404] & b[395])^(a[403] & b[396])^(a[402] & b[397])^(a[401] & b[398])^(a[400] & b[399])^(a[399] & b[400])^(a[398] & b[401])^(a[397] & b[402])^(a[396] & b[403])^(a[395] & b[404])^(a[394] & b[405])^(a[393] & b[406])^(a[392] & b[407])^(a[391] & b[408]);
assign y[800] = (a[408] & b[392])^(a[407] & b[393])^(a[406] & b[394])^(a[405] & b[395])^(a[404] & b[396])^(a[403] & b[397])^(a[402] & b[398])^(a[401] & b[399])^(a[400] & b[400])^(a[399] & b[401])^(a[398] & b[402])^(a[397] & b[403])^(a[396] & b[404])^(a[395] & b[405])^(a[394] & b[406])^(a[393] & b[407])^(a[392] & b[408]);
assign y[801] = (a[408] & b[393])^(a[407] & b[394])^(a[406] & b[395])^(a[405] & b[396])^(a[404] & b[397])^(a[403] & b[398])^(a[402] & b[399])^(a[401] & b[400])^(a[400] & b[401])^(a[399] & b[402])^(a[398] & b[403])^(a[397] & b[404])^(a[396] & b[405])^(a[395] & b[406])^(a[394] & b[407])^(a[393] & b[408]);
assign y[802] = (a[408] & b[394])^(a[407] & b[395])^(a[406] & b[396])^(a[405] & b[397])^(a[404] & b[398])^(a[403] & b[399])^(a[402] & b[400])^(a[401] & b[401])^(a[400] & b[402])^(a[399] & b[403])^(a[398] & b[404])^(a[397] & b[405])^(a[396] & b[406])^(a[395] & b[407])^(a[394] & b[408]);
assign y[803] = (a[408] & b[395])^(a[407] & b[396])^(a[406] & b[397])^(a[405] & b[398])^(a[404] & b[399])^(a[403] & b[400])^(a[402] & b[401])^(a[401] & b[402])^(a[400] & b[403])^(a[399] & b[404])^(a[398] & b[405])^(a[397] & b[406])^(a[396] & b[407])^(a[395] & b[408]);
assign y[804] = (a[408] & b[396])^(a[407] & b[397])^(a[406] & b[398])^(a[405] & b[399])^(a[404] & b[400])^(a[403] & b[401])^(a[402] & b[402])^(a[401] & b[403])^(a[400] & b[404])^(a[399] & b[405])^(a[398] & b[406])^(a[397] & b[407])^(a[396] & b[408]);
assign y[805] = (a[408] & b[397])^(a[407] & b[398])^(a[406] & b[399])^(a[405] & b[400])^(a[404] & b[401])^(a[403] & b[402])^(a[402] & b[403])^(a[401] & b[404])^(a[400] & b[405])^(a[399] & b[406])^(a[398] & b[407])^(a[397] & b[408]);
assign y[806] = (a[408] & b[398])^(a[407] & b[399])^(a[406] & b[400])^(a[405] & b[401])^(a[404] & b[402])^(a[403] & b[403])^(a[402] & b[404])^(a[401] & b[405])^(a[400] & b[406])^(a[399] & b[407])^(a[398] & b[408]);
assign y[807] = (a[408] & b[399])^(a[407] & b[400])^(a[406] & b[401])^(a[405] & b[402])^(a[404] & b[403])^(a[403] & b[404])^(a[402] & b[405])^(a[401] & b[406])^(a[400] & b[407])^(a[399] & b[408]);
assign y[808] = (a[408] & b[400])^(a[407] & b[401])^(a[406] & b[402])^(a[405] & b[403])^(a[404] & b[404])^(a[403] & b[405])^(a[402] & b[406])^(a[401] & b[407])^(a[400] & b[408]);
assign y[809] = (a[408] & b[401])^(a[407] & b[402])^(a[406] & b[403])^(a[405] & b[404])^(a[404] & b[405])^(a[403] & b[406])^(a[402] & b[407])^(a[401] & b[408]);
assign y[810] = (a[408] & b[402])^(a[407] & b[403])^(a[406] & b[404])^(a[405] & b[405])^(a[404] & b[406])^(a[403] & b[407])^(a[402] & b[408]);
assign y[811] = (a[408] & b[403])^(a[407] & b[404])^(a[406] & b[405])^(a[405] & b[406])^(a[404] & b[407])^(a[403] & b[408]);
assign y[812] = (a[408] & b[404])^(a[407] & b[405])^(a[406] & b[406])^(a[405] & b[407])^(a[404] & b[408]);
assign y[813] = (a[408] & b[405])^(a[407] & b[406])^(a[406] & b[407])^(a[405] & b[408]);
assign y[814] = (a[408] & b[406])^(a[407] & b[407])^(a[406] & b[408]);
assign y[815] = (a[408] & b[407])^(a[407] & b[408]);
assign y[816] = (a[408] & b[408]);


endmodule
