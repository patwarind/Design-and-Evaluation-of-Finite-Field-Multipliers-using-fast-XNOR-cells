`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Nitin D. Patwari
// 
// Create Date: 20.01.2022 22:17:47
// Design Name: 
// Module Name: CA_163bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CA_163bit(
    a,
    b,
    y
    );

input [162:0] a;
input [162:0] b;

output [324:0] y;


assign y[0] = (a[0] & b[0]);
assign y[1] = (a[1] & b[0])^(a[0] & b[1]);
assign y[2] = (a[2] & b[0])^(a[1] & b[1])^(a[0] & b[2]);
assign y[3] = (a[3] & b[0])^(a[2] & b[1])^(a[1] & b[2])^(a[0] & b[3]);
assign y[4] = (a[4] & b[0])^(a[3] & b[1])^(a[2] & b[2])^(a[1] & b[3])^(a[0] & b[4]);
assign y[5] = (a[5] & b[0])^(a[4] & b[1])^(a[3] & b[2])^(a[2] & b[3])^(a[1] & b[4])^(a[0] & b[5]);
assign y[6] = (a[6] & b[0])^(a[5] & b[1])^(a[4] & b[2])^(a[3] & b[3])^(a[2] & b[4])^(a[1] & b[5])^(a[0] & b[6]);
assign y[7] = (a[7] & b[0])^(a[6] & b[1])^(a[5] & b[2])^(a[4] & b[3])^(a[3] & b[4])^(a[2] & b[5])^(a[1] & b[6])^(a[0] & b[7]);
assign y[8] = (a[8] & b[0])^(a[7] & b[1])^(a[6] & b[2])^(a[5] & b[3])^(a[4] & b[4])^(a[3] & b[5])^(a[2] & b[6])^(a[1] & b[7])^(a[0] & b[8]);
assign y[9] = (a[9] & b[0])^(a[8] & b[1])^(a[7] & b[2])^(a[6] & b[3])^(a[5] & b[4])^(a[4] & b[5])^(a[3] & b[6])^(a[2] & b[7])^(a[1] & b[8])^(a[0] & b[9]);
assign y[10] = (a[10] & b[0])^(a[9] & b[1])^(a[8] & b[2])^(a[7] & b[3])^(a[6] & b[4])^(a[5] & b[5])^(a[4] & b[6])^(a[3] & b[7])^(a[2] & b[8])^(a[1] & b[9])^(a[0] & b[10]);
assign y[11] = (a[11] & b[0])^(a[10] & b[1])^(a[9] & b[2])^(a[8] & b[3])^(a[7] & b[4])^(a[6] & b[5])^(a[5] & b[6])^(a[4] & b[7])^(a[3] & b[8])^(a[2] & b[9])^(a[1] & b[10])^(a[0] & b[11]);
assign y[12] = (a[12] & b[0])^(a[11] & b[1])^(a[10] & b[2])^(a[9] & b[3])^(a[8] & b[4])^(a[7] & b[5])^(a[6] & b[6])^(a[5] & b[7])^(a[4] & b[8])^(a[3] & b[9])^(a[2] & b[10])^(a[1] & b[11])^(a[0] & b[12]);
assign y[13] = (a[13] & b[0])^(a[12] & b[1])^(a[11] & b[2])^(a[10] & b[3])^(a[9] & b[4])^(a[8] & b[5])^(a[7] & b[6])^(a[6] & b[7])^(a[5] & b[8])^(a[4] & b[9])^(a[3] & b[10])^(a[2] & b[11])^(a[1] & b[12])^(a[0] & b[13]);
assign y[14] = (a[14] & b[0])^(a[13] & b[1])^(a[12] & b[2])^(a[11] & b[3])^(a[10] & b[4])^(a[9] & b[5])^(a[8] & b[6])^(a[7] & b[7])^(a[6] & b[8])^(a[5] & b[9])^(a[4] & b[10])^(a[3] & b[11])^(a[2] & b[12])^(a[1] & b[13])^(a[0] & b[14]);
assign y[15] = (a[15] & b[0])^(a[14] & b[1])^(a[13] & b[2])^(a[12] & b[3])^(a[11] & b[4])^(a[10] & b[5])^(a[9] & b[6])^(a[8] & b[7])^(a[7] & b[8])^(a[6] & b[9])^(a[5] & b[10])^(a[4] & b[11])^(a[3] & b[12])^(a[2] & b[13])^(a[1] & b[14])^(a[0] & b[15]);
assign y[16] = (a[16] & b[0])^(a[15] & b[1])^(a[14] & b[2])^(a[13] & b[3])^(a[12] & b[4])^(a[11] & b[5])^(a[10] & b[6])^(a[9] & b[7])^(a[8] & b[8])^(a[7] & b[9])^(a[6] & b[10])^(a[5] & b[11])^(a[4] & b[12])^(a[3] & b[13])^(a[2] & b[14])^(a[1] & b[15])^(a[0] & b[16]);
assign y[17] = (a[17] & b[0])^(a[16] & b[1])^(a[15] & b[2])^(a[14] & b[3])^(a[13] & b[4])^(a[12] & b[5])^(a[11] & b[6])^(a[10] & b[7])^(a[9] & b[8])^(a[8] & b[9])^(a[7] & b[10])^(a[6] & b[11])^(a[5] & b[12])^(a[4] & b[13])^(a[3] & b[14])^(a[2] & b[15])^(a[1] & b[16])^(a[0] & b[17]);
assign y[18] = (a[18] & b[0])^(a[17] & b[1])^(a[16] & b[2])^(a[15] & b[3])^(a[14] & b[4])^(a[13] & b[5])^(a[12] & b[6])^(a[11] & b[7])^(a[10] & b[8])^(a[9] & b[9])^(a[8] & b[10])^(a[7] & b[11])^(a[6] & b[12])^(a[5] & b[13])^(a[4] & b[14])^(a[3] & b[15])^(a[2] & b[16])^(a[1] & b[17])^(a[0] & b[18]);
assign y[19] = (a[19] & b[0])^(a[18] & b[1])^(a[17] & b[2])^(a[16] & b[3])^(a[15] & b[4])^(a[14] & b[5])^(a[13] & b[6])^(a[12] & b[7])^(a[11] & b[8])^(a[10] & b[9])^(a[9] & b[10])^(a[8] & b[11])^(a[7] & b[12])^(a[6] & b[13])^(a[5] & b[14])^(a[4] & b[15])^(a[3] & b[16])^(a[2] & b[17])^(a[1] & b[18])^(a[0] & b[19]);
assign y[20] = (a[20] & b[0])^(a[19] & b[1])^(a[18] & b[2])^(a[17] & b[3])^(a[16] & b[4])^(a[15] & b[5])^(a[14] & b[6])^(a[13] & b[7])^(a[12] & b[8])^(a[11] & b[9])^(a[10] & b[10])^(a[9] & b[11])^(a[8] & b[12])^(a[7] & b[13])^(a[6] & b[14])^(a[5] & b[15])^(a[4] & b[16])^(a[3] & b[17])^(a[2] & b[18])^(a[1] & b[19])^(a[0] & b[20]);
assign y[21] = (a[21] & b[0])^(a[20] & b[1])^(a[19] & b[2])^(a[18] & b[3])^(a[17] & b[4])^(a[16] & b[5])^(a[15] & b[6])^(a[14] & b[7])^(a[13] & b[8])^(a[12] & b[9])^(a[11] & b[10])^(a[10] & b[11])^(a[9] & b[12])^(a[8] & b[13])^(a[7] & b[14])^(a[6] & b[15])^(a[5] & b[16])^(a[4] & b[17])^(a[3] & b[18])^(a[2] & b[19])^(a[1] & b[20])^(a[0] & b[21]);
assign y[22] = (a[22] & b[0])^(a[21] & b[1])^(a[20] & b[2])^(a[19] & b[3])^(a[18] & b[4])^(a[17] & b[5])^(a[16] & b[6])^(a[15] & b[7])^(a[14] & b[8])^(a[13] & b[9])^(a[12] & b[10])^(a[11] & b[11])^(a[10] & b[12])^(a[9] & b[13])^(a[8] & b[14])^(a[7] & b[15])^(a[6] & b[16])^(a[5] & b[17])^(a[4] & b[18])^(a[3] & b[19])^(a[2] & b[20])^(a[1] & b[21])^(a[0] & b[22]);
assign y[23] = (a[23] & b[0])^(a[22] & b[1])^(a[21] & b[2])^(a[20] & b[3])^(a[19] & b[4])^(a[18] & b[5])^(a[17] & b[6])^(a[16] & b[7])^(a[15] & b[8])^(a[14] & b[9])^(a[13] & b[10])^(a[12] & b[11])^(a[11] & b[12])^(a[10] & b[13])^(a[9] & b[14])^(a[8] & b[15])^(a[7] & b[16])^(a[6] & b[17])^(a[5] & b[18])^(a[4] & b[19])^(a[3] & b[20])^(a[2] & b[21])^(a[1] & b[22])^(a[0] & b[23]);
assign y[24] = (a[24] & b[0])^(a[23] & b[1])^(a[22] & b[2])^(a[21] & b[3])^(a[20] & b[4])^(a[19] & b[5])^(a[18] & b[6])^(a[17] & b[7])^(a[16] & b[8])^(a[15] & b[9])^(a[14] & b[10])^(a[13] & b[11])^(a[12] & b[12])^(a[11] & b[13])^(a[10] & b[14])^(a[9] & b[15])^(a[8] & b[16])^(a[7] & b[17])^(a[6] & b[18])^(a[5] & b[19])^(a[4] & b[20])^(a[3] & b[21])^(a[2] & b[22])^(a[1] & b[23])^(a[0] & b[24]);
assign y[25] = (a[25] & b[0])^(a[24] & b[1])^(a[23] & b[2])^(a[22] & b[3])^(a[21] & b[4])^(a[20] & b[5])^(a[19] & b[6])^(a[18] & b[7])^(a[17] & b[8])^(a[16] & b[9])^(a[15] & b[10])^(a[14] & b[11])^(a[13] & b[12])^(a[12] & b[13])^(a[11] & b[14])^(a[10] & b[15])^(a[9] & b[16])^(a[8] & b[17])^(a[7] & b[18])^(a[6] & b[19])^(a[5] & b[20])^(a[4] & b[21])^(a[3] & b[22])^(a[2] & b[23])^(a[1] & b[24])^(a[0] & b[25]);
assign y[26] = (a[26] & b[0])^(a[25] & b[1])^(a[24] & b[2])^(a[23] & b[3])^(a[22] & b[4])^(a[21] & b[5])^(a[20] & b[6])^(a[19] & b[7])^(a[18] & b[8])^(a[17] & b[9])^(a[16] & b[10])^(a[15] & b[11])^(a[14] & b[12])^(a[13] & b[13])^(a[12] & b[14])^(a[11] & b[15])^(a[10] & b[16])^(a[9] & b[17])^(a[8] & b[18])^(a[7] & b[19])^(a[6] & b[20])^(a[5] & b[21])^(a[4] & b[22])^(a[3] & b[23])^(a[2] & b[24])^(a[1] & b[25])^(a[0] & b[26]);
assign y[27] = (a[27] & b[0])^(a[26] & b[1])^(a[25] & b[2])^(a[24] & b[3])^(a[23] & b[4])^(a[22] & b[5])^(a[21] & b[6])^(a[20] & b[7])^(a[19] & b[8])^(a[18] & b[9])^(a[17] & b[10])^(a[16] & b[11])^(a[15] & b[12])^(a[14] & b[13])^(a[13] & b[14])^(a[12] & b[15])^(a[11] & b[16])^(a[10] & b[17])^(a[9] & b[18])^(a[8] & b[19])^(a[7] & b[20])^(a[6] & b[21])^(a[5] & b[22])^(a[4] & b[23])^(a[3] & b[24])^(a[2] & b[25])^(a[1] & b[26])^(a[0] & b[27]);
assign y[28] = (a[28] & b[0])^(a[27] & b[1])^(a[26] & b[2])^(a[25] & b[3])^(a[24] & b[4])^(a[23] & b[5])^(a[22] & b[6])^(a[21] & b[7])^(a[20] & b[8])^(a[19] & b[9])^(a[18] & b[10])^(a[17] & b[11])^(a[16] & b[12])^(a[15] & b[13])^(a[14] & b[14])^(a[13] & b[15])^(a[12] & b[16])^(a[11] & b[17])^(a[10] & b[18])^(a[9] & b[19])^(a[8] & b[20])^(a[7] & b[21])^(a[6] & b[22])^(a[5] & b[23])^(a[4] & b[24])^(a[3] & b[25])^(a[2] & b[26])^(a[1] & b[27])^(a[0] & b[28]);
assign y[29] = (a[29] & b[0])^(a[28] & b[1])^(a[27] & b[2])^(a[26] & b[3])^(a[25] & b[4])^(a[24] & b[5])^(a[23] & b[6])^(a[22] & b[7])^(a[21] & b[8])^(a[20] & b[9])^(a[19] & b[10])^(a[18] & b[11])^(a[17] & b[12])^(a[16] & b[13])^(a[15] & b[14])^(a[14] & b[15])^(a[13] & b[16])^(a[12] & b[17])^(a[11] & b[18])^(a[10] & b[19])^(a[9] & b[20])^(a[8] & b[21])^(a[7] & b[22])^(a[6] & b[23])^(a[5] & b[24])^(a[4] & b[25])^(a[3] & b[26])^(a[2] & b[27])^(a[1] & b[28])^(a[0] & b[29]);
assign y[30] = (a[30] & b[0])^(a[29] & b[1])^(a[28] & b[2])^(a[27] & b[3])^(a[26] & b[4])^(a[25] & b[5])^(a[24] & b[6])^(a[23] & b[7])^(a[22] & b[8])^(a[21] & b[9])^(a[20] & b[10])^(a[19] & b[11])^(a[18] & b[12])^(a[17] & b[13])^(a[16] & b[14])^(a[15] & b[15])^(a[14] & b[16])^(a[13] & b[17])^(a[12] & b[18])^(a[11] & b[19])^(a[10] & b[20])^(a[9] & b[21])^(a[8] & b[22])^(a[7] & b[23])^(a[6] & b[24])^(a[5] & b[25])^(a[4] & b[26])^(a[3] & b[27])^(a[2] & b[28])^(a[1] & b[29])^(a[0] & b[30]);
assign y[31] = (a[31] & b[0])^(a[30] & b[1])^(a[29] & b[2])^(a[28] & b[3])^(a[27] & b[4])^(a[26] & b[5])^(a[25] & b[6])^(a[24] & b[7])^(a[23] & b[8])^(a[22] & b[9])^(a[21] & b[10])^(a[20] & b[11])^(a[19] & b[12])^(a[18] & b[13])^(a[17] & b[14])^(a[16] & b[15])^(a[15] & b[16])^(a[14] & b[17])^(a[13] & b[18])^(a[12] & b[19])^(a[11] & b[20])^(a[10] & b[21])^(a[9] & b[22])^(a[8] & b[23])^(a[7] & b[24])^(a[6] & b[25])^(a[5] & b[26])^(a[4] & b[27])^(a[3] & b[28])^(a[2] & b[29])^(a[1] & b[30])^(a[0] & b[31]);
assign y[32] = (a[32] & b[0])^(a[31] & b[1])^(a[30] & b[2])^(a[29] & b[3])^(a[28] & b[4])^(a[27] & b[5])^(a[26] & b[6])^(a[25] & b[7])^(a[24] & b[8])^(a[23] & b[9])^(a[22] & b[10])^(a[21] & b[11])^(a[20] & b[12])^(a[19] & b[13])^(a[18] & b[14])^(a[17] & b[15])^(a[16] & b[16])^(a[15] & b[17])^(a[14] & b[18])^(a[13] & b[19])^(a[12] & b[20])^(a[11] & b[21])^(a[10] & b[22])^(a[9] & b[23])^(a[8] & b[24])^(a[7] & b[25])^(a[6] & b[26])^(a[5] & b[27])^(a[4] & b[28])^(a[3] & b[29])^(a[2] & b[30])^(a[1] & b[31])^(a[0] & b[32]);
assign y[33] = (a[33] & b[0])^(a[32] & b[1])^(a[31] & b[2])^(a[30] & b[3])^(a[29] & b[4])^(a[28] & b[5])^(a[27] & b[6])^(a[26] & b[7])^(a[25] & b[8])^(a[24] & b[9])^(a[23] & b[10])^(a[22] & b[11])^(a[21] & b[12])^(a[20] & b[13])^(a[19] & b[14])^(a[18] & b[15])^(a[17] & b[16])^(a[16] & b[17])^(a[15] & b[18])^(a[14] & b[19])^(a[13] & b[20])^(a[12] & b[21])^(a[11] & b[22])^(a[10] & b[23])^(a[9] & b[24])^(a[8] & b[25])^(a[7] & b[26])^(a[6] & b[27])^(a[5] & b[28])^(a[4] & b[29])^(a[3] & b[30])^(a[2] & b[31])^(a[1] & b[32])^(a[0] & b[33]);
assign y[34] = (a[34] & b[0])^(a[33] & b[1])^(a[32] & b[2])^(a[31] & b[3])^(a[30] & b[4])^(a[29] & b[5])^(a[28] & b[6])^(a[27] & b[7])^(a[26] & b[8])^(a[25] & b[9])^(a[24] & b[10])^(a[23] & b[11])^(a[22] & b[12])^(a[21] & b[13])^(a[20] & b[14])^(a[19] & b[15])^(a[18] & b[16])^(a[17] & b[17])^(a[16] & b[18])^(a[15] & b[19])^(a[14] & b[20])^(a[13] & b[21])^(a[12] & b[22])^(a[11] & b[23])^(a[10] & b[24])^(a[9] & b[25])^(a[8] & b[26])^(a[7] & b[27])^(a[6] & b[28])^(a[5] & b[29])^(a[4] & b[30])^(a[3] & b[31])^(a[2] & b[32])^(a[1] & b[33])^(a[0] & b[34]);
assign y[35] = (a[35] & b[0])^(a[34] & b[1])^(a[33] & b[2])^(a[32] & b[3])^(a[31] & b[4])^(a[30] & b[5])^(a[29] & b[6])^(a[28] & b[7])^(a[27] & b[8])^(a[26] & b[9])^(a[25] & b[10])^(a[24] & b[11])^(a[23] & b[12])^(a[22] & b[13])^(a[21] & b[14])^(a[20] & b[15])^(a[19] & b[16])^(a[18] & b[17])^(a[17] & b[18])^(a[16] & b[19])^(a[15] & b[20])^(a[14] & b[21])^(a[13] & b[22])^(a[12] & b[23])^(a[11] & b[24])^(a[10] & b[25])^(a[9] & b[26])^(a[8] & b[27])^(a[7] & b[28])^(a[6] & b[29])^(a[5] & b[30])^(a[4] & b[31])^(a[3] & b[32])^(a[2] & b[33])^(a[1] & b[34])^(a[0] & b[35]);
assign y[36] = (a[36] & b[0])^(a[35] & b[1])^(a[34] & b[2])^(a[33] & b[3])^(a[32] & b[4])^(a[31] & b[5])^(a[30] & b[6])^(a[29] & b[7])^(a[28] & b[8])^(a[27] & b[9])^(a[26] & b[10])^(a[25] & b[11])^(a[24] & b[12])^(a[23] & b[13])^(a[22] & b[14])^(a[21] & b[15])^(a[20] & b[16])^(a[19] & b[17])^(a[18] & b[18])^(a[17] & b[19])^(a[16] & b[20])^(a[15] & b[21])^(a[14] & b[22])^(a[13] & b[23])^(a[12] & b[24])^(a[11] & b[25])^(a[10] & b[26])^(a[9] & b[27])^(a[8] & b[28])^(a[7] & b[29])^(a[6] & b[30])^(a[5] & b[31])^(a[4] & b[32])^(a[3] & b[33])^(a[2] & b[34])^(a[1] & b[35])^(a[0] & b[36]);
assign y[37] = (a[37] & b[0])^(a[36] & b[1])^(a[35] & b[2])^(a[34] & b[3])^(a[33] & b[4])^(a[32] & b[5])^(a[31] & b[6])^(a[30] & b[7])^(a[29] & b[8])^(a[28] & b[9])^(a[27] & b[10])^(a[26] & b[11])^(a[25] & b[12])^(a[24] & b[13])^(a[23] & b[14])^(a[22] & b[15])^(a[21] & b[16])^(a[20] & b[17])^(a[19] & b[18])^(a[18] & b[19])^(a[17] & b[20])^(a[16] & b[21])^(a[15] & b[22])^(a[14] & b[23])^(a[13] & b[24])^(a[12] & b[25])^(a[11] & b[26])^(a[10] & b[27])^(a[9] & b[28])^(a[8] & b[29])^(a[7] & b[30])^(a[6] & b[31])^(a[5] & b[32])^(a[4] & b[33])^(a[3] & b[34])^(a[2] & b[35])^(a[1] & b[36])^(a[0] & b[37]);
assign y[38] = (a[38] & b[0])^(a[37] & b[1])^(a[36] & b[2])^(a[35] & b[3])^(a[34] & b[4])^(a[33] & b[5])^(a[32] & b[6])^(a[31] & b[7])^(a[30] & b[8])^(a[29] & b[9])^(a[28] & b[10])^(a[27] & b[11])^(a[26] & b[12])^(a[25] & b[13])^(a[24] & b[14])^(a[23] & b[15])^(a[22] & b[16])^(a[21] & b[17])^(a[20] & b[18])^(a[19] & b[19])^(a[18] & b[20])^(a[17] & b[21])^(a[16] & b[22])^(a[15] & b[23])^(a[14] & b[24])^(a[13] & b[25])^(a[12] & b[26])^(a[11] & b[27])^(a[10] & b[28])^(a[9] & b[29])^(a[8] & b[30])^(a[7] & b[31])^(a[6] & b[32])^(a[5] & b[33])^(a[4] & b[34])^(a[3] & b[35])^(a[2] & b[36])^(a[1] & b[37])^(a[0] & b[38]);
assign y[39] = (a[39] & b[0])^(a[38] & b[1])^(a[37] & b[2])^(a[36] & b[3])^(a[35] & b[4])^(a[34] & b[5])^(a[33] & b[6])^(a[32] & b[7])^(a[31] & b[8])^(a[30] & b[9])^(a[29] & b[10])^(a[28] & b[11])^(a[27] & b[12])^(a[26] & b[13])^(a[25] & b[14])^(a[24] & b[15])^(a[23] & b[16])^(a[22] & b[17])^(a[21] & b[18])^(a[20] & b[19])^(a[19] & b[20])^(a[18] & b[21])^(a[17] & b[22])^(a[16] & b[23])^(a[15] & b[24])^(a[14] & b[25])^(a[13] & b[26])^(a[12] & b[27])^(a[11] & b[28])^(a[10] & b[29])^(a[9] & b[30])^(a[8] & b[31])^(a[7] & b[32])^(a[6] & b[33])^(a[5] & b[34])^(a[4] & b[35])^(a[3] & b[36])^(a[2] & b[37])^(a[1] & b[38])^(a[0] & b[39]);
assign y[40] = (a[40] & b[0])^(a[39] & b[1])^(a[38] & b[2])^(a[37] & b[3])^(a[36] & b[4])^(a[35] & b[5])^(a[34] & b[6])^(a[33] & b[7])^(a[32] & b[8])^(a[31] & b[9])^(a[30] & b[10])^(a[29] & b[11])^(a[28] & b[12])^(a[27] & b[13])^(a[26] & b[14])^(a[25] & b[15])^(a[24] & b[16])^(a[23] & b[17])^(a[22] & b[18])^(a[21] & b[19])^(a[20] & b[20])^(a[19] & b[21])^(a[18] & b[22])^(a[17] & b[23])^(a[16] & b[24])^(a[15] & b[25])^(a[14] & b[26])^(a[13] & b[27])^(a[12] & b[28])^(a[11] & b[29])^(a[10] & b[30])^(a[9] & b[31])^(a[8] & b[32])^(a[7] & b[33])^(a[6] & b[34])^(a[5] & b[35])^(a[4] & b[36])^(a[3] & b[37])^(a[2] & b[38])^(a[1] & b[39])^(a[0] & b[40]);
assign y[41] = (a[41] & b[0])^(a[40] & b[1])^(a[39] & b[2])^(a[38] & b[3])^(a[37] & b[4])^(a[36] & b[5])^(a[35] & b[6])^(a[34] & b[7])^(a[33] & b[8])^(a[32] & b[9])^(a[31] & b[10])^(a[30] & b[11])^(a[29] & b[12])^(a[28] & b[13])^(a[27] & b[14])^(a[26] & b[15])^(a[25] & b[16])^(a[24] & b[17])^(a[23] & b[18])^(a[22] & b[19])^(a[21] & b[20])^(a[20] & b[21])^(a[19] & b[22])^(a[18] & b[23])^(a[17] & b[24])^(a[16] & b[25])^(a[15] & b[26])^(a[14] & b[27])^(a[13] & b[28])^(a[12] & b[29])^(a[11] & b[30])^(a[10] & b[31])^(a[9] & b[32])^(a[8] & b[33])^(a[7] & b[34])^(a[6] & b[35])^(a[5] & b[36])^(a[4] & b[37])^(a[3] & b[38])^(a[2] & b[39])^(a[1] & b[40])^(a[0] & b[41]);
assign y[42] = (a[42] & b[0])^(a[41] & b[1])^(a[40] & b[2])^(a[39] & b[3])^(a[38] & b[4])^(a[37] & b[5])^(a[36] & b[6])^(a[35] & b[7])^(a[34] & b[8])^(a[33] & b[9])^(a[32] & b[10])^(a[31] & b[11])^(a[30] & b[12])^(a[29] & b[13])^(a[28] & b[14])^(a[27] & b[15])^(a[26] & b[16])^(a[25] & b[17])^(a[24] & b[18])^(a[23] & b[19])^(a[22] & b[20])^(a[21] & b[21])^(a[20] & b[22])^(a[19] & b[23])^(a[18] & b[24])^(a[17] & b[25])^(a[16] & b[26])^(a[15] & b[27])^(a[14] & b[28])^(a[13] & b[29])^(a[12] & b[30])^(a[11] & b[31])^(a[10] & b[32])^(a[9] & b[33])^(a[8] & b[34])^(a[7] & b[35])^(a[6] & b[36])^(a[5] & b[37])^(a[4] & b[38])^(a[3] & b[39])^(a[2] & b[40])^(a[1] & b[41])^(a[0] & b[42]);
assign y[43] = (a[43] & b[0])^(a[42] & b[1])^(a[41] & b[2])^(a[40] & b[3])^(a[39] & b[4])^(a[38] & b[5])^(a[37] & b[6])^(a[36] & b[7])^(a[35] & b[8])^(a[34] & b[9])^(a[33] & b[10])^(a[32] & b[11])^(a[31] & b[12])^(a[30] & b[13])^(a[29] & b[14])^(a[28] & b[15])^(a[27] & b[16])^(a[26] & b[17])^(a[25] & b[18])^(a[24] & b[19])^(a[23] & b[20])^(a[22] & b[21])^(a[21] & b[22])^(a[20] & b[23])^(a[19] & b[24])^(a[18] & b[25])^(a[17] & b[26])^(a[16] & b[27])^(a[15] & b[28])^(a[14] & b[29])^(a[13] & b[30])^(a[12] & b[31])^(a[11] & b[32])^(a[10] & b[33])^(a[9] & b[34])^(a[8] & b[35])^(a[7] & b[36])^(a[6] & b[37])^(a[5] & b[38])^(a[4] & b[39])^(a[3] & b[40])^(a[2] & b[41])^(a[1] & b[42])^(a[0] & b[43]);
assign y[44] = (a[44] & b[0])^(a[43] & b[1])^(a[42] & b[2])^(a[41] & b[3])^(a[40] & b[4])^(a[39] & b[5])^(a[38] & b[6])^(a[37] & b[7])^(a[36] & b[8])^(a[35] & b[9])^(a[34] & b[10])^(a[33] & b[11])^(a[32] & b[12])^(a[31] & b[13])^(a[30] & b[14])^(a[29] & b[15])^(a[28] & b[16])^(a[27] & b[17])^(a[26] & b[18])^(a[25] & b[19])^(a[24] & b[20])^(a[23] & b[21])^(a[22] & b[22])^(a[21] & b[23])^(a[20] & b[24])^(a[19] & b[25])^(a[18] & b[26])^(a[17] & b[27])^(a[16] & b[28])^(a[15] & b[29])^(a[14] & b[30])^(a[13] & b[31])^(a[12] & b[32])^(a[11] & b[33])^(a[10] & b[34])^(a[9] & b[35])^(a[8] & b[36])^(a[7] & b[37])^(a[6] & b[38])^(a[5] & b[39])^(a[4] & b[40])^(a[3] & b[41])^(a[2] & b[42])^(a[1] & b[43])^(a[0] & b[44]);
assign y[45] = (a[45] & b[0])^(a[44] & b[1])^(a[43] & b[2])^(a[42] & b[3])^(a[41] & b[4])^(a[40] & b[5])^(a[39] & b[6])^(a[38] & b[7])^(a[37] & b[8])^(a[36] & b[9])^(a[35] & b[10])^(a[34] & b[11])^(a[33] & b[12])^(a[32] & b[13])^(a[31] & b[14])^(a[30] & b[15])^(a[29] & b[16])^(a[28] & b[17])^(a[27] & b[18])^(a[26] & b[19])^(a[25] & b[20])^(a[24] & b[21])^(a[23] & b[22])^(a[22] & b[23])^(a[21] & b[24])^(a[20] & b[25])^(a[19] & b[26])^(a[18] & b[27])^(a[17] & b[28])^(a[16] & b[29])^(a[15] & b[30])^(a[14] & b[31])^(a[13] & b[32])^(a[12] & b[33])^(a[11] & b[34])^(a[10] & b[35])^(a[9] & b[36])^(a[8] & b[37])^(a[7] & b[38])^(a[6] & b[39])^(a[5] & b[40])^(a[4] & b[41])^(a[3] & b[42])^(a[2] & b[43])^(a[1] & b[44])^(a[0] & b[45]);
assign y[46] = (a[46] & b[0])^(a[45] & b[1])^(a[44] & b[2])^(a[43] & b[3])^(a[42] & b[4])^(a[41] & b[5])^(a[40] & b[6])^(a[39] & b[7])^(a[38] & b[8])^(a[37] & b[9])^(a[36] & b[10])^(a[35] & b[11])^(a[34] & b[12])^(a[33] & b[13])^(a[32] & b[14])^(a[31] & b[15])^(a[30] & b[16])^(a[29] & b[17])^(a[28] & b[18])^(a[27] & b[19])^(a[26] & b[20])^(a[25] & b[21])^(a[24] & b[22])^(a[23] & b[23])^(a[22] & b[24])^(a[21] & b[25])^(a[20] & b[26])^(a[19] & b[27])^(a[18] & b[28])^(a[17] & b[29])^(a[16] & b[30])^(a[15] & b[31])^(a[14] & b[32])^(a[13] & b[33])^(a[12] & b[34])^(a[11] & b[35])^(a[10] & b[36])^(a[9] & b[37])^(a[8] & b[38])^(a[7] & b[39])^(a[6] & b[40])^(a[5] & b[41])^(a[4] & b[42])^(a[3] & b[43])^(a[2] & b[44])^(a[1] & b[45])^(a[0] & b[46]);
assign y[47] = (a[47] & b[0])^(a[46] & b[1])^(a[45] & b[2])^(a[44] & b[3])^(a[43] & b[4])^(a[42] & b[5])^(a[41] & b[6])^(a[40] & b[7])^(a[39] & b[8])^(a[38] & b[9])^(a[37] & b[10])^(a[36] & b[11])^(a[35] & b[12])^(a[34] & b[13])^(a[33] & b[14])^(a[32] & b[15])^(a[31] & b[16])^(a[30] & b[17])^(a[29] & b[18])^(a[28] & b[19])^(a[27] & b[20])^(a[26] & b[21])^(a[25] & b[22])^(a[24] & b[23])^(a[23] & b[24])^(a[22] & b[25])^(a[21] & b[26])^(a[20] & b[27])^(a[19] & b[28])^(a[18] & b[29])^(a[17] & b[30])^(a[16] & b[31])^(a[15] & b[32])^(a[14] & b[33])^(a[13] & b[34])^(a[12] & b[35])^(a[11] & b[36])^(a[10] & b[37])^(a[9] & b[38])^(a[8] & b[39])^(a[7] & b[40])^(a[6] & b[41])^(a[5] & b[42])^(a[4] & b[43])^(a[3] & b[44])^(a[2] & b[45])^(a[1] & b[46])^(a[0] & b[47]);
assign y[48] = (a[48] & b[0])^(a[47] & b[1])^(a[46] & b[2])^(a[45] & b[3])^(a[44] & b[4])^(a[43] & b[5])^(a[42] & b[6])^(a[41] & b[7])^(a[40] & b[8])^(a[39] & b[9])^(a[38] & b[10])^(a[37] & b[11])^(a[36] & b[12])^(a[35] & b[13])^(a[34] & b[14])^(a[33] & b[15])^(a[32] & b[16])^(a[31] & b[17])^(a[30] & b[18])^(a[29] & b[19])^(a[28] & b[20])^(a[27] & b[21])^(a[26] & b[22])^(a[25] & b[23])^(a[24] & b[24])^(a[23] & b[25])^(a[22] & b[26])^(a[21] & b[27])^(a[20] & b[28])^(a[19] & b[29])^(a[18] & b[30])^(a[17] & b[31])^(a[16] & b[32])^(a[15] & b[33])^(a[14] & b[34])^(a[13] & b[35])^(a[12] & b[36])^(a[11] & b[37])^(a[10] & b[38])^(a[9] & b[39])^(a[8] & b[40])^(a[7] & b[41])^(a[6] & b[42])^(a[5] & b[43])^(a[4] & b[44])^(a[3] & b[45])^(a[2] & b[46])^(a[1] & b[47])^(a[0] & b[48]);
assign y[49] = (a[49] & b[0])^(a[48] & b[1])^(a[47] & b[2])^(a[46] & b[3])^(a[45] & b[4])^(a[44] & b[5])^(a[43] & b[6])^(a[42] & b[7])^(a[41] & b[8])^(a[40] & b[9])^(a[39] & b[10])^(a[38] & b[11])^(a[37] & b[12])^(a[36] & b[13])^(a[35] & b[14])^(a[34] & b[15])^(a[33] & b[16])^(a[32] & b[17])^(a[31] & b[18])^(a[30] & b[19])^(a[29] & b[20])^(a[28] & b[21])^(a[27] & b[22])^(a[26] & b[23])^(a[25] & b[24])^(a[24] & b[25])^(a[23] & b[26])^(a[22] & b[27])^(a[21] & b[28])^(a[20] & b[29])^(a[19] & b[30])^(a[18] & b[31])^(a[17] & b[32])^(a[16] & b[33])^(a[15] & b[34])^(a[14] & b[35])^(a[13] & b[36])^(a[12] & b[37])^(a[11] & b[38])^(a[10] & b[39])^(a[9] & b[40])^(a[8] & b[41])^(a[7] & b[42])^(a[6] & b[43])^(a[5] & b[44])^(a[4] & b[45])^(a[3] & b[46])^(a[2] & b[47])^(a[1] & b[48])^(a[0] & b[49]);
assign y[50] = (a[50] & b[0])^(a[49] & b[1])^(a[48] & b[2])^(a[47] & b[3])^(a[46] & b[4])^(a[45] & b[5])^(a[44] & b[6])^(a[43] & b[7])^(a[42] & b[8])^(a[41] & b[9])^(a[40] & b[10])^(a[39] & b[11])^(a[38] & b[12])^(a[37] & b[13])^(a[36] & b[14])^(a[35] & b[15])^(a[34] & b[16])^(a[33] & b[17])^(a[32] & b[18])^(a[31] & b[19])^(a[30] & b[20])^(a[29] & b[21])^(a[28] & b[22])^(a[27] & b[23])^(a[26] & b[24])^(a[25] & b[25])^(a[24] & b[26])^(a[23] & b[27])^(a[22] & b[28])^(a[21] & b[29])^(a[20] & b[30])^(a[19] & b[31])^(a[18] & b[32])^(a[17] & b[33])^(a[16] & b[34])^(a[15] & b[35])^(a[14] & b[36])^(a[13] & b[37])^(a[12] & b[38])^(a[11] & b[39])^(a[10] & b[40])^(a[9] & b[41])^(a[8] & b[42])^(a[7] & b[43])^(a[6] & b[44])^(a[5] & b[45])^(a[4] & b[46])^(a[3] & b[47])^(a[2] & b[48])^(a[1] & b[49])^(a[0] & b[50]);
assign y[51] = (a[51] & b[0])^(a[50] & b[1])^(a[49] & b[2])^(a[48] & b[3])^(a[47] & b[4])^(a[46] & b[5])^(a[45] & b[6])^(a[44] & b[7])^(a[43] & b[8])^(a[42] & b[9])^(a[41] & b[10])^(a[40] & b[11])^(a[39] & b[12])^(a[38] & b[13])^(a[37] & b[14])^(a[36] & b[15])^(a[35] & b[16])^(a[34] & b[17])^(a[33] & b[18])^(a[32] & b[19])^(a[31] & b[20])^(a[30] & b[21])^(a[29] & b[22])^(a[28] & b[23])^(a[27] & b[24])^(a[26] & b[25])^(a[25] & b[26])^(a[24] & b[27])^(a[23] & b[28])^(a[22] & b[29])^(a[21] & b[30])^(a[20] & b[31])^(a[19] & b[32])^(a[18] & b[33])^(a[17] & b[34])^(a[16] & b[35])^(a[15] & b[36])^(a[14] & b[37])^(a[13] & b[38])^(a[12] & b[39])^(a[11] & b[40])^(a[10] & b[41])^(a[9] & b[42])^(a[8] & b[43])^(a[7] & b[44])^(a[6] & b[45])^(a[5] & b[46])^(a[4] & b[47])^(a[3] & b[48])^(a[2] & b[49])^(a[1] & b[50])^(a[0] & b[51]);
assign y[52] = (a[52] & b[0])^(a[51] & b[1])^(a[50] & b[2])^(a[49] & b[3])^(a[48] & b[4])^(a[47] & b[5])^(a[46] & b[6])^(a[45] & b[7])^(a[44] & b[8])^(a[43] & b[9])^(a[42] & b[10])^(a[41] & b[11])^(a[40] & b[12])^(a[39] & b[13])^(a[38] & b[14])^(a[37] & b[15])^(a[36] & b[16])^(a[35] & b[17])^(a[34] & b[18])^(a[33] & b[19])^(a[32] & b[20])^(a[31] & b[21])^(a[30] & b[22])^(a[29] & b[23])^(a[28] & b[24])^(a[27] & b[25])^(a[26] & b[26])^(a[25] & b[27])^(a[24] & b[28])^(a[23] & b[29])^(a[22] & b[30])^(a[21] & b[31])^(a[20] & b[32])^(a[19] & b[33])^(a[18] & b[34])^(a[17] & b[35])^(a[16] & b[36])^(a[15] & b[37])^(a[14] & b[38])^(a[13] & b[39])^(a[12] & b[40])^(a[11] & b[41])^(a[10] & b[42])^(a[9] & b[43])^(a[8] & b[44])^(a[7] & b[45])^(a[6] & b[46])^(a[5] & b[47])^(a[4] & b[48])^(a[3] & b[49])^(a[2] & b[50])^(a[1] & b[51])^(a[0] & b[52]);
assign y[53] = (a[53] & b[0])^(a[52] & b[1])^(a[51] & b[2])^(a[50] & b[3])^(a[49] & b[4])^(a[48] & b[5])^(a[47] & b[6])^(a[46] & b[7])^(a[45] & b[8])^(a[44] & b[9])^(a[43] & b[10])^(a[42] & b[11])^(a[41] & b[12])^(a[40] & b[13])^(a[39] & b[14])^(a[38] & b[15])^(a[37] & b[16])^(a[36] & b[17])^(a[35] & b[18])^(a[34] & b[19])^(a[33] & b[20])^(a[32] & b[21])^(a[31] & b[22])^(a[30] & b[23])^(a[29] & b[24])^(a[28] & b[25])^(a[27] & b[26])^(a[26] & b[27])^(a[25] & b[28])^(a[24] & b[29])^(a[23] & b[30])^(a[22] & b[31])^(a[21] & b[32])^(a[20] & b[33])^(a[19] & b[34])^(a[18] & b[35])^(a[17] & b[36])^(a[16] & b[37])^(a[15] & b[38])^(a[14] & b[39])^(a[13] & b[40])^(a[12] & b[41])^(a[11] & b[42])^(a[10] & b[43])^(a[9] & b[44])^(a[8] & b[45])^(a[7] & b[46])^(a[6] & b[47])^(a[5] & b[48])^(a[4] & b[49])^(a[3] & b[50])^(a[2] & b[51])^(a[1] & b[52])^(a[0] & b[53]);
assign y[54] = (a[54] & b[0])^(a[53] & b[1])^(a[52] & b[2])^(a[51] & b[3])^(a[50] & b[4])^(a[49] & b[5])^(a[48] & b[6])^(a[47] & b[7])^(a[46] & b[8])^(a[45] & b[9])^(a[44] & b[10])^(a[43] & b[11])^(a[42] & b[12])^(a[41] & b[13])^(a[40] & b[14])^(a[39] & b[15])^(a[38] & b[16])^(a[37] & b[17])^(a[36] & b[18])^(a[35] & b[19])^(a[34] & b[20])^(a[33] & b[21])^(a[32] & b[22])^(a[31] & b[23])^(a[30] & b[24])^(a[29] & b[25])^(a[28] & b[26])^(a[27] & b[27])^(a[26] & b[28])^(a[25] & b[29])^(a[24] & b[30])^(a[23] & b[31])^(a[22] & b[32])^(a[21] & b[33])^(a[20] & b[34])^(a[19] & b[35])^(a[18] & b[36])^(a[17] & b[37])^(a[16] & b[38])^(a[15] & b[39])^(a[14] & b[40])^(a[13] & b[41])^(a[12] & b[42])^(a[11] & b[43])^(a[10] & b[44])^(a[9] & b[45])^(a[8] & b[46])^(a[7] & b[47])^(a[6] & b[48])^(a[5] & b[49])^(a[4] & b[50])^(a[3] & b[51])^(a[2] & b[52])^(a[1] & b[53])^(a[0] & b[54]);
assign y[55] = (a[55] & b[0])^(a[54] & b[1])^(a[53] & b[2])^(a[52] & b[3])^(a[51] & b[4])^(a[50] & b[5])^(a[49] & b[6])^(a[48] & b[7])^(a[47] & b[8])^(a[46] & b[9])^(a[45] & b[10])^(a[44] & b[11])^(a[43] & b[12])^(a[42] & b[13])^(a[41] & b[14])^(a[40] & b[15])^(a[39] & b[16])^(a[38] & b[17])^(a[37] & b[18])^(a[36] & b[19])^(a[35] & b[20])^(a[34] & b[21])^(a[33] & b[22])^(a[32] & b[23])^(a[31] & b[24])^(a[30] & b[25])^(a[29] & b[26])^(a[28] & b[27])^(a[27] & b[28])^(a[26] & b[29])^(a[25] & b[30])^(a[24] & b[31])^(a[23] & b[32])^(a[22] & b[33])^(a[21] & b[34])^(a[20] & b[35])^(a[19] & b[36])^(a[18] & b[37])^(a[17] & b[38])^(a[16] & b[39])^(a[15] & b[40])^(a[14] & b[41])^(a[13] & b[42])^(a[12] & b[43])^(a[11] & b[44])^(a[10] & b[45])^(a[9] & b[46])^(a[8] & b[47])^(a[7] & b[48])^(a[6] & b[49])^(a[5] & b[50])^(a[4] & b[51])^(a[3] & b[52])^(a[2] & b[53])^(a[1] & b[54])^(a[0] & b[55]);
assign y[56] = (a[56] & b[0])^(a[55] & b[1])^(a[54] & b[2])^(a[53] & b[3])^(a[52] & b[4])^(a[51] & b[5])^(a[50] & b[6])^(a[49] & b[7])^(a[48] & b[8])^(a[47] & b[9])^(a[46] & b[10])^(a[45] & b[11])^(a[44] & b[12])^(a[43] & b[13])^(a[42] & b[14])^(a[41] & b[15])^(a[40] & b[16])^(a[39] & b[17])^(a[38] & b[18])^(a[37] & b[19])^(a[36] & b[20])^(a[35] & b[21])^(a[34] & b[22])^(a[33] & b[23])^(a[32] & b[24])^(a[31] & b[25])^(a[30] & b[26])^(a[29] & b[27])^(a[28] & b[28])^(a[27] & b[29])^(a[26] & b[30])^(a[25] & b[31])^(a[24] & b[32])^(a[23] & b[33])^(a[22] & b[34])^(a[21] & b[35])^(a[20] & b[36])^(a[19] & b[37])^(a[18] & b[38])^(a[17] & b[39])^(a[16] & b[40])^(a[15] & b[41])^(a[14] & b[42])^(a[13] & b[43])^(a[12] & b[44])^(a[11] & b[45])^(a[10] & b[46])^(a[9] & b[47])^(a[8] & b[48])^(a[7] & b[49])^(a[6] & b[50])^(a[5] & b[51])^(a[4] & b[52])^(a[3] & b[53])^(a[2] & b[54])^(a[1] & b[55])^(a[0] & b[56]);
assign y[57] = (a[57] & b[0])^(a[56] & b[1])^(a[55] & b[2])^(a[54] & b[3])^(a[53] & b[4])^(a[52] & b[5])^(a[51] & b[6])^(a[50] & b[7])^(a[49] & b[8])^(a[48] & b[9])^(a[47] & b[10])^(a[46] & b[11])^(a[45] & b[12])^(a[44] & b[13])^(a[43] & b[14])^(a[42] & b[15])^(a[41] & b[16])^(a[40] & b[17])^(a[39] & b[18])^(a[38] & b[19])^(a[37] & b[20])^(a[36] & b[21])^(a[35] & b[22])^(a[34] & b[23])^(a[33] & b[24])^(a[32] & b[25])^(a[31] & b[26])^(a[30] & b[27])^(a[29] & b[28])^(a[28] & b[29])^(a[27] & b[30])^(a[26] & b[31])^(a[25] & b[32])^(a[24] & b[33])^(a[23] & b[34])^(a[22] & b[35])^(a[21] & b[36])^(a[20] & b[37])^(a[19] & b[38])^(a[18] & b[39])^(a[17] & b[40])^(a[16] & b[41])^(a[15] & b[42])^(a[14] & b[43])^(a[13] & b[44])^(a[12] & b[45])^(a[11] & b[46])^(a[10] & b[47])^(a[9] & b[48])^(a[8] & b[49])^(a[7] & b[50])^(a[6] & b[51])^(a[5] & b[52])^(a[4] & b[53])^(a[3] & b[54])^(a[2] & b[55])^(a[1] & b[56])^(a[0] & b[57]);
assign y[58] = (a[58] & b[0])^(a[57] & b[1])^(a[56] & b[2])^(a[55] & b[3])^(a[54] & b[4])^(a[53] & b[5])^(a[52] & b[6])^(a[51] & b[7])^(a[50] & b[8])^(a[49] & b[9])^(a[48] & b[10])^(a[47] & b[11])^(a[46] & b[12])^(a[45] & b[13])^(a[44] & b[14])^(a[43] & b[15])^(a[42] & b[16])^(a[41] & b[17])^(a[40] & b[18])^(a[39] & b[19])^(a[38] & b[20])^(a[37] & b[21])^(a[36] & b[22])^(a[35] & b[23])^(a[34] & b[24])^(a[33] & b[25])^(a[32] & b[26])^(a[31] & b[27])^(a[30] & b[28])^(a[29] & b[29])^(a[28] & b[30])^(a[27] & b[31])^(a[26] & b[32])^(a[25] & b[33])^(a[24] & b[34])^(a[23] & b[35])^(a[22] & b[36])^(a[21] & b[37])^(a[20] & b[38])^(a[19] & b[39])^(a[18] & b[40])^(a[17] & b[41])^(a[16] & b[42])^(a[15] & b[43])^(a[14] & b[44])^(a[13] & b[45])^(a[12] & b[46])^(a[11] & b[47])^(a[10] & b[48])^(a[9] & b[49])^(a[8] & b[50])^(a[7] & b[51])^(a[6] & b[52])^(a[5] & b[53])^(a[4] & b[54])^(a[3] & b[55])^(a[2] & b[56])^(a[1] & b[57])^(a[0] & b[58]);
assign y[59] = (a[59] & b[0])^(a[58] & b[1])^(a[57] & b[2])^(a[56] & b[3])^(a[55] & b[4])^(a[54] & b[5])^(a[53] & b[6])^(a[52] & b[7])^(a[51] & b[8])^(a[50] & b[9])^(a[49] & b[10])^(a[48] & b[11])^(a[47] & b[12])^(a[46] & b[13])^(a[45] & b[14])^(a[44] & b[15])^(a[43] & b[16])^(a[42] & b[17])^(a[41] & b[18])^(a[40] & b[19])^(a[39] & b[20])^(a[38] & b[21])^(a[37] & b[22])^(a[36] & b[23])^(a[35] & b[24])^(a[34] & b[25])^(a[33] & b[26])^(a[32] & b[27])^(a[31] & b[28])^(a[30] & b[29])^(a[29] & b[30])^(a[28] & b[31])^(a[27] & b[32])^(a[26] & b[33])^(a[25] & b[34])^(a[24] & b[35])^(a[23] & b[36])^(a[22] & b[37])^(a[21] & b[38])^(a[20] & b[39])^(a[19] & b[40])^(a[18] & b[41])^(a[17] & b[42])^(a[16] & b[43])^(a[15] & b[44])^(a[14] & b[45])^(a[13] & b[46])^(a[12] & b[47])^(a[11] & b[48])^(a[10] & b[49])^(a[9] & b[50])^(a[8] & b[51])^(a[7] & b[52])^(a[6] & b[53])^(a[5] & b[54])^(a[4] & b[55])^(a[3] & b[56])^(a[2] & b[57])^(a[1] & b[58])^(a[0] & b[59]);
assign y[60] = (a[60] & b[0])^(a[59] & b[1])^(a[58] & b[2])^(a[57] & b[3])^(a[56] & b[4])^(a[55] & b[5])^(a[54] & b[6])^(a[53] & b[7])^(a[52] & b[8])^(a[51] & b[9])^(a[50] & b[10])^(a[49] & b[11])^(a[48] & b[12])^(a[47] & b[13])^(a[46] & b[14])^(a[45] & b[15])^(a[44] & b[16])^(a[43] & b[17])^(a[42] & b[18])^(a[41] & b[19])^(a[40] & b[20])^(a[39] & b[21])^(a[38] & b[22])^(a[37] & b[23])^(a[36] & b[24])^(a[35] & b[25])^(a[34] & b[26])^(a[33] & b[27])^(a[32] & b[28])^(a[31] & b[29])^(a[30] & b[30])^(a[29] & b[31])^(a[28] & b[32])^(a[27] & b[33])^(a[26] & b[34])^(a[25] & b[35])^(a[24] & b[36])^(a[23] & b[37])^(a[22] & b[38])^(a[21] & b[39])^(a[20] & b[40])^(a[19] & b[41])^(a[18] & b[42])^(a[17] & b[43])^(a[16] & b[44])^(a[15] & b[45])^(a[14] & b[46])^(a[13] & b[47])^(a[12] & b[48])^(a[11] & b[49])^(a[10] & b[50])^(a[9] & b[51])^(a[8] & b[52])^(a[7] & b[53])^(a[6] & b[54])^(a[5] & b[55])^(a[4] & b[56])^(a[3] & b[57])^(a[2] & b[58])^(a[1] & b[59])^(a[0] & b[60]);
assign y[61] = (a[61] & b[0])^(a[60] & b[1])^(a[59] & b[2])^(a[58] & b[3])^(a[57] & b[4])^(a[56] & b[5])^(a[55] & b[6])^(a[54] & b[7])^(a[53] & b[8])^(a[52] & b[9])^(a[51] & b[10])^(a[50] & b[11])^(a[49] & b[12])^(a[48] & b[13])^(a[47] & b[14])^(a[46] & b[15])^(a[45] & b[16])^(a[44] & b[17])^(a[43] & b[18])^(a[42] & b[19])^(a[41] & b[20])^(a[40] & b[21])^(a[39] & b[22])^(a[38] & b[23])^(a[37] & b[24])^(a[36] & b[25])^(a[35] & b[26])^(a[34] & b[27])^(a[33] & b[28])^(a[32] & b[29])^(a[31] & b[30])^(a[30] & b[31])^(a[29] & b[32])^(a[28] & b[33])^(a[27] & b[34])^(a[26] & b[35])^(a[25] & b[36])^(a[24] & b[37])^(a[23] & b[38])^(a[22] & b[39])^(a[21] & b[40])^(a[20] & b[41])^(a[19] & b[42])^(a[18] & b[43])^(a[17] & b[44])^(a[16] & b[45])^(a[15] & b[46])^(a[14] & b[47])^(a[13] & b[48])^(a[12] & b[49])^(a[11] & b[50])^(a[10] & b[51])^(a[9] & b[52])^(a[8] & b[53])^(a[7] & b[54])^(a[6] & b[55])^(a[5] & b[56])^(a[4] & b[57])^(a[3] & b[58])^(a[2] & b[59])^(a[1] & b[60])^(a[0] & b[61]);
assign y[62] = (a[62] & b[0])^(a[61] & b[1])^(a[60] & b[2])^(a[59] & b[3])^(a[58] & b[4])^(a[57] & b[5])^(a[56] & b[6])^(a[55] & b[7])^(a[54] & b[8])^(a[53] & b[9])^(a[52] & b[10])^(a[51] & b[11])^(a[50] & b[12])^(a[49] & b[13])^(a[48] & b[14])^(a[47] & b[15])^(a[46] & b[16])^(a[45] & b[17])^(a[44] & b[18])^(a[43] & b[19])^(a[42] & b[20])^(a[41] & b[21])^(a[40] & b[22])^(a[39] & b[23])^(a[38] & b[24])^(a[37] & b[25])^(a[36] & b[26])^(a[35] & b[27])^(a[34] & b[28])^(a[33] & b[29])^(a[32] & b[30])^(a[31] & b[31])^(a[30] & b[32])^(a[29] & b[33])^(a[28] & b[34])^(a[27] & b[35])^(a[26] & b[36])^(a[25] & b[37])^(a[24] & b[38])^(a[23] & b[39])^(a[22] & b[40])^(a[21] & b[41])^(a[20] & b[42])^(a[19] & b[43])^(a[18] & b[44])^(a[17] & b[45])^(a[16] & b[46])^(a[15] & b[47])^(a[14] & b[48])^(a[13] & b[49])^(a[12] & b[50])^(a[11] & b[51])^(a[10] & b[52])^(a[9] & b[53])^(a[8] & b[54])^(a[7] & b[55])^(a[6] & b[56])^(a[5] & b[57])^(a[4] & b[58])^(a[3] & b[59])^(a[2] & b[60])^(a[1] & b[61])^(a[0] & b[62]);
assign y[63] = (a[63] & b[0])^(a[62] & b[1])^(a[61] & b[2])^(a[60] & b[3])^(a[59] & b[4])^(a[58] & b[5])^(a[57] & b[6])^(a[56] & b[7])^(a[55] & b[8])^(a[54] & b[9])^(a[53] & b[10])^(a[52] & b[11])^(a[51] & b[12])^(a[50] & b[13])^(a[49] & b[14])^(a[48] & b[15])^(a[47] & b[16])^(a[46] & b[17])^(a[45] & b[18])^(a[44] & b[19])^(a[43] & b[20])^(a[42] & b[21])^(a[41] & b[22])^(a[40] & b[23])^(a[39] & b[24])^(a[38] & b[25])^(a[37] & b[26])^(a[36] & b[27])^(a[35] & b[28])^(a[34] & b[29])^(a[33] & b[30])^(a[32] & b[31])^(a[31] & b[32])^(a[30] & b[33])^(a[29] & b[34])^(a[28] & b[35])^(a[27] & b[36])^(a[26] & b[37])^(a[25] & b[38])^(a[24] & b[39])^(a[23] & b[40])^(a[22] & b[41])^(a[21] & b[42])^(a[20] & b[43])^(a[19] & b[44])^(a[18] & b[45])^(a[17] & b[46])^(a[16] & b[47])^(a[15] & b[48])^(a[14] & b[49])^(a[13] & b[50])^(a[12] & b[51])^(a[11] & b[52])^(a[10] & b[53])^(a[9] & b[54])^(a[8] & b[55])^(a[7] & b[56])^(a[6] & b[57])^(a[5] & b[58])^(a[4] & b[59])^(a[3] & b[60])^(a[2] & b[61])^(a[1] & b[62])^(a[0] & b[63]);
assign y[64] = (a[64] & b[0])^(a[63] & b[1])^(a[62] & b[2])^(a[61] & b[3])^(a[60] & b[4])^(a[59] & b[5])^(a[58] & b[6])^(a[57] & b[7])^(a[56] & b[8])^(a[55] & b[9])^(a[54] & b[10])^(a[53] & b[11])^(a[52] & b[12])^(a[51] & b[13])^(a[50] & b[14])^(a[49] & b[15])^(a[48] & b[16])^(a[47] & b[17])^(a[46] & b[18])^(a[45] & b[19])^(a[44] & b[20])^(a[43] & b[21])^(a[42] & b[22])^(a[41] & b[23])^(a[40] & b[24])^(a[39] & b[25])^(a[38] & b[26])^(a[37] & b[27])^(a[36] & b[28])^(a[35] & b[29])^(a[34] & b[30])^(a[33] & b[31])^(a[32] & b[32])^(a[31] & b[33])^(a[30] & b[34])^(a[29] & b[35])^(a[28] & b[36])^(a[27] & b[37])^(a[26] & b[38])^(a[25] & b[39])^(a[24] & b[40])^(a[23] & b[41])^(a[22] & b[42])^(a[21] & b[43])^(a[20] & b[44])^(a[19] & b[45])^(a[18] & b[46])^(a[17] & b[47])^(a[16] & b[48])^(a[15] & b[49])^(a[14] & b[50])^(a[13] & b[51])^(a[12] & b[52])^(a[11] & b[53])^(a[10] & b[54])^(a[9] & b[55])^(a[8] & b[56])^(a[7] & b[57])^(a[6] & b[58])^(a[5] & b[59])^(a[4] & b[60])^(a[3] & b[61])^(a[2] & b[62])^(a[1] & b[63])^(a[0] & b[64]);
assign y[65] = (a[65] & b[0])^(a[64] & b[1])^(a[63] & b[2])^(a[62] & b[3])^(a[61] & b[4])^(a[60] & b[5])^(a[59] & b[6])^(a[58] & b[7])^(a[57] & b[8])^(a[56] & b[9])^(a[55] & b[10])^(a[54] & b[11])^(a[53] & b[12])^(a[52] & b[13])^(a[51] & b[14])^(a[50] & b[15])^(a[49] & b[16])^(a[48] & b[17])^(a[47] & b[18])^(a[46] & b[19])^(a[45] & b[20])^(a[44] & b[21])^(a[43] & b[22])^(a[42] & b[23])^(a[41] & b[24])^(a[40] & b[25])^(a[39] & b[26])^(a[38] & b[27])^(a[37] & b[28])^(a[36] & b[29])^(a[35] & b[30])^(a[34] & b[31])^(a[33] & b[32])^(a[32] & b[33])^(a[31] & b[34])^(a[30] & b[35])^(a[29] & b[36])^(a[28] & b[37])^(a[27] & b[38])^(a[26] & b[39])^(a[25] & b[40])^(a[24] & b[41])^(a[23] & b[42])^(a[22] & b[43])^(a[21] & b[44])^(a[20] & b[45])^(a[19] & b[46])^(a[18] & b[47])^(a[17] & b[48])^(a[16] & b[49])^(a[15] & b[50])^(a[14] & b[51])^(a[13] & b[52])^(a[12] & b[53])^(a[11] & b[54])^(a[10] & b[55])^(a[9] & b[56])^(a[8] & b[57])^(a[7] & b[58])^(a[6] & b[59])^(a[5] & b[60])^(a[4] & b[61])^(a[3] & b[62])^(a[2] & b[63])^(a[1] & b[64])^(a[0] & b[65]);
assign y[66] = (a[66] & b[0])^(a[65] & b[1])^(a[64] & b[2])^(a[63] & b[3])^(a[62] & b[4])^(a[61] & b[5])^(a[60] & b[6])^(a[59] & b[7])^(a[58] & b[8])^(a[57] & b[9])^(a[56] & b[10])^(a[55] & b[11])^(a[54] & b[12])^(a[53] & b[13])^(a[52] & b[14])^(a[51] & b[15])^(a[50] & b[16])^(a[49] & b[17])^(a[48] & b[18])^(a[47] & b[19])^(a[46] & b[20])^(a[45] & b[21])^(a[44] & b[22])^(a[43] & b[23])^(a[42] & b[24])^(a[41] & b[25])^(a[40] & b[26])^(a[39] & b[27])^(a[38] & b[28])^(a[37] & b[29])^(a[36] & b[30])^(a[35] & b[31])^(a[34] & b[32])^(a[33] & b[33])^(a[32] & b[34])^(a[31] & b[35])^(a[30] & b[36])^(a[29] & b[37])^(a[28] & b[38])^(a[27] & b[39])^(a[26] & b[40])^(a[25] & b[41])^(a[24] & b[42])^(a[23] & b[43])^(a[22] & b[44])^(a[21] & b[45])^(a[20] & b[46])^(a[19] & b[47])^(a[18] & b[48])^(a[17] & b[49])^(a[16] & b[50])^(a[15] & b[51])^(a[14] & b[52])^(a[13] & b[53])^(a[12] & b[54])^(a[11] & b[55])^(a[10] & b[56])^(a[9] & b[57])^(a[8] & b[58])^(a[7] & b[59])^(a[6] & b[60])^(a[5] & b[61])^(a[4] & b[62])^(a[3] & b[63])^(a[2] & b[64])^(a[1] & b[65])^(a[0] & b[66]);
assign y[67] = (a[67] & b[0])^(a[66] & b[1])^(a[65] & b[2])^(a[64] & b[3])^(a[63] & b[4])^(a[62] & b[5])^(a[61] & b[6])^(a[60] & b[7])^(a[59] & b[8])^(a[58] & b[9])^(a[57] & b[10])^(a[56] & b[11])^(a[55] & b[12])^(a[54] & b[13])^(a[53] & b[14])^(a[52] & b[15])^(a[51] & b[16])^(a[50] & b[17])^(a[49] & b[18])^(a[48] & b[19])^(a[47] & b[20])^(a[46] & b[21])^(a[45] & b[22])^(a[44] & b[23])^(a[43] & b[24])^(a[42] & b[25])^(a[41] & b[26])^(a[40] & b[27])^(a[39] & b[28])^(a[38] & b[29])^(a[37] & b[30])^(a[36] & b[31])^(a[35] & b[32])^(a[34] & b[33])^(a[33] & b[34])^(a[32] & b[35])^(a[31] & b[36])^(a[30] & b[37])^(a[29] & b[38])^(a[28] & b[39])^(a[27] & b[40])^(a[26] & b[41])^(a[25] & b[42])^(a[24] & b[43])^(a[23] & b[44])^(a[22] & b[45])^(a[21] & b[46])^(a[20] & b[47])^(a[19] & b[48])^(a[18] & b[49])^(a[17] & b[50])^(a[16] & b[51])^(a[15] & b[52])^(a[14] & b[53])^(a[13] & b[54])^(a[12] & b[55])^(a[11] & b[56])^(a[10] & b[57])^(a[9] & b[58])^(a[8] & b[59])^(a[7] & b[60])^(a[6] & b[61])^(a[5] & b[62])^(a[4] & b[63])^(a[3] & b[64])^(a[2] & b[65])^(a[1] & b[66])^(a[0] & b[67]);
assign y[68] = (a[68] & b[0])^(a[67] & b[1])^(a[66] & b[2])^(a[65] & b[3])^(a[64] & b[4])^(a[63] & b[5])^(a[62] & b[6])^(a[61] & b[7])^(a[60] & b[8])^(a[59] & b[9])^(a[58] & b[10])^(a[57] & b[11])^(a[56] & b[12])^(a[55] & b[13])^(a[54] & b[14])^(a[53] & b[15])^(a[52] & b[16])^(a[51] & b[17])^(a[50] & b[18])^(a[49] & b[19])^(a[48] & b[20])^(a[47] & b[21])^(a[46] & b[22])^(a[45] & b[23])^(a[44] & b[24])^(a[43] & b[25])^(a[42] & b[26])^(a[41] & b[27])^(a[40] & b[28])^(a[39] & b[29])^(a[38] & b[30])^(a[37] & b[31])^(a[36] & b[32])^(a[35] & b[33])^(a[34] & b[34])^(a[33] & b[35])^(a[32] & b[36])^(a[31] & b[37])^(a[30] & b[38])^(a[29] & b[39])^(a[28] & b[40])^(a[27] & b[41])^(a[26] & b[42])^(a[25] & b[43])^(a[24] & b[44])^(a[23] & b[45])^(a[22] & b[46])^(a[21] & b[47])^(a[20] & b[48])^(a[19] & b[49])^(a[18] & b[50])^(a[17] & b[51])^(a[16] & b[52])^(a[15] & b[53])^(a[14] & b[54])^(a[13] & b[55])^(a[12] & b[56])^(a[11] & b[57])^(a[10] & b[58])^(a[9] & b[59])^(a[8] & b[60])^(a[7] & b[61])^(a[6] & b[62])^(a[5] & b[63])^(a[4] & b[64])^(a[3] & b[65])^(a[2] & b[66])^(a[1] & b[67])^(a[0] & b[68]);
assign y[69] = (a[69] & b[0])^(a[68] & b[1])^(a[67] & b[2])^(a[66] & b[3])^(a[65] & b[4])^(a[64] & b[5])^(a[63] & b[6])^(a[62] & b[7])^(a[61] & b[8])^(a[60] & b[9])^(a[59] & b[10])^(a[58] & b[11])^(a[57] & b[12])^(a[56] & b[13])^(a[55] & b[14])^(a[54] & b[15])^(a[53] & b[16])^(a[52] & b[17])^(a[51] & b[18])^(a[50] & b[19])^(a[49] & b[20])^(a[48] & b[21])^(a[47] & b[22])^(a[46] & b[23])^(a[45] & b[24])^(a[44] & b[25])^(a[43] & b[26])^(a[42] & b[27])^(a[41] & b[28])^(a[40] & b[29])^(a[39] & b[30])^(a[38] & b[31])^(a[37] & b[32])^(a[36] & b[33])^(a[35] & b[34])^(a[34] & b[35])^(a[33] & b[36])^(a[32] & b[37])^(a[31] & b[38])^(a[30] & b[39])^(a[29] & b[40])^(a[28] & b[41])^(a[27] & b[42])^(a[26] & b[43])^(a[25] & b[44])^(a[24] & b[45])^(a[23] & b[46])^(a[22] & b[47])^(a[21] & b[48])^(a[20] & b[49])^(a[19] & b[50])^(a[18] & b[51])^(a[17] & b[52])^(a[16] & b[53])^(a[15] & b[54])^(a[14] & b[55])^(a[13] & b[56])^(a[12] & b[57])^(a[11] & b[58])^(a[10] & b[59])^(a[9] & b[60])^(a[8] & b[61])^(a[7] & b[62])^(a[6] & b[63])^(a[5] & b[64])^(a[4] & b[65])^(a[3] & b[66])^(a[2] & b[67])^(a[1] & b[68])^(a[0] & b[69]);
assign y[70] = (a[70] & b[0])^(a[69] & b[1])^(a[68] & b[2])^(a[67] & b[3])^(a[66] & b[4])^(a[65] & b[5])^(a[64] & b[6])^(a[63] & b[7])^(a[62] & b[8])^(a[61] & b[9])^(a[60] & b[10])^(a[59] & b[11])^(a[58] & b[12])^(a[57] & b[13])^(a[56] & b[14])^(a[55] & b[15])^(a[54] & b[16])^(a[53] & b[17])^(a[52] & b[18])^(a[51] & b[19])^(a[50] & b[20])^(a[49] & b[21])^(a[48] & b[22])^(a[47] & b[23])^(a[46] & b[24])^(a[45] & b[25])^(a[44] & b[26])^(a[43] & b[27])^(a[42] & b[28])^(a[41] & b[29])^(a[40] & b[30])^(a[39] & b[31])^(a[38] & b[32])^(a[37] & b[33])^(a[36] & b[34])^(a[35] & b[35])^(a[34] & b[36])^(a[33] & b[37])^(a[32] & b[38])^(a[31] & b[39])^(a[30] & b[40])^(a[29] & b[41])^(a[28] & b[42])^(a[27] & b[43])^(a[26] & b[44])^(a[25] & b[45])^(a[24] & b[46])^(a[23] & b[47])^(a[22] & b[48])^(a[21] & b[49])^(a[20] & b[50])^(a[19] & b[51])^(a[18] & b[52])^(a[17] & b[53])^(a[16] & b[54])^(a[15] & b[55])^(a[14] & b[56])^(a[13] & b[57])^(a[12] & b[58])^(a[11] & b[59])^(a[10] & b[60])^(a[9] & b[61])^(a[8] & b[62])^(a[7] & b[63])^(a[6] & b[64])^(a[5] & b[65])^(a[4] & b[66])^(a[3] & b[67])^(a[2] & b[68])^(a[1] & b[69])^(a[0] & b[70]);
assign y[71] = (a[71] & b[0])^(a[70] & b[1])^(a[69] & b[2])^(a[68] & b[3])^(a[67] & b[4])^(a[66] & b[5])^(a[65] & b[6])^(a[64] & b[7])^(a[63] & b[8])^(a[62] & b[9])^(a[61] & b[10])^(a[60] & b[11])^(a[59] & b[12])^(a[58] & b[13])^(a[57] & b[14])^(a[56] & b[15])^(a[55] & b[16])^(a[54] & b[17])^(a[53] & b[18])^(a[52] & b[19])^(a[51] & b[20])^(a[50] & b[21])^(a[49] & b[22])^(a[48] & b[23])^(a[47] & b[24])^(a[46] & b[25])^(a[45] & b[26])^(a[44] & b[27])^(a[43] & b[28])^(a[42] & b[29])^(a[41] & b[30])^(a[40] & b[31])^(a[39] & b[32])^(a[38] & b[33])^(a[37] & b[34])^(a[36] & b[35])^(a[35] & b[36])^(a[34] & b[37])^(a[33] & b[38])^(a[32] & b[39])^(a[31] & b[40])^(a[30] & b[41])^(a[29] & b[42])^(a[28] & b[43])^(a[27] & b[44])^(a[26] & b[45])^(a[25] & b[46])^(a[24] & b[47])^(a[23] & b[48])^(a[22] & b[49])^(a[21] & b[50])^(a[20] & b[51])^(a[19] & b[52])^(a[18] & b[53])^(a[17] & b[54])^(a[16] & b[55])^(a[15] & b[56])^(a[14] & b[57])^(a[13] & b[58])^(a[12] & b[59])^(a[11] & b[60])^(a[10] & b[61])^(a[9] & b[62])^(a[8] & b[63])^(a[7] & b[64])^(a[6] & b[65])^(a[5] & b[66])^(a[4] & b[67])^(a[3] & b[68])^(a[2] & b[69])^(a[1] & b[70])^(a[0] & b[71]);
assign y[72] = (a[72] & b[0])^(a[71] & b[1])^(a[70] & b[2])^(a[69] & b[3])^(a[68] & b[4])^(a[67] & b[5])^(a[66] & b[6])^(a[65] & b[7])^(a[64] & b[8])^(a[63] & b[9])^(a[62] & b[10])^(a[61] & b[11])^(a[60] & b[12])^(a[59] & b[13])^(a[58] & b[14])^(a[57] & b[15])^(a[56] & b[16])^(a[55] & b[17])^(a[54] & b[18])^(a[53] & b[19])^(a[52] & b[20])^(a[51] & b[21])^(a[50] & b[22])^(a[49] & b[23])^(a[48] & b[24])^(a[47] & b[25])^(a[46] & b[26])^(a[45] & b[27])^(a[44] & b[28])^(a[43] & b[29])^(a[42] & b[30])^(a[41] & b[31])^(a[40] & b[32])^(a[39] & b[33])^(a[38] & b[34])^(a[37] & b[35])^(a[36] & b[36])^(a[35] & b[37])^(a[34] & b[38])^(a[33] & b[39])^(a[32] & b[40])^(a[31] & b[41])^(a[30] & b[42])^(a[29] & b[43])^(a[28] & b[44])^(a[27] & b[45])^(a[26] & b[46])^(a[25] & b[47])^(a[24] & b[48])^(a[23] & b[49])^(a[22] & b[50])^(a[21] & b[51])^(a[20] & b[52])^(a[19] & b[53])^(a[18] & b[54])^(a[17] & b[55])^(a[16] & b[56])^(a[15] & b[57])^(a[14] & b[58])^(a[13] & b[59])^(a[12] & b[60])^(a[11] & b[61])^(a[10] & b[62])^(a[9] & b[63])^(a[8] & b[64])^(a[7] & b[65])^(a[6] & b[66])^(a[5] & b[67])^(a[4] & b[68])^(a[3] & b[69])^(a[2] & b[70])^(a[1] & b[71])^(a[0] & b[72]);
assign y[73] = (a[73] & b[0])^(a[72] & b[1])^(a[71] & b[2])^(a[70] & b[3])^(a[69] & b[4])^(a[68] & b[5])^(a[67] & b[6])^(a[66] & b[7])^(a[65] & b[8])^(a[64] & b[9])^(a[63] & b[10])^(a[62] & b[11])^(a[61] & b[12])^(a[60] & b[13])^(a[59] & b[14])^(a[58] & b[15])^(a[57] & b[16])^(a[56] & b[17])^(a[55] & b[18])^(a[54] & b[19])^(a[53] & b[20])^(a[52] & b[21])^(a[51] & b[22])^(a[50] & b[23])^(a[49] & b[24])^(a[48] & b[25])^(a[47] & b[26])^(a[46] & b[27])^(a[45] & b[28])^(a[44] & b[29])^(a[43] & b[30])^(a[42] & b[31])^(a[41] & b[32])^(a[40] & b[33])^(a[39] & b[34])^(a[38] & b[35])^(a[37] & b[36])^(a[36] & b[37])^(a[35] & b[38])^(a[34] & b[39])^(a[33] & b[40])^(a[32] & b[41])^(a[31] & b[42])^(a[30] & b[43])^(a[29] & b[44])^(a[28] & b[45])^(a[27] & b[46])^(a[26] & b[47])^(a[25] & b[48])^(a[24] & b[49])^(a[23] & b[50])^(a[22] & b[51])^(a[21] & b[52])^(a[20] & b[53])^(a[19] & b[54])^(a[18] & b[55])^(a[17] & b[56])^(a[16] & b[57])^(a[15] & b[58])^(a[14] & b[59])^(a[13] & b[60])^(a[12] & b[61])^(a[11] & b[62])^(a[10] & b[63])^(a[9] & b[64])^(a[8] & b[65])^(a[7] & b[66])^(a[6] & b[67])^(a[5] & b[68])^(a[4] & b[69])^(a[3] & b[70])^(a[2] & b[71])^(a[1] & b[72])^(a[0] & b[73]);
assign y[74] = (a[74] & b[0])^(a[73] & b[1])^(a[72] & b[2])^(a[71] & b[3])^(a[70] & b[4])^(a[69] & b[5])^(a[68] & b[6])^(a[67] & b[7])^(a[66] & b[8])^(a[65] & b[9])^(a[64] & b[10])^(a[63] & b[11])^(a[62] & b[12])^(a[61] & b[13])^(a[60] & b[14])^(a[59] & b[15])^(a[58] & b[16])^(a[57] & b[17])^(a[56] & b[18])^(a[55] & b[19])^(a[54] & b[20])^(a[53] & b[21])^(a[52] & b[22])^(a[51] & b[23])^(a[50] & b[24])^(a[49] & b[25])^(a[48] & b[26])^(a[47] & b[27])^(a[46] & b[28])^(a[45] & b[29])^(a[44] & b[30])^(a[43] & b[31])^(a[42] & b[32])^(a[41] & b[33])^(a[40] & b[34])^(a[39] & b[35])^(a[38] & b[36])^(a[37] & b[37])^(a[36] & b[38])^(a[35] & b[39])^(a[34] & b[40])^(a[33] & b[41])^(a[32] & b[42])^(a[31] & b[43])^(a[30] & b[44])^(a[29] & b[45])^(a[28] & b[46])^(a[27] & b[47])^(a[26] & b[48])^(a[25] & b[49])^(a[24] & b[50])^(a[23] & b[51])^(a[22] & b[52])^(a[21] & b[53])^(a[20] & b[54])^(a[19] & b[55])^(a[18] & b[56])^(a[17] & b[57])^(a[16] & b[58])^(a[15] & b[59])^(a[14] & b[60])^(a[13] & b[61])^(a[12] & b[62])^(a[11] & b[63])^(a[10] & b[64])^(a[9] & b[65])^(a[8] & b[66])^(a[7] & b[67])^(a[6] & b[68])^(a[5] & b[69])^(a[4] & b[70])^(a[3] & b[71])^(a[2] & b[72])^(a[1] & b[73])^(a[0] & b[74]);
assign y[75] = (a[75] & b[0])^(a[74] & b[1])^(a[73] & b[2])^(a[72] & b[3])^(a[71] & b[4])^(a[70] & b[5])^(a[69] & b[6])^(a[68] & b[7])^(a[67] & b[8])^(a[66] & b[9])^(a[65] & b[10])^(a[64] & b[11])^(a[63] & b[12])^(a[62] & b[13])^(a[61] & b[14])^(a[60] & b[15])^(a[59] & b[16])^(a[58] & b[17])^(a[57] & b[18])^(a[56] & b[19])^(a[55] & b[20])^(a[54] & b[21])^(a[53] & b[22])^(a[52] & b[23])^(a[51] & b[24])^(a[50] & b[25])^(a[49] & b[26])^(a[48] & b[27])^(a[47] & b[28])^(a[46] & b[29])^(a[45] & b[30])^(a[44] & b[31])^(a[43] & b[32])^(a[42] & b[33])^(a[41] & b[34])^(a[40] & b[35])^(a[39] & b[36])^(a[38] & b[37])^(a[37] & b[38])^(a[36] & b[39])^(a[35] & b[40])^(a[34] & b[41])^(a[33] & b[42])^(a[32] & b[43])^(a[31] & b[44])^(a[30] & b[45])^(a[29] & b[46])^(a[28] & b[47])^(a[27] & b[48])^(a[26] & b[49])^(a[25] & b[50])^(a[24] & b[51])^(a[23] & b[52])^(a[22] & b[53])^(a[21] & b[54])^(a[20] & b[55])^(a[19] & b[56])^(a[18] & b[57])^(a[17] & b[58])^(a[16] & b[59])^(a[15] & b[60])^(a[14] & b[61])^(a[13] & b[62])^(a[12] & b[63])^(a[11] & b[64])^(a[10] & b[65])^(a[9] & b[66])^(a[8] & b[67])^(a[7] & b[68])^(a[6] & b[69])^(a[5] & b[70])^(a[4] & b[71])^(a[3] & b[72])^(a[2] & b[73])^(a[1] & b[74])^(a[0] & b[75]);
assign y[76] = (a[76] & b[0])^(a[75] & b[1])^(a[74] & b[2])^(a[73] & b[3])^(a[72] & b[4])^(a[71] & b[5])^(a[70] & b[6])^(a[69] & b[7])^(a[68] & b[8])^(a[67] & b[9])^(a[66] & b[10])^(a[65] & b[11])^(a[64] & b[12])^(a[63] & b[13])^(a[62] & b[14])^(a[61] & b[15])^(a[60] & b[16])^(a[59] & b[17])^(a[58] & b[18])^(a[57] & b[19])^(a[56] & b[20])^(a[55] & b[21])^(a[54] & b[22])^(a[53] & b[23])^(a[52] & b[24])^(a[51] & b[25])^(a[50] & b[26])^(a[49] & b[27])^(a[48] & b[28])^(a[47] & b[29])^(a[46] & b[30])^(a[45] & b[31])^(a[44] & b[32])^(a[43] & b[33])^(a[42] & b[34])^(a[41] & b[35])^(a[40] & b[36])^(a[39] & b[37])^(a[38] & b[38])^(a[37] & b[39])^(a[36] & b[40])^(a[35] & b[41])^(a[34] & b[42])^(a[33] & b[43])^(a[32] & b[44])^(a[31] & b[45])^(a[30] & b[46])^(a[29] & b[47])^(a[28] & b[48])^(a[27] & b[49])^(a[26] & b[50])^(a[25] & b[51])^(a[24] & b[52])^(a[23] & b[53])^(a[22] & b[54])^(a[21] & b[55])^(a[20] & b[56])^(a[19] & b[57])^(a[18] & b[58])^(a[17] & b[59])^(a[16] & b[60])^(a[15] & b[61])^(a[14] & b[62])^(a[13] & b[63])^(a[12] & b[64])^(a[11] & b[65])^(a[10] & b[66])^(a[9] & b[67])^(a[8] & b[68])^(a[7] & b[69])^(a[6] & b[70])^(a[5] & b[71])^(a[4] & b[72])^(a[3] & b[73])^(a[2] & b[74])^(a[1] & b[75])^(a[0] & b[76]);
assign y[77] = (a[77] & b[0])^(a[76] & b[1])^(a[75] & b[2])^(a[74] & b[3])^(a[73] & b[4])^(a[72] & b[5])^(a[71] & b[6])^(a[70] & b[7])^(a[69] & b[8])^(a[68] & b[9])^(a[67] & b[10])^(a[66] & b[11])^(a[65] & b[12])^(a[64] & b[13])^(a[63] & b[14])^(a[62] & b[15])^(a[61] & b[16])^(a[60] & b[17])^(a[59] & b[18])^(a[58] & b[19])^(a[57] & b[20])^(a[56] & b[21])^(a[55] & b[22])^(a[54] & b[23])^(a[53] & b[24])^(a[52] & b[25])^(a[51] & b[26])^(a[50] & b[27])^(a[49] & b[28])^(a[48] & b[29])^(a[47] & b[30])^(a[46] & b[31])^(a[45] & b[32])^(a[44] & b[33])^(a[43] & b[34])^(a[42] & b[35])^(a[41] & b[36])^(a[40] & b[37])^(a[39] & b[38])^(a[38] & b[39])^(a[37] & b[40])^(a[36] & b[41])^(a[35] & b[42])^(a[34] & b[43])^(a[33] & b[44])^(a[32] & b[45])^(a[31] & b[46])^(a[30] & b[47])^(a[29] & b[48])^(a[28] & b[49])^(a[27] & b[50])^(a[26] & b[51])^(a[25] & b[52])^(a[24] & b[53])^(a[23] & b[54])^(a[22] & b[55])^(a[21] & b[56])^(a[20] & b[57])^(a[19] & b[58])^(a[18] & b[59])^(a[17] & b[60])^(a[16] & b[61])^(a[15] & b[62])^(a[14] & b[63])^(a[13] & b[64])^(a[12] & b[65])^(a[11] & b[66])^(a[10] & b[67])^(a[9] & b[68])^(a[8] & b[69])^(a[7] & b[70])^(a[6] & b[71])^(a[5] & b[72])^(a[4] & b[73])^(a[3] & b[74])^(a[2] & b[75])^(a[1] & b[76])^(a[0] & b[77]);
assign y[78] = (a[78] & b[0])^(a[77] & b[1])^(a[76] & b[2])^(a[75] & b[3])^(a[74] & b[4])^(a[73] & b[5])^(a[72] & b[6])^(a[71] & b[7])^(a[70] & b[8])^(a[69] & b[9])^(a[68] & b[10])^(a[67] & b[11])^(a[66] & b[12])^(a[65] & b[13])^(a[64] & b[14])^(a[63] & b[15])^(a[62] & b[16])^(a[61] & b[17])^(a[60] & b[18])^(a[59] & b[19])^(a[58] & b[20])^(a[57] & b[21])^(a[56] & b[22])^(a[55] & b[23])^(a[54] & b[24])^(a[53] & b[25])^(a[52] & b[26])^(a[51] & b[27])^(a[50] & b[28])^(a[49] & b[29])^(a[48] & b[30])^(a[47] & b[31])^(a[46] & b[32])^(a[45] & b[33])^(a[44] & b[34])^(a[43] & b[35])^(a[42] & b[36])^(a[41] & b[37])^(a[40] & b[38])^(a[39] & b[39])^(a[38] & b[40])^(a[37] & b[41])^(a[36] & b[42])^(a[35] & b[43])^(a[34] & b[44])^(a[33] & b[45])^(a[32] & b[46])^(a[31] & b[47])^(a[30] & b[48])^(a[29] & b[49])^(a[28] & b[50])^(a[27] & b[51])^(a[26] & b[52])^(a[25] & b[53])^(a[24] & b[54])^(a[23] & b[55])^(a[22] & b[56])^(a[21] & b[57])^(a[20] & b[58])^(a[19] & b[59])^(a[18] & b[60])^(a[17] & b[61])^(a[16] & b[62])^(a[15] & b[63])^(a[14] & b[64])^(a[13] & b[65])^(a[12] & b[66])^(a[11] & b[67])^(a[10] & b[68])^(a[9] & b[69])^(a[8] & b[70])^(a[7] & b[71])^(a[6] & b[72])^(a[5] & b[73])^(a[4] & b[74])^(a[3] & b[75])^(a[2] & b[76])^(a[1] & b[77])^(a[0] & b[78]);
assign y[79] = (a[79] & b[0])^(a[78] & b[1])^(a[77] & b[2])^(a[76] & b[3])^(a[75] & b[4])^(a[74] & b[5])^(a[73] & b[6])^(a[72] & b[7])^(a[71] & b[8])^(a[70] & b[9])^(a[69] & b[10])^(a[68] & b[11])^(a[67] & b[12])^(a[66] & b[13])^(a[65] & b[14])^(a[64] & b[15])^(a[63] & b[16])^(a[62] & b[17])^(a[61] & b[18])^(a[60] & b[19])^(a[59] & b[20])^(a[58] & b[21])^(a[57] & b[22])^(a[56] & b[23])^(a[55] & b[24])^(a[54] & b[25])^(a[53] & b[26])^(a[52] & b[27])^(a[51] & b[28])^(a[50] & b[29])^(a[49] & b[30])^(a[48] & b[31])^(a[47] & b[32])^(a[46] & b[33])^(a[45] & b[34])^(a[44] & b[35])^(a[43] & b[36])^(a[42] & b[37])^(a[41] & b[38])^(a[40] & b[39])^(a[39] & b[40])^(a[38] & b[41])^(a[37] & b[42])^(a[36] & b[43])^(a[35] & b[44])^(a[34] & b[45])^(a[33] & b[46])^(a[32] & b[47])^(a[31] & b[48])^(a[30] & b[49])^(a[29] & b[50])^(a[28] & b[51])^(a[27] & b[52])^(a[26] & b[53])^(a[25] & b[54])^(a[24] & b[55])^(a[23] & b[56])^(a[22] & b[57])^(a[21] & b[58])^(a[20] & b[59])^(a[19] & b[60])^(a[18] & b[61])^(a[17] & b[62])^(a[16] & b[63])^(a[15] & b[64])^(a[14] & b[65])^(a[13] & b[66])^(a[12] & b[67])^(a[11] & b[68])^(a[10] & b[69])^(a[9] & b[70])^(a[8] & b[71])^(a[7] & b[72])^(a[6] & b[73])^(a[5] & b[74])^(a[4] & b[75])^(a[3] & b[76])^(a[2] & b[77])^(a[1] & b[78])^(a[0] & b[79]);
assign y[80] = (a[80] & b[0])^(a[79] & b[1])^(a[78] & b[2])^(a[77] & b[3])^(a[76] & b[4])^(a[75] & b[5])^(a[74] & b[6])^(a[73] & b[7])^(a[72] & b[8])^(a[71] & b[9])^(a[70] & b[10])^(a[69] & b[11])^(a[68] & b[12])^(a[67] & b[13])^(a[66] & b[14])^(a[65] & b[15])^(a[64] & b[16])^(a[63] & b[17])^(a[62] & b[18])^(a[61] & b[19])^(a[60] & b[20])^(a[59] & b[21])^(a[58] & b[22])^(a[57] & b[23])^(a[56] & b[24])^(a[55] & b[25])^(a[54] & b[26])^(a[53] & b[27])^(a[52] & b[28])^(a[51] & b[29])^(a[50] & b[30])^(a[49] & b[31])^(a[48] & b[32])^(a[47] & b[33])^(a[46] & b[34])^(a[45] & b[35])^(a[44] & b[36])^(a[43] & b[37])^(a[42] & b[38])^(a[41] & b[39])^(a[40] & b[40])^(a[39] & b[41])^(a[38] & b[42])^(a[37] & b[43])^(a[36] & b[44])^(a[35] & b[45])^(a[34] & b[46])^(a[33] & b[47])^(a[32] & b[48])^(a[31] & b[49])^(a[30] & b[50])^(a[29] & b[51])^(a[28] & b[52])^(a[27] & b[53])^(a[26] & b[54])^(a[25] & b[55])^(a[24] & b[56])^(a[23] & b[57])^(a[22] & b[58])^(a[21] & b[59])^(a[20] & b[60])^(a[19] & b[61])^(a[18] & b[62])^(a[17] & b[63])^(a[16] & b[64])^(a[15] & b[65])^(a[14] & b[66])^(a[13] & b[67])^(a[12] & b[68])^(a[11] & b[69])^(a[10] & b[70])^(a[9] & b[71])^(a[8] & b[72])^(a[7] & b[73])^(a[6] & b[74])^(a[5] & b[75])^(a[4] & b[76])^(a[3] & b[77])^(a[2] & b[78])^(a[1] & b[79])^(a[0] & b[80]);
assign y[81] = (a[81] & b[0])^(a[80] & b[1])^(a[79] & b[2])^(a[78] & b[3])^(a[77] & b[4])^(a[76] & b[5])^(a[75] & b[6])^(a[74] & b[7])^(a[73] & b[8])^(a[72] & b[9])^(a[71] & b[10])^(a[70] & b[11])^(a[69] & b[12])^(a[68] & b[13])^(a[67] & b[14])^(a[66] & b[15])^(a[65] & b[16])^(a[64] & b[17])^(a[63] & b[18])^(a[62] & b[19])^(a[61] & b[20])^(a[60] & b[21])^(a[59] & b[22])^(a[58] & b[23])^(a[57] & b[24])^(a[56] & b[25])^(a[55] & b[26])^(a[54] & b[27])^(a[53] & b[28])^(a[52] & b[29])^(a[51] & b[30])^(a[50] & b[31])^(a[49] & b[32])^(a[48] & b[33])^(a[47] & b[34])^(a[46] & b[35])^(a[45] & b[36])^(a[44] & b[37])^(a[43] & b[38])^(a[42] & b[39])^(a[41] & b[40])^(a[40] & b[41])^(a[39] & b[42])^(a[38] & b[43])^(a[37] & b[44])^(a[36] & b[45])^(a[35] & b[46])^(a[34] & b[47])^(a[33] & b[48])^(a[32] & b[49])^(a[31] & b[50])^(a[30] & b[51])^(a[29] & b[52])^(a[28] & b[53])^(a[27] & b[54])^(a[26] & b[55])^(a[25] & b[56])^(a[24] & b[57])^(a[23] & b[58])^(a[22] & b[59])^(a[21] & b[60])^(a[20] & b[61])^(a[19] & b[62])^(a[18] & b[63])^(a[17] & b[64])^(a[16] & b[65])^(a[15] & b[66])^(a[14] & b[67])^(a[13] & b[68])^(a[12] & b[69])^(a[11] & b[70])^(a[10] & b[71])^(a[9] & b[72])^(a[8] & b[73])^(a[7] & b[74])^(a[6] & b[75])^(a[5] & b[76])^(a[4] & b[77])^(a[3] & b[78])^(a[2] & b[79])^(a[1] & b[80])^(a[0] & b[81]);
assign y[82] = (a[82] & b[0])^(a[81] & b[1])^(a[80] & b[2])^(a[79] & b[3])^(a[78] & b[4])^(a[77] & b[5])^(a[76] & b[6])^(a[75] & b[7])^(a[74] & b[8])^(a[73] & b[9])^(a[72] & b[10])^(a[71] & b[11])^(a[70] & b[12])^(a[69] & b[13])^(a[68] & b[14])^(a[67] & b[15])^(a[66] & b[16])^(a[65] & b[17])^(a[64] & b[18])^(a[63] & b[19])^(a[62] & b[20])^(a[61] & b[21])^(a[60] & b[22])^(a[59] & b[23])^(a[58] & b[24])^(a[57] & b[25])^(a[56] & b[26])^(a[55] & b[27])^(a[54] & b[28])^(a[53] & b[29])^(a[52] & b[30])^(a[51] & b[31])^(a[50] & b[32])^(a[49] & b[33])^(a[48] & b[34])^(a[47] & b[35])^(a[46] & b[36])^(a[45] & b[37])^(a[44] & b[38])^(a[43] & b[39])^(a[42] & b[40])^(a[41] & b[41])^(a[40] & b[42])^(a[39] & b[43])^(a[38] & b[44])^(a[37] & b[45])^(a[36] & b[46])^(a[35] & b[47])^(a[34] & b[48])^(a[33] & b[49])^(a[32] & b[50])^(a[31] & b[51])^(a[30] & b[52])^(a[29] & b[53])^(a[28] & b[54])^(a[27] & b[55])^(a[26] & b[56])^(a[25] & b[57])^(a[24] & b[58])^(a[23] & b[59])^(a[22] & b[60])^(a[21] & b[61])^(a[20] & b[62])^(a[19] & b[63])^(a[18] & b[64])^(a[17] & b[65])^(a[16] & b[66])^(a[15] & b[67])^(a[14] & b[68])^(a[13] & b[69])^(a[12] & b[70])^(a[11] & b[71])^(a[10] & b[72])^(a[9] & b[73])^(a[8] & b[74])^(a[7] & b[75])^(a[6] & b[76])^(a[5] & b[77])^(a[4] & b[78])^(a[3] & b[79])^(a[2] & b[80])^(a[1] & b[81])^(a[0] & b[82]);
assign y[83] = (a[83] & b[0])^(a[82] & b[1])^(a[81] & b[2])^(a[80] & b[3])^(a[79] & b[4])^(a[78] & b[5])^(a[77] & b[6])^(a[76] & b[7])^(a[75] & b[8])^(a[74] & b[9])^(a[73] & b[10])^(a[72] & b[11])^(a[71] & b[12])^(a[70] & b[13])^(a[69] & b[14])^(a[68] & b[15])^(a[67] & b[16])^(a[66] & b[17])^(a[65] & b[18])^(a[64] & b[19])^(a[63] & b[20])^(a[62] & b[21])^(a[61] & b[22])^(a[60] & b[23])^(a[59] & b[24])^(a[58] & b[25])^(a[57] & b[26])^(a[56] & b[27])^(a[55] & b[28])^(a[54] & b[29])^(a[53] & b[30])^(a[52] & b[31])^(a[51] & b[32])^(a[50] & b[33])^(a[49] & b[34])^(a[48] & b[35])^(a[47] & b[36])^(a[46] & b[37])^(a[45] & b[38])^(a[44] & b[39])^(a[43] & b[40])^(a[42] & b[41])^(a[41] & b[42])^(a[40] & b[43])^(a[39] & b[44])^(a[38] & b[45])^(a[37] & b[46])^(a[36] & b[47])^(a[35] & b[48])^(a[34] & b[49])^(a[33] & b[50])^(a[32] & b[51])^(a[31] & b[52])^(a[30] & b[53])^(a[29] & b[54])^(a[28] & b[55])^(a[27] & b[56])^(a[26] & b[57])^(a[25] & b[58])^(a[24] & b[59])^(a[23] & b[60])^(a[22] & b[61])^(a[21] & b[62])^(a[20] & b[63])^(a[19] & b[64])^(a[18] & b[65])^(a[17] & b[66])^(a[16] & b[67])^(a[15] & b[68])^(a[14] & b[69])^(a[13] & b[70])^(a[12] & b[71])^(a[11] & b[72])^(a[10] & b[73])^(a[9] & b[74])^(a[8] & b[75])^(a[7] & b[76])^(a[6] & b[77])^(a[5] & b[78])^(a[4] & b[79])^(a[3] & b[80])^(a[2] & b[81])^(a[1] & b[82])^(a[0] & b[83]);
assign y[84] = (a[84] & b[0])^(a[83] & b[1])^(a[82] & b[2])^(a[81] & b[3])^(a[80] & b[4])^(a[79] & b[5])^(a[78] & b[6])^(a[77] & b[7])^(a[76] & b[8])^(a[75] & b[9])^(a[74] & b[10])^(a[73] & b[11])^(a[72] & b[12])^(a[71] & b[13])^(a[70] & b[14])^(a[69] & b[15])^(a[68] & b[16])^(a[67] & b[17])^(a[66] & b[18])^(a[65] & b[19])^(a[64] & b[20])^(a[63] & b[21])^(a[62] & b[22])^(a[61] & b[23])^(a[60] & b[24])^(a[59] & b[25])^(a[58] & b[26])^(a[57] & b[27])^(a[56] & b[28])^(a[55] & b[29])^(a[54] & b[30])^(a[53] & b[31])^(a[52] & b[32])^(a[51] & b[33])^(a[50] & b[34])^(a[49] & b[35])^(a[48] & b[36])^(a[47] & b[37])^(a[46] & b[38])^(a[45] & b[39])^(a[44] & b[40])^(a[43] & b[41])^(a[42] & b[42])^(a[41] & b[43])^(a[40] & b[44])^(a[39] & b[45])^(a[38] & b[46])^(a[37] & b[47])^(a[36] & b[48])^(a[35] & b[49])^(a[34] & b[50])^(a[33] & b[51])^(a[32] & b[52])^(a[31] & b[53])^(a[30] & b[54])^(a[29] & b[55])^(a[28] & b[56])^(a[27] & b[57])^(a[26] & b[58])^(a[25] & b[59])^(a[24] & b[60])^(a[23] & b[61])^(a[22] & b[62])^(a[21] & b[63])^(a[20] & b[64])^(a[19] & b[65])^(a[18] & b[66])^(a[17] & b[67])^(a[16] & b[68])^(a[15] & b[69])^(a[14] & b[70])^(a[13] & b[71])^(a[12] & b[72])^(a[11] & b[73])^(a[10] & b[74])^(a[9] & b[75])^(a[8] & b[76])^(a[7] & b[77])^(a[6] & b[78])^(a[5] & b[79])^(a[4] & b[80])^(a[3] & b[81])^(a[2] & b[82])^(a[1] & b[83])^(a[0] & b[84]);
assign y[85] = (a[85] & b[0])^(a[84] & b[1])^(a[83] & b[2])^(a[82] & b[3])^(a[81] & b[4])^(a[80] & b[5])^(a[79] & b[6])^(a[78] & b[7])^(a[77] & b[8])^(a[76] & b[9])^(a[75] & b[10])^(a[74] & b[11])^(a[73] & b[12])^(a[72] & b[13])^(a[71] & b[14])^(a[70] & b[15])^(a[69] & b[16])^(a[68] & b[17])^(a[67] & b[18])^(a[66] & b[19])^(a[65] & b[20])^(a[64] & b[21])^(a[63] & b[22])^(a[62] & b[23])^(a[61] & b[24])^(a[60] & b[25])^(a[59] & b[26])^(a[58] & b[27])^(a[57] & b[28])^(a[56] & b[29])^(a[55] & b[30])^(a[54] & b[31])^(a[53] & b[32])^(a[52] & b[33])^(a[51] & b[34])^(a[50] & b[35])^(a[49] & b[36])^(a[48] & b[37])^(a[47] & b[38])^(a[46] & b[39])^(a[45] & b[40])^(a[44] & b[41])^(a[43] & b[42])^(a[42] & b[43])^(a[41] & b[44])^(a[40] & b[45])^(a[39] & b[46])^(a[38] & b[47])^(a[37] & b[48])^(a[36] & b[49])^(a[35] & b[50])^(a[34] & b[51])^(a[33] & b[52])^(a[32] & b[53])^(a[31] & b[54])^(a[30] & b[55])^(a[29] & b[56])^(a[28] & b[57])^(a[27] & b[58])^(a[26] & b[59])^(a[25] & b[60])^(a[24] & b[61])^(a[23] & b[62])^(a[22] & b[63])^(a[21] & b[64])^(a[20] & b[65])^(a[19] & b[66])^(a[18] & b[67])^(a[17] & b[68])^(a[16] & b[69])^(a[15] & b[70])^(a[14] & b[71])^(a[13] & b[72])^(a[12] & b[73])^(a[11] & b[74])^(a[10] & b[75])^(a[9] & b[76])^(a[8] & b[77])^(a[7] & b[78])^(a[6] & b[79])^(a[5] & b[80])^(a[4] & b[81])^(a[3] & b[82])^(a[2] & b[83])^(a[1] & b[84])^(a[0] & b[85]);
assign y[86] = (a[86] & b[0])^(a[85] & b[1])^(a[84] & b[2])^(a[83] & b[3])^(a[82] & b[4])^(a[81] & b[5])^(a[80] & b[6])^(a[79] & b[7])^(a[78] & b[8])^(a[77] & b[9])^(a[76] & b[10])^(a[75] & b[11])^(a[74] & b[12])^(a[73] & b[13])^(a[72] & b[14])^(a[71] & b[15])^(a[70] & b[16])^(a[69] & b[17])^(a[68] & b[18])^(a[67] & b[19])^(a[66] & b[20])^(a[65] & b[21])^(a[64] & b[22])^(a[63] & b[23])^(a[62] & b[24])^(a[61] & b[25])^(a[60] & b[26])^(a[59] & b[27])^(a[58] & b[28])^(a[57] & b[29])^(a[56] & b[30])^(a[55] & b[31])^(a[54] & b[32])^(a[53] & b[33])^(a[52] & b[34])^(a[51] & b[35])^(a[50] & b[36])^(a[49] & b[37])^(a[48] & b[38])^(a[47] & b[39])^(a[46] & b[40])^(a[45] & b[41])^(a[44] & b[42])^(a[43] & b[43])^(a[42] & b[44])^(a[41] & b[45])^(a[40] & b[46])^(a[39] & b[47])^(a[38] & b[48])^(a[37] & b[49])^(a[36] & b[50])^(a[35] & b[51])^(a[34] & b[52])^(a[33] & b[53])^(a[32] & b[54])^(a[31] & b[55])^(a[30] & b[56])^(a[29] & b[57])^(a[28] & b[58])^(a[27] & b[59])^(a[26] & b[60])^(a[25] & b[61])^(a[24] & b[62])^(a[23] & b[63])^(a[22] & b[64])^(a[21] & b[65])^(a[20] & b[66])^(a[19] & b[67])^(a[18] & b[68])^(a[17] & b[69])^(a[16] & b[70])^(a[15] & b[71])^(a[14] & b[72])^(a[13] & b[73])^(a[12] & b[74])^(a[11] & b[75])^(a[10] & b[76])^(a[9] & b[77])^(a[8] & b[78])^(a[7] & b[79])^(a[6] & b[80])^(a[5] & b[81])^(a[4] & b[82])^(a[3] & b[83])^(a[2] & b[84])^(a[1] & b[85])^(a[0] & b[86]);
assign y[87] = (a[87] & b[0])^(a[86] & b[1])^(a[85] & b[2])^(a[84] & b[3])^(a[83] & b[4])^(a[82] & b[5])^(a[81] & b[6])^(a[80] & b[7])^(a[79] & b[8])^(a[78] & b[9])^(a[77] & b[10])^(a[76] & b[11])^(a[75] & b[12])^(a[74] & b[13])^(a[73] & b[14])^(a[72] & b[15])^(a[71] & b[16])^(a[70] & b[17])^(a[69] & b[18])^(a[68] & b[19])^(a[67] & b[20])^(a[66] & b[21])^(a[65] & b[22])^(a[64] & b[23])^(a[63] & b[24])^(a[62] & b[25])^(a[61] & b[26])^(a[60] & b[27])^(a[59] & b[28])^(a[58] & b[29])^(a[57] & b[30])^(a[56] & b[31])^(a[55] & b[32])^(a[54] & b[33])^(a[53] & b[34])^(a[52] & b[35])^(a[51] & b[36])^(a[50] & b[37])^(a[49] & b[38])^(a[48] & b[39])^(a[47] & b[40])^(a[46] & b[41])^(a[45] & b[42])^(a[44] & b[43])^(a[43] & b[44])^(a[42] & b[45])^(a[41] & b[46])^(a[40] & b[47])^(a[39] & b[48])^(a[38] & b[49])^(a[37] & b[50])^(a[36] & b[51])^(a[35] & b[52])^(a[34] & b[53])^(a[33] & b[54])^(a[32] & b[55])^(a[31] & b[56])^(a[30] & b[57])^(a[29] & b[58])^(a[28] & b[59])^(a[27] & b[60])^(a[26] & b[61])^(a[25] & b[62])^(a[24] & b[63])^(a[23] & b[64])^(a[22] & b[65])^(a[21] & b[66])^(a[20] & b[67])^(a[19] & b[68])^(a[18] & b[69])^(a[17] & b[70])^(a[16] & b[71])^(a[15] & b[72])^(a[14] & b[73])^(a[13] & b[74])^(a[12] & b[75])^(a[11] & b[76])^(a[10] & b[77])^(a[9] & b[78])^(a[8] & b[79])^(a[7] & b[80])^(a[6] & b[81])^(a[5] & b[82])^(a[4] & b[83])^(a[3] & b[84])^(a[2] & b[85])^(a[1] & b[86])^(a[0] & b[87]);
assign y[88] = (a[88] & b[0])^(a[87] & b[1])^(a[86] & b[2])^(a[85] & b[3])^(a[84] & b[4])^(a[83] & b[5])^(a[82] & b[6])^(a[81] & b[7])^(a[80] & b[8])^(a[79] & b[9])^(a[78] & b[10])^(a[77] & b[11])^(a[76] & b[12])^(a[75] & b[13])^(a[74] & b[14])^(a[73] & b[15])^(a[72] & b[16])^(a[71] & b[17])^(a[70] & b[18])^(a[69] & b[19])^(a[68] & b[20])^(a[67] & b[21])^(a[66] & b[22])^(a[65] & b[23])^(a[64] & b[24])^(a[63] & b[25])^(a[62] & b[26])^(a[61] & b[27])^(a[60] & b[28])^(a[59] & b[29])^(a[58] & b[30])^(a[57] & b[31])^(a[56] & b[32])^(a[55] & b[33])^(a[54] & b[34])^(a[53] & b[35])^(a[52] & b[36])^(a[51] & b[37])^(a[50] & b[38])^(a[49] & b[39])^(a[48] & b[40])^(a[47] & b[41])^(a[46] & b[42])^(a[45] & b[43])^(a[44] & b[44])^(a[43] & b[45])^(a[42] & b[46])^(a[41] & b[47])^(a[40] & b[48])^(a[39] & b[49])^(a[38] & b[50])^(a[37] & b[51])^(a[36] & b[52])^(a[35] & b[53])^(a[34] & b[54])^(a[33] & b[55])^(a[32] & b[56])^(a[31] & b[57])^(a[30] & b[58])^(a[29] & b[59])^(a[28] & b[60])^(a[27] & b[61])^(a[26] & b[62])^(a[25] & b[63])^(a[24] & b[64])^(a[23] & b[65])^(a[22] & b[66])^(a[21] & b[67])^(a[20] & b[68])^(a[19] & b[69])^(a[18] & b[70])^(a[17] & b[71])^(a[16] & b[72])^(a[15] & b[73])^(a[14] & b[74])^(a[13] & b[75])^(a[12] & b[76])^(a[11] & b[77])^(a[10] & b[78])^(a[9] & b[79])^(a[8] & b[80])^(a[7] & b[81])^(a[6] & b[82])^(a[5] & b[83])^(a[4] & b[84])^(a[3] & b[85])^(a[2] & b[86])^(a[1] & b[87])^(a[0] & b[88]);
assign y[89] = (a[89] & b[0])^(a[88] & b[1])^(a[87] & b[2])^(a[86] & b[3])^(a[85] & b[4])^(a[84] & b[5])^(a[83] & b[6])^(a[82] & b[7])^(a[81] & b[8])^(a[80] & b[9])^(a[79] & b[10])^(a[78] & b[11])^(a[77] & b[12])^(a[76] & b[13])^(a[75] & b[14])^(a[74] & b[15])^(a[73] & b[16])^(a[72] & b[17])^(a[71] & b[18])^(a[70] & b[19])^(a[69] & b[20])^(a[68] & b[21])^(a[67] & b[22])^(a[66] & b[23])^(a[65] & b[24])^(a[64] & b[25])^(a[63] & b[26])^(a[62] & b[27])^(a[61] & b[28])^(a[60] & b[29])^(a[59] & b[30])^(a[58] & b[31])^(a[57] & b[32])^(a[56] & b[33])^(a[55] & b[34])^(a[54] & b[35])^(a[53] & b[36])^(a[52] & b[37])^(a[51] & b[38])^(a[50] & b[39])^(a[49] & b[40])^(a[48] & b[41])^(a[47] & b[42])^(a[46] & b[43])^(a[45] & b[44])^(a[44] & b[45])^(a[43] & b[46])^(a[42] & b[47])^(a[41] & b[48])^(a[40] & b[49])^(a[39] & b[50])^(a[38] & b[51])^(a[37] & b[52])^(a[36] & b[53])^(a[35] & b[54])^(a[34] & b[55])^(a[33] & b[56])^(a[32] & b[57])^(a[31] & b[58])^(a[30] & b[59])^(a[29] & b[60])^(a[28] & b[61])^(a[27] & b[62])^(a[26] & b[63])^(a[25] & b[64])^(a[24] & b[65])^(a[23] & b[66])^(a[22] & b[67])^(a[21] & b[68])^(a[20] & b[69])^(a[19] & b[70])^(a[18] & b[71])^(a[17] & b[72])^(a[16] & b[73])^(a[15] & b[74])^(a[14] & b[75])^(a[13] & b[76])^(a[12] & b[77])^(a[11] & b[78])^(a[10] & b[79])^(a[9] & b[80])^(a[8] & b[81])^(a[7] & b[82])^(a[6] & b[83])^(a[5] & b[84])^(a[4] & b[85])^(a[3] & b[86])^(a[2] & b[87])^(a[1] & b[88])^(a[0] & b[89]);
assign y[90] = (a[90] & b[0])^(a[89] & b[1])^(a[88] & b[2])^(a[87] & b[3])^(a[86] & b[4])^(a[85] & b[5])^(a[84] & b[6])^(a[83] & b[7])^(a[82] & b[8])^(a[81] & b[9])^(a[80] & b[10])^(a[79] & b[11])^(a[78] & b[12])^(a[77] & b[13])^(a[76] & b[14])^(a[75] & b[15])^(a[74] & b[16])^(a[73] & b[17])^(a[72] & b[18])^(a[71] & b[19])^(a[70] & b[20])^(a[69] & b[21])^(a[68] & b[22])^(a[67] & b[23])^(a[66] & b[24])^(a[65] & b[25])^(a[64] & b[26])^(a[63] & b[27])^(a[62] & b[28])^(a[61] & b[29])^(a[60] & b[30])^(a[59] & b[31])^(a[58] & b[32])^(a[57] & b[33])^(a[56] & b[34])^(a[55] & b[35])^(a[54] & b[36])^(a[53] & b[37])^(a[52] & b[38])^(a[51] & b[39])^(a[50] & b[40])^(a[49] & b[41])^(a[48] & b[42])^(a[47] & b[43])^(a[46] & b[44])^(a[45] & b[45])^(a[44] & b[46])^(a[43] & b[47])^(a[42] & b[48])^(a[41] & b[49])^(a[40] & b[50])^(a[39] & b[51])^(a[38] & b[52])^(a[37] & b[53])^(a[36] & b[54])^(a[35] & b[55])^(a[34] & b[56])^(a[33] & b[57])^(a[32] & b[58])^(a[31] & b[59])^(a[30] & b[60])^(a[29] & b[61])^(a[28] & b[62])^(a[27] & b[63])^(a[26] & b[64])^(a[25] & b[65])^(a[24] & b[66])^(a[23] & b[67])^(a[22] & b[68])^(a[21] & b[69])^(a[20] & b[70])^(a[19] & b[71])^(a[18] & b[72])^(a[17] & b[73])^(a[16] & b[74])^(a[15] & b[75])^(a[14] & b[76])^(a[13] & b[77])^(a[12] & b[78])^(a[11] & b[79])^(a[10] & b[80])^(a[9] & b[81])^(a[8] & b[82])^(a[7] & b[83])^(a[6] & b[84])^(a[5] & b[85])^(a[4] & b[86])^(a[3] & b[87])^(a[2] & b[88])^(a[1] & b[89])^(a[0] & b[90]);
assign y[91] = (a[91] & b[0])^(a[90] & b[1])^(a[89] & b[2])^(a[88] & b[3])^(a[87] & b[4])^(a[86] & b[5])^(a[85] & b[6])^(a[84] & b[7])^(a[83] & b[8])^(a[82] & b[9])^(a[81] & b[10])^(a[80] & b[11])^(a[79] & b[12])^(a[78] & b[13])^(a[77] & b[14])^(a[76] & b[15])^(a[75] & b[16])^(a[74] & b[17])^(a[73] & b[18])^(a[72] & b[19])^(a[71] & b[20])^(a[70] & b[21])^(a[69] & b[22])^(a[68] & b[23])^(a[67] & b[24])^(a[66] & b[25])^(a[65] & b[26])^(a[64] & b[27])^(a[63] & b[28])^(a[62] & b[29])^(a[61] & b[30])^(a[60] & b[31])^(a[59] & b[32])^(a[58] & b[33])^(a[57] & b[34])^(a[56] & b[35])^(a[55] & b[36])^(a[54] & b[37])^(a[53] & b[38])^(a[52] & b[39])^(a[51] & b[40])^(a[50] & b[41])^(a[49] & b[42])^(a[48] & b[43])^(a[47] & b[44])^(a[46] & b[45])^(a[45] & b[46])^(a[44] & b[47])^(a[43] & b[48])^(a[42] & b[49])^(a[41] & b[50])^(a[40] & b[51])^(a[39] & b[52])^(a[38] & b[53])^(a[37] & b[54])^(a[36] & b[55])^(a[35] & b[56])^(a[34] & b[57])^(a[33] & b[58])^(a[32] & b[59])^(a[31] & b[60])^(a[30] & b[61])^(a[29] & b[62])^(a[28] & b[63])^(a[27] & b[64])^(a[26] & b[65])^(a[25] & b[66])^(a[24] & b[67])^(a[23] & b[68])^(a[22] & b[69])^(a[21] & b[70])^(a[20] & b[71])^(a[19] & b[72])^(a[18] & b[73])^(a[17] & b[74])^(a[16] & b[75])^(a[15] & b[76])^(a[14] & b[77])^(a[13] & b[78])^(a[12] & b[79])^(a[11] & b[80])^(a[10] & b[81])^(a[9] & b[82])^(a[8] & b[83])^(a[7] & b[84])^(a[6] & b[85])^(a[5] & b[86])^(a[4] & b[87])^(a[3] & b[88])^(a[2] & b[89])^(a[1] & b[90])^(a[0] & b[91]);
assign y[92] = (a[92] & b[0])^(a[91] & b[1])^(a[90] & b[2])^(a[89] & b[3])^(a[88] & b[4])^(a[87] & b[5])^(a[86] & b[6])^(a[85] & b[7])^(a[84] & b[8])^(a[83] & b[9])^(a[82] & b[10])^(a[81] & b[11])^(a[80] & b[12])^(a[79] & b[13])^(a[78] & b[14])^(a[77] & b[15])^(a[76] & b[16])^(a[75] & b[17])^(a[74] & b[18])^(a[73] & b[19])^(a[72] & b[20])^(a[71] & b[21])^(a[70] & b[22])^(a[69] & b[23])^(a[68] & b[24])^(a[67] & b[25])^(a[66] & b[26])^(a[65] & b[27])^(a[64] & b[28])^(a[63] & b[29])^(a[62] & b[30])^(a[61] & b[31])^(a[60] & b[32])^(a[59] & b[33])^(a[58] & b[34])^(a[57] & b[35])^(a[56] & b[36])^(a[55] & b[37])^(a[54] & b[38])^(a[53] & b[39])^(a[52] & b[40])^(a[51] & b[41])^(a[50] & b[42])^(a[49] & b[43])^(a[48] & b[44])^(a[47] & b[45])^(a[46] & b[46])^(a[45] & b[47])^(a[44] & b[48])^(a[43] & b[49])^(a[42] & b[50])^(a[41] & b[51])^(a[40] & b[52])^(a[39] & b[53])^(a[38] & b[54])^(a[37] & b[55])^(a[36] & b[56])^(a[35] & b[57])^(a[34] & b[58])^(a[33] & b[59])^(a[32] & b[60])^(a[31] & b[61])^(a[30] & b[62])^(a[29] & b[63])^(a[28] & b[64])^(a[27] & b[65])^(a[26] & b[66])^(a[25] & b[67])^(a[24] & b[68])^(a[23] & b[69])^(a[22] & b[70])^(a[21] & b[71])^(a[20] & b[72])^(a[19] & b[73])^(a[18] & b[74])^(a[17] & b[75])^(a[16] & b[76])^(a[15] & b[77])^(a[14] & b[78])^(a[13] & b[79])^(a[12] & b[80])^(a[11] & b[81])^(a[10] & b[82])^(a[9] & b[83])^(a[8] & b[84])^(a[7] & b[85])^(a[6] & b[86])^(a[5] & b[87])^(a[4] & b[88])^(a[3] & b[89])^(a[2] & b[90])^(a[1] & b[91])^(a[0] & b[92]);
assign y[93] = (a[93] & b[0])^(a[92] & b[1])^(a[91] & b[2])^(a[90] & b[3])^(a[89] & b[4])^(a[88] & b[5])^(a[87] & b[6])^(a[86] & b[7])^(a[85] & b[8])^(a[84] & b[9])^(a[83] & b[10])^(a[82] & b[11])^(a[81] & b[12])^(a[80] & b[13])^(a[79] & b[14])^(a[78] & b[15])^(a[77] & b[16])^(a[76] & b[17])^(a[75] & b[18])^(a[74] & b[19])^(a[73] & b[20])^(a[72] & b[21])^(a[71] & b[22])^(a[70] & b[23])^(a[69] & b[24])^(a[68] & b[25])^(a[67] & b[26])^(a[66] & b[27])^(a[65] & b[28])^(a[64] & b[29])^(a[63] & b[30])^(a[62] & b[31])^(a[61] & b[32])^(a[60] & b[33])^(a[59] & b[34])^(a[58] & b[35])^(a[57] & b[36])^(a[56] & b[37])^(a[55] & b[38])^(a[54] & b[39])^(a[53] & b[40])^(a[52] & b[41])^(a[51] & b[42])^(a[50] & b[43])^(a[49] & b[44])^(a[48] & b[45])^(a[47] & b[46])^(a[46] & b[47])^(a[45] & b[48])^(a[44] & b[49])^(a[43] & b[50])^(a[42] & b[51])^(a[41] & b[52])^(a[40] & b[53])^(a[39] & b[54])^(a[38] & b[55])^(a[37] & b[56])^(a[36] & b[57])^(a[35] & b[58])^(a[34] & b[59])^(a[33] & b[60])^(a[32] & b[61])^(a[31] & b[62])^(a[30] & b[63])^(a[29] & b[64])^(a[28] & b[65])^(a[27] & b[66])^(a[26] & b[67])^(a[25] & b[68])^(a[24] & b[69])^(a[23] & b[70])^(a[22] & b[71])^(a[21] & b[72])^(a[20] & b[73])^(a[19] & b[74])^(a[18] & b[75])^(a[17] & b[76])^(a[16] & b[77])^(a[15] & b[78])^(a[14] & b[79])^(a[13] & b[80])^(a[12] & b[81])^(a[11] & b[82])^(a[10] & b[83])^(a[9] & b[84])^(a[8] & b[85])^(a[7] & b[86])^(a[6] & b[87])^(a[5] & b[88])^(a[4] & b[89])^(a[3] & b[90])^(a[2] & b[91])^(a[1] & b[92])^(a[0] & b[93]);
assign y[94] = (a[94] & b[0])^(a[93] & b[1])^(a[92] & b[2])^(a[91] & b[3])^(a[90] & b[4])^(a[89] & b[5])^(a[88] & b[6])^(a[87] & b[7])^(a[86] & b[8])^(a[85] & b[9])^(a[84] & b[10])^(a[83] & b[11])^(a[82] & b[12])^(a[81] & b[13])^(a[80] & b[14])^(a[79] & b[15])^(a[78] & b[16])^(a[77] & b[17])^(a[76] & b[18])^(a[75] & b[19])^(a[74] & b[20])^(a[73] & b[21])^(a[72] & b[22])^(a[71] & b[23])^(a[70] & b[24])^(a[69] & b[25])^(a[68] & b[26])^(a[67] & b[27])^(a[66] & b[28])^(a[65] & b[29])^(a[64] & b[30])^(a[63] & b[31])^(a[62] & b[32])^(a[61] & b[33])^(a[60] & b[34])^(a[59] & b[35])^(a[58] & b[36])^(a[57] & b[37])^(a[56] & b[38])^(a[55] & b[39])^(a[54] & b[40])^(a[53] & b[41])^(a[52] & b[42])^(a[51] & b[43])^(a[50] & b[44])^(a[49] & b[45])^(a[48] & b[46])^(a[47] & b[47])^(a[46] & b[48])^(a[45] & b[49])^(a[44] & b[50])^(a[43] & b[51])^(a[42] & b[52])^(a[41] & b[53])^(a[40] & b[54])^(a[39] & b[55])^(a[38] & b[56])^(a[37] & b[57])^(a[36] & b[58])^(a[35] & b[59])^(a[34] & b[60])^(a[33] & b[61])^(a[32] & b[62])^(a[31] & b[63])^(a[30] & b[64])^(a[29] & b[65])^(a[28] & b[66])^(a[27] & b[67])^(a[26] & b[68])^(a[25] & b[69])^(a[24] & b[70])^(a[23] & b[71])^(a[22] & b[72])^(a[21] & b[73])^(a[20] & b[74])^(a[19] & b[75])^(a[18] & b[76])^(a[17] & b[77])^(a[16] & b[78])^(a[15] & b[79])^(a[14] & b[80])^(a[13] & b[81])^(a[12] & b[82])^(a[11] & b[83])^(a[10] & b[84])^(a[9] & b[85])^(a[8] & b[86])^(a[7] & b[87])^(a[6] & b[88])^(a[5] & b[89])^(a[4] & b[90])^(a[3] & b[91])^(a[2] & b[92])^(a[1] & b[93])^(a[0] & b[94]);
assign y[95] = (a[95] & b[0])^(a[94] & b[1])^(a[93] & b[2])^(a[92] & b[3])^(a[91] & b[4])^(a[90] & b[5])^(a[89] & b[6])^(a[88] & b[7])^(a[87] & b[8])^(a[86] & b[9])^(a[85] & b[10])^(a[84] & b[11])^(a[83] & b[12])^(a[82] & b[13])^(a[81] & b[14])^(a[80] & b[15])^(a[79] & b[16])^(a[78] & b[17])^(a[77] & b[18])^(a[76] & b[19])^(a[75] & b[20])^(a[74] & b[21])^(a[73] & b[22])^(a[72] & b[23])^(a[71] & b[24])^(a[70] & b[25])^(a[69] & b[26])^(a[68] & b[27])^(a[67] & b[28])^(a[66] & b[29])^(a[65] & b[30])^(a[64] & b[31])^(a[63] & b[32])^(a[62] & b[33])^(a[61] & b[34])^(a[60] & b[35])^(a[59] & b[36])^(a[58] & b[37])^(a[57] & b[38])^(a[56] & b[39])^(a[55] & b[40])^(a[54] & b[41])^(a[53] & b[42])^(a[52] & b[43])^(a[51] & b[44])^(a[50] & b[45])^(a[49] & b[46])^(a[48] & b[47])^(a[47] & b[48])^(a[46] & b[49])^(a[45] & b[50])^(a[44] & b[51])^(a[43] & b[52])^(a[42] & b[53])^(a[41] & b[54])^(a[40] & b[55])^(a[39] & b[56])^(a[38] & b[57])^(a[37] & b[58])^(a[36] & b[59])^(a[35] & b[60])^(a[34] & b[61])^(a[33] & b[62])^(a[32] & b[63])^(a[31] & b[64])^(a[30] & b[65])^(a[29] & b[66])^(a[28] & b[67])^(a[27] & b[68])^(a[26] & b[69])^(a[25] & b[70])^(a[24] & b[71])^(a[23] & b[72])^(a[22] & b[73])^(a[21] & b[74])^(a[20] & b[75])^(a[19] & b[76])^(a[18] & b[77])^(a[17] & b[78])^(a[16] & b[79])^(a[15] & b[80])^(a[14] & b[81])^(a[13] & b[82])^(a[12] & b[83])^(a[11] & b[84])^(a[10] & b[85])^(a[9] & b[86])^(a[8] & b[87])^(a[7] & b[88])^(a[6] & b[89])^(a[5] & b[90])^(a[4] & b[91])^(a[3] & b[92])^(a[2] & b[93])^(a[1] & b[94])^(a[0] & b[95]);
assign y[96] = (a[96] & b[0])^(a[95] & b[1])^(a[94] & b[2])^(a[93] & b[3])^(a[92] & b[4])^(a[91] & b[5])^(a[90] & b[6])^(a[89] & b[7])^(a[88] & b[8])^(a[87] & b[9])^(a[86] & b[10])^(a[85] & b[11])^(a[84] & b[12])^(a[83] & b[13])^(a[82] & b[14])^(a[81] & b[15])^(a[80] & b[16])^(a[79] & b[17])^(a[78] & b[18])^(a[77] & b[19])^(a[76] & b[20])^(a[75] & b[21])^(a[74] & b[22])^(a[73] & b[23])^(a[72] & b[24])^(a[71] & b[25])^(a[70] & b[26])^(a[69] & b[27])^(a[68] & b[28])^(a[67] & b[29])^(a[66] & b[30])^(a[65] & b[31])^(a[64] & b[32])^(a[63] & b[33])^(a[62] & b[34])^(a[61] & b[35])^(a[60] & b[36])^(a[59] & b[37])^(a[58] & b[38])^(a[57] & b[39])^(a[56] & b[40])^(a[55] & b[41])^(a[54] & b[42])^(a[53] & b[43])^(a[52] & b[44])^(a[51] & b[45])^(a[50] & b[46])^(a[49] & b[47])^(a[48] & b[48])^(a[47] & b[49])^(a[46] & b[50])^(a[45] & b[51])^(a[44] & b[52])^(a[43] & b[53])^(a[42] & b[54])^(a[41] & b[55])^(a[40] & b[56])^(a[39] & b[57])^(a[38] & b[58])^(a[37] & b[59])^(a[36] & b[60])^(a[35] & b[61])^(a[34] & b[62])^(a[33] & b[63])^(a[32] & b[64])^(a[31] & b[65])^(a[30] & b[66])^(a[29] & b[67])^(a[28] & b[68])^(a[27] & b[69])^(a[26] & b[70])^(a[25] & b[71])^(a[24] & b[72])^(a[23] & b[73])^(a[22] & b[74])^(a[21] & b[75])^(a[20] & b[76])^(a[19] & b[77])^(a[18] & b[78])^(a[17] & b[79])^(a[16] & b[80])^(a[15] & b[81])^(a[14] & b[82])^(a[13] & b[83])^(a[12] & b[84])^(a[11] & b[85])^(a[10] & b[86])^(a[9] & b[87])^(a[8] & b[88])^(a[7] & b[89])^(a[6] & b[90])^(a[5] & b[91])^(a[4] & b[92])^(a[3] & b[93])^(a[2] & b[94])^(a[1] & b[95])^(a[0] & b[96]);
assign y[97] = (a[97] & b[0])^(a[96] & b[1])^(a[95] & b[2])^(a[94] & b[3])^(a[93] & b[4])^(a[92] & b[5])^(a[91] & b[6])^(a[90] & b[7])^(a[89] & b[8])^(a[88] & b[9])^(a[87] & b[10])^(a[86] & b[11])^(a[85] & b[12])^(a[84] & b[13])^(a[83] & b[14])^(a[82] & b[15])^(a[81] & b[16])^(a[80] & b[17])^(a[79] & b[18])^(a[78] & b[19])^(a[77] & b[20])^(a[76] & b[21])^(a[75] & b[22])^(a[74] & b[23])^(a[73] & b[24])^(a[72] & b[25])^(a[71] & b[26])^(a[70] & b[27])^(a[69] & b[28])^(a[68] & b[29])^(a[67] & b[30])^(a[66] & b[31])^(a[65] & b[32])^(a[64] & b[33])^(a[63] & b[34])^(a[62] & b[35])^(a[61] & b[36])^(a[60] & b[37])^(a[59] & b[38])^(a[58] & b[39])^(a[57] & b[40])^(a[56] & b[41])^(a[55] & b[42])^(a[54] & b[43])^(a[53] & b[44])^(a[52] & b[45])^(a[51] & b[46])^(a[50] & b[47])^(a[49] & b[48])^(a[48] & b[49])^(a[47] & b[50])^(a[46] & b[51])^(a[45] & b[52])^(a[44] & b[53])^(a[43] & b[54])^(a[42] & b[55])^(a[41] & b[56])^(a[40] & b[57])^(a[39] & b[58])^(a[38] & b[59])^(a[37] & b[60])^(a[36] & b[61])^(a[35] & b[62])^(a[34] & b[63])^(a[33] & b[64])^(a[32] & b[65])^(a[31] & b[66])^(a[30] & b[67])^(a[29] & b[68])^(a[28] & b[69])^(a[27] & b[70])^(a[26] & b[71])^(a[25] & b[72])^(a[24] & b[73])^(a[23] & b[74])^(a[22] & b[75])^(a[21] & b[76])^(a[20] & b[77])^(a[19] & b[78])^(a[18] & b[79])^(a[17] & b[80])^(a[16] & b[81])^(a[15] & b[82])^(a[14] & b[83])^(a[13] & b[84])^(a[12] & b[85])^(a[11] & b[86])^(a[10] & b[87])^(a[9] & b[88])^(a[8] & b[89])^(a[7] & b[90])^(a[6] & b[91])^(a[5] & b[92])^(a[4] & b[93])^(a[3] & b[94])^(a[2] & b[95])^(a[1] & b[96])^(a[0] & b[97]);
assign y[98] = (a[98] & b[0])^(a[97] & b[1])^(a[96] & b[2])^(a[95] & b[3])^(a[94] & b[4])^(a[93] & b[5])^(a[92] & b[6])^(a[91] & b[7])^(a[90] & b[8])^(a[89] & b[9])^(a[88] & b[10])^(a[87] & b[11])^(a[86] & b[12])^(a[85] & b[13])^(a[84] & b[14])^(a[83] & b[15])^(a[82] & b[16])^(a[81] & b[17])^(a[80] & b[18])^(a[79] & b[19])^(a[78] & b[20])^(a[77] & b[21])^(a[76] & b[22])^(a[75] & b[23])^(a[74] & b[24])^(a[73] & b[25])^(a[72] & b[26])^(a[71] & b[27])^(a[70] & b[28])^(a[69] & b[29])^(a[68] & b[30])^(a[67] & b[31])^(a[66] & b[32])^(a[65] & b[33])^(a[64] & b[34])^(a[63] & b[35])^(a[62] & b[36])^(a[61] & b[37])^(a[60] & b[38])^(a[59] & b[39])^(a[58] & b[40])^(a[57] & b[41])^(a[56] & b[42])^(a[55] & b[43])^(a[54] & b[44])^(a[53] & b[45])^(a[52] & b[46])^(a[51] & b[47])^(a[50] & b[48])^(a[49] & b[49])^(a[48] & b[50])^(a[47] & b[51])^(a[46] & b[52])^(a[45] & b[53])^(a[44] & b[54])^(a[43] & b[55])^(a[42] & b[56])^(a[41] & b[57])^(a[40] & b[58])^(a[39] & b[59])^(a[38] & b[60])^(a[37] & b[61])^(a[36] & b[62])^(a[35] & b[63])^(a[34] & b[64])^(a[33] & b[65])^(a[32] & b[66])^(a[31] & b[67])^(a[30] & b[68])^(a[29] & b[69])^(a[28] & b[70])^(a[27] & b[71])^(a[26] & b[72])^(a[25] & b[73])^(a[24] & b[74])^(a[23] & b[75])^(a[22] & b[76])^(a[21] & b[77])^(a[20] & b[78])^(a[19] & b[79])^(a[18] & b[80])^(a[17] & b[81])^(a[16] & b[82])^(a[15] & b[83])^(a[14] & b[84])^(a[13] & b[85])^(a[12] & b[86])^(a[11] & b[87])^(a[10] & b[88])^(a[9] & b[89])^(a[8] & b[90])^(a[7] & b[91])^(a[6] & b[92])^(a[5] & b[93])^(a[4] & b[94])^(a[3] & b[95])^(a[2] & b[96])^(a[1] & b[97])^(a[0] & b[98]);
assign y[99] = (a[99] & b[0])^(a[98] & b[1])^(a[97] & b[2])^(a[96] & b[3])^(a[95] & b[4])^(a[94] & b[5])^(a[93] & b[6])^(a[92] & b[7])^(a[91] & b[8])^(a[90] & b[9])^(a[89] & b[10])^(a[88] & b[11])^(a[87] & b[12])^(a[86] & b[13])^(a[85] & b[14])^(a[84] & b[15])^(a[83] & b[16])^(a[82] & b[17])^(a[81] & b[18])^(a[80] & b[19])^(a[79] & b[20])^(a[78] & b[21])^(a[77] & b[22])^(a[76] & b[23])^(a[75] & b[24])^(a[74] & b[25])^(a[73] & b[26])^(a[72] & b[27])^(a[71] & b[28])^(a[70] & b[29])^(a[69] & b[30])^(a[68] & b[31])^(a[67] & b[32])^(a[66] & b[33])^(a[65] & b[34])^(a[64] & b[35])^(a[63] & b[36])^(a[62] & b[37])^(a[61] & b[38])^(a[60] & b[39])^(a[59] & b[40])^(a[58] & b[41])^(a[57] & b[42])^(a[56] & b[43])^(a[55] & b[44])^(a[54] & b[45])^(a[53] & b[46])^(a[52] & b[47])^(a[51] & b[48])^(a[50] & b[49])^(a[49] & b[50])^(a[48] & b[51])^(a[47] & b[52])^(a[46] & b[53])^(a[45] & b[54])^(a[44] & b[55])^(a[43] & b[56])^(a[42] & b[57])^(a[41] & b[58])^(a[40] & b[59])^(a[39] & b[60])^(a[38] & b[61])^(a[37] & b[62])^(a[36] & b[63])^(a[35] & b[64])^(a[34] & b[65])^(a[33] & b[66])^(a[32] & b[67])^(a[31] & b[68])^(a[30] & b[69])^(a[29] & b[70])^(a[28] & b[71])^(a[27] & b[72])^(a[26] & b[73])^(a[25] & b[74])^(a[24] & b[75])^(a[23] & b[76])^(a[22] & b[77])^(a[21] & b[78])^(a[20] & b[79])^(a[19] & b[80])^(a[18] & b[81])^(a[17] & b[82])^(a[16] & b[83])^(a[15] & b[84])^(a[14] & b[85])^(a[13] & b[86])^(a[12] & b[87])^(a[11] & b[88])^(a[10] & b[89])^(a[9] & b[90])^(a[8] & b[91])^(a[7] & b[92])^(a[6] & b[93])^(a[5] & b[94])^(a[4] & b[95])^(a[3] & b[96])^(a[2] & b[97])^(a[1] & b[98])^(a[0] & b[99]);
assign y[100] = (a[100] & b[0])^(a[99] & b[1])^(a[98] & b[2])^(a[97] & b[3])^(a[96] & b[4])^(a[95] & b[5])^(a[94] & b[6])^(a[93] & b[7])^(a[92] & b[8])^(a[91] & b[9])^(a[90] & b[10])^(a[89] & b[11])^(a[88] & b[12])^(a[87] & b[13])^(a[86] & b[14])^(a[85] & b[15])^(a[84] & b[16])^(a[83] & b[17])^(a[82] & b[18])^(a[81] & b[19])^(a[80] & b[20])^(a[79] & b[21])^(a[78] & b[22])^(a[77] & b[23])^(a[76] & b[24])^(a[75] & b[25])^(a[74] & b[26])^(a[73] & b[27])^(a[72] & b[28])^(a[71] & b[29])^(a[70] & b[30])^(a[69] & b[31])^(a[68] & b[32])^(a[67] & b[33])^(a[66] & b[34])^(a[65] & b[35])^(a[64] & b[36])^(a[63] & b[37])^(a[62] & b[38])^(a[61] & b[39])^(a[60] & b[40])^(a[59] & b[41])^(a[58] & b[42])^(a[57] & b[43])^(a[56] & b[44])^(a[55] & b[45])^(a[54] & b[46])^(a[53] & b[47])^(a[52] & b[48])^(a[51] & b[49])^(a[50] & b[50])^(a[49] & b[51])^(a[48] & b[52])^(a[47] & b[53])^(a[46] & b[54])^(a[45] & b[55])^(a[44] & b[56])^(a[43] & b[57])^(a[42] & b[58])^(a[41] & b[59])^(a[40] & b[60])^(a[39] & b[61])^(a[38] & b[62])^(a[37] & b[63])^(a[36] & b[64])^(a[35] & b[65])^(a[34] & b[66])^(a[33] & b[67])^(a[32] & b[68])^(a[31] & b[69])^(a[30] & b[70])^(a[29] & b[71])^(a[28] & b[72])^(a[27] & b[73])^(a[26] & b[74])^(a[25] & b[75])^(a[24] & b[76])^(a[23] & b[77])^(a[22] & b[78])^(a[21] & b[79])^(a[20] & b[80])^(a[19] & b[81])^(a[18] & b[82])^(a[17] & b[83])^(a[16] & b[84])^(a[15] & b[85])^(a[14] & b[86])^(a[13] & b[87])^(a[12] & b[88])^(a[11] & b[89])^(a[10] & b[90])^(a[9] & b[91])^(a[8] & b[92])^(a[7] & b[93])^(a[6] & b[94])^(a[5] & b[95])^(a[4] & b[96])^(a[3] & b[97])^(a[2] & b[98])^(a[1] & b[99])^(a[0] & b[100]);
assign y[101] = (a[101] & b[0])^(a[100] & b[1])^(a[99] & b[2])^(a[98] & b[3])^(a[97] & b[4])^(a[96] & b[5])^(a[95] & b[6])^(a[94] & b[7])^(a[93] & b[8])^(a[92] & b[9])^(a[91] & b[10])^(a[90] & b[11])^(a[89] & b[12])^(a[88] & b[13])^(a[87] & b[14])^(a[86] & b[15])^(a[85] & b[16])^(a[84] & b[17])^(a[83] & b[18])^(a[82] & b[19])^(a[81] & b[20])^(a[80] & b[21])^(a[79] & b[22])^(a[78] & b[23])^(a[77] & b[24])^(a[76] & b[25])^(a[75] & b[26])^(a[74] & b[27])^(a[73] & b[28])^(a[72] & b[29])^(a[71] & b[30])^(a[70] & b[31])^(a[69] & b[32])^(a[68] & b[33])^(a[67] & b[34])^(a[66] & b[35])^(a[65] & b[36])^(a[64] & b[37])^(a[63] & b[38])^(a[62] & b[39])^(a[61] & b[40])^(a[60] & b[41])^(a[59] & b[42])^(a[58] & b[43])^(a[57] & b[44])^(a[56] & b[45])^(a[55] & b[46])^(a[54] & b[47])^(a[53] & b[48])^(a[52] & b[49])^(a[51] & b[50])^(a[50] & b[51])^(a[49] & b[52])^(a[48] & b[53])^(a[47] & b[54])^(a[46] & b[55])^(a[45] & b[56])^(a[44] & b[57])^(a[43] & b[58])^(a[42] & b[59])^(a[41] & b[60])^(a[40] & b[61])^(a[39] & b[62])^(a[38] & b[63])^(a[37] & b[64])^(a[36] & b[65])^(a[35] & b[66])^(a[34] & b[67])^(a[33] & b[68])^(a[32] & b[69])^(a[31] & b[70])^(a[30] & b[71])^(a[29] & b[72])^(a[28] & b[73])^(a[27] & b[74])^(a[26] & b[75])^(a[25] & b[76])^(a[24] & b[77])^(a[23] & b[78])^(a[22] & b[79])^(a[21] & b[80])^(a[20] & b[81])^(a[19] & b[82])^(a[18] & b[83])^(a[17] & b[84])^(a[16] & b[85])^(a[15] & b[86])^(a[14] & b[87])^(a[13] & b[88])^(a[12] & b[89])^(a[11] & b[90])^(a[10] & b[91])^(a[9] & b[92])^(a[8] & b[93])^(a[7] & b[94])^(a[6] & b[95])^(a[5] & b[96])^(a[4] & b[97])^(a[3] & b[98])^(a[2] & b[99])^(a[1] & b[100])^(a[0] & b[101]);
assign y[102] = (a[102] & b[0])^(a[101] & b[1])^(a[100] & b[2])^(a[99] & b[3])^(a[98] & b[4])^(a[97] & b[5])^(a[96] & b[6])^(a[95] & b[7])^(a[94] & b[8])^(a[93] & b[9])^(a[92] & b[10])^(a[91] & b[11])^(a[90] & b[12])^(a[89] & b[13])^(a[88] & b[14])^(a[87] & b[15])^(a[86] & b[16])^(a[85] & b[17])^(a[84] & b[18])^(a[83] & b[19])^(a[82] & b[20])^(a[81] & b[21])^(a[80] & b[22])^(a[79] & b[23])^(a[78] & b[24])^(a[77] & b[25])^(a[76] & b[26])^(a[75] & b[27])^(a[74] & b[28])^(a[73] & b[29])^(a[72] & b[30])^(a[71] & b[31])^(a[70] & b[32])^(a[69] & b[33])^(a[68] & b[34])^(a[67] & b[35])^(a[66] & b[36])^(a[65] & b[37])^(a[64] & b[38])^(a[63] & b[39])^(a[62] & b[40])^(a[61] & b[41])^(a[60] & b[42])^(a[59] & b[43])^(a[58] & b[44])^(a[57] & b[45])^(a[56] & b[46])^(a[55] & b[47])^(a[54] & b[48])^(a[53] & b[49])^(a[52] & b[50])^(a[51] & b[51])^(a[50] & b[52])^(a[49] & b[53])^(a[48] & b[54])^(a[47] & b[55])^(a[46] & b[56])^(a[45] & b[57])^(a[44] & b[58])^(a[43] & b[59])^(a[42] & b[60])^(a[41] & b[61])^(a[40] & b[62])^(a[39] & b[63])^(a[38] & b[64])^(a[37] & b[65])^(a[36] & b[66])^(a[35] & b[67])^(a[34] & b[68])^(a[33] & b[69])^(a[32] & b[70])^(a[31] & b[71])^(a[30] & b[72])^(a[29] & b[73])^(a[28] & b[74])^(a[27] & b[75])^(a[26] & b[76])^(a[25] & b[77])^(a[24] & b[78])^(a[23] & b[79])^(a[22] & b[80])^(a[21] & b[81])^(a[20] & b[82])^(a[19] & b[83])^(a[18] & b[84])^(a[17] & b[85])^(a[16] & b[86])^(a[15] & b[87])^(a[14] & b[88])^(a[13] & b[89])^(a[12] & b[90])^(a[11] & b[91])^(a[10] & b[92])^(a[9] & b[93])^(a[8] & b[94])^(a[7] & b[95])^(a[6] & b[96])^(a[5] & b[97])^(a[4] & b[98])^(a[3] & b[99])^(a[2] & b[100])^(a[1] & b[101])^(a[0] & b[102]);
assign y[103] = (a[103] & b[0])^(a[102] & b[1])^(a[101] & b[2])^(a[100] & b[3])^(a[99] & b[4])^(a[98] & b[5])^(a[97] & b[6])^(a[96] & b[7])^(a[95] & b[8])^(a[94] & b[9])^(a[93] & b[10])^(a[92] & b[11])^(a[91] & b[12])^(a[90] & b[13])^(a[89] & b[14])^(a[88] & b[15])^(a[87] & b[16])^(a[86] & b[17])^(a[85] & b[18])^(a[84] & b[19])^(a[83] & b[20])^(a[82] & b[21])^(a[81] & b[22])^(a[80] & b[23])^(a[79] & b[24])^(a[78] & b[25])^(a[77] & b[26])^(a[76] & b[27])^(a[75] & b[28])^(a[74] & b[29])^(a[73] & b[30])^(a[72] & b[31])^(a[71] & b[32])^(a[70] & b[33])^(a[69] & b[34])^(a[68] & b[35])^(a[67] & b[36])^(a[66] & b[37])^(a[65] & b[38])^(a[64] & b[39])^(a[63] & b[40])^(a[62] & b[41])^(a[61] & b[42])^(a[60] & b[43])^(a[59] & b[44])^(a[58] & b[45])^(a[57] & b[46])^(a[56] & b[47])^(a[55] & b[48])^(a[54] & b[49])^(a[53] & b[50])^(a[52] & b[51])^(a[51] & b[52])^(a[50] & b[53])^(a[49] & b[54])^(a[48] & b[55])^(a[47] & b[56])^(a[46] & b[57])^(a[45] & b[58])^(a[44] & b[59])^(a[43] & b[60])^(a[42] & b[61])^(a[41] & b[62])^(a[40] & b[63])^(a[39] & b[64])^(a[38] & b[65])^(a[37] & b[66])^(a[36] & b[67])^(a[35] & b[68])^(a[34] & b[69])^(a[33] & b[70])^(a[32] & b[71])^(a[31] & b[72])^(a[30] & b[73])^(a[29] & b[74])^(a[28] & b[75])^(a[27] & b[76])^(a[26] & b[77])^(a[25] & b[78])^(a[24] & b[79])^(a[23] & b[80])^(a[22] & b[81])^(a[21] & b[82])^(a[20] & b[83])^(a[19] & b[84])^(a[18] & b[85])^(a[17] & b[86])^(a[16] & b[87])^(a[15] & b[88])^(a[14] & b[89])^(a[13] & b[90])^(a[12] & b[91])^(a[11] & b[92])^(a[10] & b[93])^(a[9] & b[94])^(a[8] & b[95])^(a[7] & b[96])^(a[6] & b[97])^(a[5] & b[98])^(a[4] & b[99])^(a[3] & b[100])^(a[2] & b[101])^(a[1] & b[102])^(a[0] & b[103]);
assign y[104] = (a[104] & b[0])^(a[103] & b[1])^(a[102] & b[2])^(a[101] & b[3])^(a[100] & b[4])^(a[99] & b[5])^(a[98] & b[6])^(a[97] & b[7])^(a[96] & b[8])^(a[95] & b[9])^(a[94] & b[10])^(a[93] & b[11])^(a[92] & b[12])^(a[91] & b[13])^(a[90] & b[14])^(a[89] & b[15])^(a[88] & b[16])^(a[87] & b[17])^(a[86] & b[18])^(a[85] & b[19])^(a[84] & b[20])^(a[83] & b[21])^(a[82] & b[22])^(a[81] & b[23])^(a[80] & b[24])^(a[79] & b[25])^(a[78] & b[26])^(a[77] & b[27])^(a[76] & b[28])^(a[75] & b[29])^(a[74] & b[30])^(a[73] & b[31])^(a[72] & b[32])^(a[71] & b[33])^(a[70] & b[34])^(a[69] & b[35])^(a[68] & b[36])^(a[67] & b[37])^(a[66] & b[38])^(a[65] & b[39])^(a[64] & b[40])^(a[63] & b[41])^(a[62] & b[42])^(a[61] & b[43])^(a[60] & b[44])^(a[59] & b[45])^(a[58] & b[46])^(a[57] & b[47])^(a[56] & b[48])^(a[55] & b[49])^(a[54] & b[50])^(a[53] & b[51])^(a[52] & b[52])^(a[51] & b[53])^(a[50] & b[54])^(a[49] & b[55])^(a[48] & b[56])^(a[47] & b[57])^(a[46] & b[58])^(a[45] & b[59])^(a[44] & b[60])^(a[43] & b[61])^(a[42] & b[62])^(a[41] & b[63])^(a[40] & b[64])^(a[39] & b[65])^(a[38] & b[66])^(a[37] & b[67])^(a[36] & b[68])^(a[35] & b[69])^(a[34] & b[70])^(a[33] & b[71])^(a[32] & b[72])^(a[31] & b[73])^(a[30] & b[74])^(a[29] & b[75])^(a[28] & b[76])^(a[27] & b[77])^(a[26] & b[78])^(a[25] & b[79])^(a[24] & b[80])^(a[23] & b[81])^(a[22] & b[82])^(a[21] & b[83])^(a[20] & b[84])^(a[19] & b[85])^(a[18] & b[86])^(a[17] & b[87])^(a[16] & b[88])^(a[15] & b[89])^(a[14] & b[90])^(a[13] & b[91])^(a[12] & b[92])^(a[11] & b[93])^(a[10] & b[94])^(a[9] & b[95])^(a[8] & b[96])^(a[7] & b[97])^(a[6] & b[98])^(a[5] & b[99])^(a[4] & b[100])^(a[3] & b[101])^(a[2] & b[102])^(a[1] & b[103])^(a[0] & b[104]);
assign y[105] = (a[105] & b[0])^(a[104] & b[1])^(a[103] & b[2])^(a[102] & b[3])^(a[101] & b[4])^(a[100] & b[5])^(a[99] & b[6])^(a[98] & b[7])^(a[97] & b[8])^(a[96] & b[9])^(a[95] & b[10])^(a[94] & b[11])^(a[93] & b[12])^(a[92] & b[13])^(a[91] & b[14])^(a[90] & b[15])^(a[89] & b[16])^(a[88] & b[17])^(a[87] & b[18])^(a[86] & b[19])^(a[85] & b[20])^(a[84] & b[21])^(a[83] & b[22])^(a[82] & b[23])^(a[81] & b[24])^(a[80] & b[25])^(a[79] & b[26])^(a[78] & b[27])^(a[77] & b[28])^(a[76] & b[29])^(a[75] & b[30])^(a[74] & b[31])^(a[73] & b[32])^(a[72] & b[33])^(a[71] & b[34])^(a[70] & b[35])^(a[69] & b[36])^(a[68] & b[37])^(a[67] & b[38])^(a[66] & b[39])^(a[65] & b[40])^(a[64] & b[41])^(a[63] & b[42])^(a[62] & b[43])^(a[61] & b[44])^(a[60] & b[45])^(a[59] & b[46])^(a[58] & b[47])^(a[57] & b[48])^(a[56] & b[49])^(a[55] & b[50])^(a[54] & b[51])^(a[53] & b[52])^(a[52] & b[53])^(a[51] & b[54])^(a[50] & b[55])^(a[49] & b[56])^(a[48] & b[57])^(a[47] & b[58])^(a[46] & b[59])^(a[45] & b[60])^(a[44] & b[61])^(a[43] & b[62])^(a[42] & b[63])^(a[41] & b[64])^(a[40] & b[65])^(a[39] & b[66])^(a[38] & b[67])^(a[37] & b[68])^(a[36] & b[69])^(a[35] & b[70])^(a[34] & b[71])^(a[33] & b[72])^(a[32] & b[73])^(a[31] & b[74])^(a[30] & b[75])^(a[29] & b[76])^(a[28] & b[77])^(a[27] & b[78])^(a[26] & b[79])^(a[25] & b[80])^(a[24] & b[81])^(a[23] & b[82])^(a[22] & b[83])^(a[21] & b[84])^(a[20] & b[85])^(a[19] & b[86])^(a[18] & b[87])^(a[17] & b[88])^(a[16] & b[89])^(a[15] & b[90])^(a[14] & b[91])^(a[13] & b[92])^(a[12] & b[93])^(a[11] & b[94])^(a[10] & b[95])^(a[9] & b[96])^(a[8] & b[97])^(a[7] & b[98])^(a[6] & b[99])^(a[5] & b[100])^(a[4] & b[101])^(a[3] & b[102])^(a[2] & b[103])^(a[1] & b[104])^(a[0] & b[105]);
assign y[106] = (a[106] & b[0])^(a[105] & b[1])^(a[104] & b[2])^(a[103] & b[3])^(a[102] & b[4])^(a[101] & b[5])^(a[100] & b[6])^(a[99] & b[7])^(a[98] & b[8])^(a[97] & b[9])^(a[96] & b[10])^(a[95] & b[11])^(a[94] & b[12])^(a[93] & b[13])^(a[92] & b[14])^(a[91] & b[15])^(a[90] & b[16])^(a[89] & b[17])^(a[88] & b[18])^(a[87] & b[19])^(a[86] & b[20])^(a[85] & b[21])^(a[84] & b[22])^(a[83] & b[23])^(a[82] & b[24])^(a[81] & b[25])^(a[80] & b[26])^(a[79] & b[27])^(a[78] & b[28])^(a[77] & b[29])^(a[76] & b[30])^(a[75] & b[31])^(a[74] & b[32])^(a[73] & b[33])^(a[72] & b[34])^(a[71] & b[35])^(a[70] & b[36])^(a[69] & b[37])^(a[68] & b[38])^(a[67] & b[39])^(a[66] & b[40])^(a[65] & b[41])^(a[64] & b[42])^(a[63] & b[43])^(a[62] & b[44])^(a[61] & b[45])^(a[60] & b[46])^(a[59] & b[47])^(a[58] & b[48])^(a[57] & b[49])^(a[56] & b[50])^(a[55] & b[51])^(a[54] & b[52])^(a[53] & b[53])^(a[52] & b[54])^(a[51] & b[55])^(a[50] & b[56])^(a[49] & b[57])^(a[48] & b[58])^(a[47] & b[59])^(a[46] & b[60])^(a[45] & b[61])^(a[44] & b[62])^(a[43] & b[63])^(a[42] & b[64])^(a[41] & b[65])^(a[40] & b[66])^(a[39] & b[67])^(a[38] & b[68])^(a[37] & b[69])^(a[36] & b[70])^(a[35] & b[71])^(a[34] & b[72])^(a[33] & b[73])^(a[32] & b[74])^(a[31] & b[75])^(a[30] & b[76])^(a[29] & b[77])^(a[28] & b[78])^(a[27] & b[79])^(a[26] & b[80])^(a[25] & b[81])^(a[24] & b[82])^(a[23] & b[83])^(a[22] & b[84])^(a[21] & b[85])^(a[20] & b[86])^(a[19] & b[87])^(a[18] & b[88])^(a[17] & b[89])^(a[16] & b[90])^(a[15] & b[91])^(a[14] & b[92])^(a[13] & b[93])^(a[12] & b[94])^(a[11] & b[95])^(a[10] & b[96])^(a[9] & b[97])^(a[8] & b[98])^(a[7] & b[99])^(a[6] & b[100])^(a[5] & b[101])^(a[4] & b[102])^(a[3] & b[103])^(a[2] & b[104])^(a[1] & b[105])^(a[0] & b[106]);
assign y[107] = (a[107] & b[0])^(a[106] & b[1])^(a[105] & b[2])^(a[104] & b[3])^(a[103] & b[4])^(a[102] & b[5])^(a[101] & b[6])^(a[100] & b[7])^(a[99] & b[8])^(a[98] & b[9])^(a[97] & b[10])^(a[96] & b[11])^(a[95] & b[12])^(a[94] & b[13])^(a[93] & b[14])^(a[92] & b[15])^(a[91] & b[16])^(a[90] & b[17])^(a[89] & b[18])^(a[88] & b[19])^(a[87] & b[20])^(a[86] & b[21])^(a[85] & b[22])^(a[84] & b[23])^(a[83] & b[24])^(a[82] & b[25])^(a[81] & b[26])^(a[80] & b[27])^(a[79] & b[28])^(a[78] & b[29])^(a[77] & b[30])^(a[76] & b[31])^(a[75] & b[32])^(a[74] & b[33])^(a[73] & b[34])^(a[72] & b[35])^(a[71] & b[36])^(a[70] & b[37])^(a[69] & b[38])^(a[68] & b[39])^(a[67] & b[40])^(a[66] & b[41])^(a[65] & b[42])^(a[64] & b[43])^(a[63] & b[44])^(a[62] & b[45])^(a[61] & b[46])^(a[60] & b[47])^(a[59] & b[48])^(a[58] & b[49])^(a[57] & b[50])^(a[56] & b[51])^(a[55] & b[52])^(a[54] & b[53])^(a[53] & b[54])^(a[52] & b[55])^(a[51] & b[56])^(a[50] & b[57])^(a[49] & b[58])^(a[48] & b[59])^(a[47] & b[60])^(a[46] & b[61])^(a[45] & b[62])^(a[44] & b[63])^(a[43] & b[64])^(a[42] & b[65])^(a[41] & b[66])^(a[40] & b[67])^(a[39] & b[68])^(a[38] & b[69])^(a[37] & b[70])^(a[36] & b[71])^(a[35] & b[72])^(a[34] & b[73])^(a[33] & b[74])^(a[32] & b[75])^(a[31] & b[76])^(a[30] & b[77])^(a[29] & b[78])^(a[28] & b[79])^(a[27] & b[80])^(a[26] & b[81])^(a[25] & b[82])^(a[24] & b[83])^(a[23] & b[84])^(a[22] & b[85])^(a[21] & b[86])^(a[20] & b[87])^(a[19] & b[88])^(a[18] & b[89])^(a[17] & b[90])^(a[16] & b[91])^(a[15] & b[92])^(a[14] & b[93])^(a[13] & b[94])^(a[12] & b[95])^(a[11] & b[96])^(a[10] & b[97])^(a[9] & b[98])^(a[8] & b[99])^(a[7] & b[100])^(a[6] & b[101])^(a[5] & b[102])^(a[4] & b[103])^(a[3] & b[104])^(a[2] & b[105])^(a[1] & b[106])^(a[0] & b[107]);
assign y[108] = (a[108] & b[0])^(a[107] & b[1])^(a[106] & b[2])^(a[105] & b[3])^(a[104] & b[4])^(a[103] & b[5])^(a[102] & b[6])^(a[101] & b[7])^(a[100] & b[8])^(a[99] & b[9])^(a[98] & b[10])^(a[97] & b[11])^(a[96] & b[12])^(a[95] & b[13])^(a[94] & b[14])^(a[93] & b[15])^(a[92] & b[16])^(a[91] & b[17])^(a[90] & b[18])^(a[89] & b[19])^(a[88] & b[20])^(a[87] & b[21])^(a[86] & b[22])^(a[85] & b[23])^(a[84] & b[24])^(a[83] & b[25])^(a[82] & b[26])^(a[81] & b[27])^(a[80] & b[28])^(a[79] & b[29])^(a[78] & b[30])^(a[77] & b[31])^(a[76] & b[32])^(a[75] & b[33])^(a[74] & b[34])^(a[73] & b[35])^(a[72] & b[36])^(a[71] & b[37])^(a[70] & b[38])^(a[69] & b[39])^(a[68] & b[40])^(a[67] & b[41])^(a[66] & b[42])^(a[65] & b[43])^(a[64] & b[44])^(a[63] & b[45])^(a[62] & b[46])^(a[61] & b[47])^(a[60] & b[48])^(a[59] & b[49])^(a[58] & b[50])^(a[57] & b[51])^(a[56] & b[52])^(a[55] & b[53])^(a[54] & b[54])^(a[53] & b[55])^(a[52] & b[56])^(a[51] & b[57])^(a[50] & b[58])^(a[49] & b[59])^(a[48] & b[60])^(a[47] & b[61])^(a[46] & b[62])^(a[45] & b[63])^(a[44] & b[64])^(a[43] & b[65])^(a[42] & b[66])^(a[41] & b[67])^(a[40] & b[68])^(a[39] & b[69])^(a[38] & b[70])^(a[37] & b[71])^(a[36] & b[72])^(a[35] & b[73])^(a[34] & b[74])^(a[33] & b[75])^(a[32] & b[76])^(a[31] & b[77])^(a[30] & b[78])^(a[29] & b[79])^(a[28] & b[80])^(a[27] & b[81])^(a[26] & b[82])^(a[25] & b[83])^(a[24] & b[84])^(a[23] & b[85])^(a[22] & b[86])^(a[21] & b[87])^(a[20] & b[88])^(a[19] & b[89])^(a[18] & b[90])^(a[17] & b[91])^(a[16] & b[92])^(a[15] & b[93])^(a[14] & b[94])^(a[13] & b[95])^(a[12] & b[96])^(a[11] & b[97])^(a[10] & b[98])^(a[9] & b[99])^(a[8] & b[100])^(a[7] & b[101])^(a[6] & b[102])^(a[5] & b[103])^(a[4] & b[104])^(a[3] & b[105])^(a[2] & b[106])^(a[1] & b[107])^(a[0] & b[108]);
assign y[109] = (a[109] & b[0])^(a[108] & b[1])^(a[107] & b[2])^(a[106] & b[3])^(a[105] & b[4])^(a[104] & b[5])^(a[103] & b[6])^(a[102] & b[7])^(a[101] & b[8])^(a[100] & b[9])^(a[99] & b[10])^(a[98] & b[11])^(a[97] & b[12])^(a[96] & b[13])^(a[95] & b[14])^(a[94] & b[15])^(a[93] & b[16])^(a[92] & b[17])^(a[91] & b[18])^(a[90] & b[19])^(a[89] & b[20])^(a[88] & b[21])^(a[87] & b[22])^(a[86] & b[23])^(a[85] & b[24])^(a[84] & b[25])^(a[83] & b[26])^(a[82] & b[27])^(a[81] & b[28])^(a[80] & b[29])^(a[79] & b[30])^(a[78] & b[31])^(a[77] & b[32])^(a[76] & b[33])^(a[75] & b[34])^(a[74] & b[35])^(a[73] & b[36])^(a[72] & b[37])^(a[71] & b[38])^(a[70] & b[39])^(a[69] & b[40])^(a[68] & b[41])^(a[67] & b[42])^(a[66] & b[43])^(a[65] & b[44])^(a[64] & b[45])^(a[63] & b[46])^(a[62] & b[47])^(a[61] & b[48])^(a[60] & b[49])^(a[59] & b[50])^(a[58] & b[51])^(a[57] & b[52])^(a[56] & b[53])^(a[55] & b[54])^(a[54] & b[55])^(a[53] & b[56])^(a[52] & b[57])^(a[51] & b[58])^(a[50] & b[59])^(a[49] & b[60])^(a[48] & b[61])^(a[47] & b[62])^(a[46] & b[63])^(a[45] & b[64])^(a[44] & b[65])^(a[43] & b[66])^(a[42] & b[67])^(a[41] & b[68])^(a[40] & b[69])^(a[39] & b[70])^(a[38] & b[71])^(a[37] & b[72])^(a[36] & b[73])^(a[35] & b[74])^(a[34] & b[75])^(a[33] & b[76])^(a[32] & b[77])^(a[31] & b[78])^(a[30] & b[79])^(a[29] & b[80])^(a[28] & b[81])^(a[27] & b[82])^(a[26] & b[83])^(a[25] & b[84])^(a[24] & b[85])^(a[23] & b[86])^(a[22] & b[87])^(a[21] & b[88])^(a[20] & b[89])^(a[19] & b[90])^(a[18] & b[91])^(a[17] & b[92])^(a[16] & b[93])^(a[15] & b[94])^(a[14] & b[95])^(a[13] & b[96])^(a[12] & b[97])^(a[11] & b[98])^(a[10] & b[99])^(a[9] & b[100])^(a[8] & b[101])^(a[7] & b[102])^(a[6] & b[103])^(a[5] & b[104])^(a[4] & b[105])^(a[3] & b[106])^(a[2] & b[107])^(a[1] & b[108])^(a[0] & b[109]);
assign y[110] = (a[110] & b[0])^(a[109] & b[1])^(a[108] & b[2])^(a[107] & b[3])^(a[106] & b[4])^(a[105] & b[5])^(a[104] & b[6])^(a[103] & b[7])^(a[102] & b[8])^(a[101] & b[9])^(a[100] & b[10])^(a[99] & b[11])^(a[98] & b[12])^(a[97] & b[13])^(a[96] & b[14])^(a[95] & b[15])^(a[94] & b[16])^(a[93] & b[17])^(a[92] & b[18])^(a[91] & b[19])^(a[90] & b[20])^(a[89] & b[21])^(a[88] & b[22])^(a[87] & b[23])^(a[86] & b[24])^(a[85] & b[25])^(a[84] & b[26])^(a[83] & b[27])^(a[82] & b[28])^(a[81] & b[29])^(a[80] & b[30])^(a[79] & b[31])^(a[78] & b[32])^(a[77] & b[33])^(a[76] & b[34])^(a[75] & b[35])^(a[74] & b[36])^(a[73] & b[37])^(a[72] & b[38])^(a[71] & b[39])^(a[70] & b[40])^(a[69] & b[41])^(a[68] & b[42])^(a[67] & b[43])^(a[66] & b[44])^(a[65] & b[45])^(a[64] & b[46])^(a[63] & b[47])^(a[62] & b[48])^(a[61] & b[49])^(a[60] & b[50])^(a[59] & b[51])^(a[58] & b[52])^(a[57] & b[53])^(a[56] & b[54])^(a[55] & b[55])^(a[54] & b[56])^(a[53] & b[57])^(a[52] & b[58])^(a[51] & b[59])^(a[50] & b[60])^(a[49] & b[61])^(a[48] & b[62])^(a[47] & b[63])^(a[46] & b[64])^(a[45] & b[65])^(a[44] & b[66])^(a[43] & b[67])^(a[42] & b[68])^(a[41] & b[69])^(a[40] & b[70])^(a[39] & b[71])^(a[38] & b[72])^(a[37] & b[73])^(a[36] & b[74])^(a[35] & b[75])^(a[34] & b[76])^(a[33] & b[77])^(a[32] & b[78])^(a[31] & b[79])^(a[30] & b[80])^(a[29] & b[81])^(a[28] & b[82])^(a[27] & b[83])^(a[26] & b[84])^(a[25] & b[85])^(a[24] & b[86])^(a[23] & b[87])^(a[22] & b[88])^(a[21] & b[89])^(a[20] & b[90])^(a[19] & b[91])^(a[18] & b[92])^(a[17] & b[93])^(a[16] & b[94])^(a[15] & b[95])^(a[14] & b[96])^(a[13] & b[97])^(a[12] & b[98])^(a[11] & b[99])^(a[10] & b[100])^(a[9] & b[101])^(a[8] & b[102])^(a[7] & b[103])^(a[6] & b[104])^(a[5] & b[105])^(a[4] & b[106])^(a[3] & b[107])^(a[2] & b[108])^(a[1] & b[109])^(a[0] & b[110]);
assign y[111] = (a[111] & b[0])^(a[110] & b[1])^(a[109] & b[2])^(a[108] & b[3])^(a[107] & b[4])^(a[106] & b[5])^(a[105] & b[6])^(a[104] & b[7])^(a[103] & b[8])^(a[102] & b[9])^(a[101] & b[10])^(a[100] & b[11])^(a[99] & b[12])^(a[98] & b[13])^(a[97] & b[14])^(a[96] & b[15])^(a[95] & b[16])^(a[94] & b[17])^(a[93] & b[18])^(a[92] & b[19])^(a[91] & b[20])^(a[90] & b[21])^(a[89] & b[22])^(a[88] & b[23])^(a[87] & b[24])^(a[86] & b[25])^(a[85] & b[26])^(a[84] & b[27])^(a[83] & b[28])^(a[82] & b[29])^(a[81] & b[30])^(a[80] & b[31])^(a[79] & b[32])^(a[78] & b[33])^(a[77] & b[34])^(a[76] & b[35])^(a[75] & b[36])^(a[74] & b[37])^(a[73] & b[38])^(a[72] & b[39])^(a[71] & b[40])^(a[70] & b[41])^(a[69] & b[42])^(a[68] & b[43])^(a[67] & b[44])^(a[66] & b[45])^(a[65] & b[46])^(a[64] & b[47])^(a[63] & b[48])^(a[62] & b[49])^(a[61] & b[50])^(a[60] & b[51])^(a[59] & b[52])^(a[58] & b[53])^(a[57] & b[54])^(a[56] & b[55])^(a[55] & b[56])^(a[54] & b[57])^(a[53] & b[58])^(a[52] & b[59])^(a[51] & b[60])^(a[50] & b[61])^(a[49] & b[62])^(a[48] & b[63])^(a[47] & b[64])^(a[46] & b[65])^(a[45] & b[66])^(a[44] & b[67])^(a[43] & b[68])^(a[42] & b[69])^(a[41] & b[70])^(a[40] & b[71])^(a[39] & b[72])^(a[38] & b[73])^(a[37] & b[74])^(a[36] & b[75])^(a[35] & b[76])^(a[34] & b[77])^(a[33] & b[78])^(a[32] & b[79])^(a[31] & b[80])^(a[30] & b[81])^(a[29] & b[82])^(a[28] & b[83])^(a[27] & b[84])^(a[26] & b[85])^(a[25] & b[86])^(a[24] & b[87])^(a[23] & b[88])^(a[22] & b[89])^(a[21] & b[90])^(a[20] & b[91])^(a[19] & b[92])^(a[18] & b[93])^(a[17] & b[94])^(a[16] & b[95])^(a[15] & b[96])^(a[14] & b[97])^(a[13] & b[98])^(a[12] & b[99])^(a[11] & b[100])^(a[10] & b[101])^(a[9] & b[102])^(a[8] & b[103])^(a[7] & b[104])^(a[6] & b[105])^(a[5] & b[106])^(a[4] & b[107])^(a[3] & b[108])^(a[2] & b[109])^(a[1] & b[110])^(a[0] & b[111]);
assign y[112] = (a[112] & b[0])^(a[111] & b[1])^(a[110] & b[2])^(a[109] & b[3])^(a[108] & b[4])^(a[107] & b[5])^(a[106] & b[6])^(a[105] & b[7])^(a[104] & b[8])^(a[103] & b[9])^(a[102] & b[10])^(a[101] & b[11])^(a[100] & b[12])^(a[99] & b[13])^(a[98] & b[14])^(a[97] & b[15])^(a[96] & b[16])^(a[95] & b[17])^(a[94] & b[18])^(a[93] & b[19])^(a[92] & b[20])^(a[91] & b[21])^(a[90] & b[22])^(a[89] & b[23])^(a[88] & b[24])^(a[87] & b[25])^(a[86] & b[26])^(a[85] & b[27])^(a[84] & b[28])^(a[83] & b[29])^(a[82] & b[30])^(a[81] & b[31])^(a[80] & b[32])^(a[79] & b[33])^(a[78] & b[34])^(a[77] & b[35])^(a[76] & b[36])^(a[75] & b[37])^(a[74] & b[38])^(a[73] & b[39])^(a[72] & b[40])^(a[71] & b[41])^(a[70] & b[42])^(a[69] & b[43])^(a[68] & b[44])^(a[67] & b[45])^(a[66] & b[46])^(a[65] & b[47])^(a[64] & b[48])^(a[63] & b[49])^(a[62] & b[50])^(a[61] & b[51])^(a[60] & b[52])^(a[59] & b[53])^(a[58] & b[54])^(a[57] & b[55])^(a[56] & b[56])^(a[55] & b[57])^(a[54] & b[58])^(a[53] & b[59])^(a[52] & b[60])^(a[51] & b[61])^(a[50] & b[62])^(a[49] & b[63])^(a[48] & b[64])^(a[47] & b[65])^(a[46] & b[66])^(a[45] & b[67])^(a[44] & b[68])^(a[43] & b[69])^(a[42] & b[70])^(a[41] & b[71])^(a[40] & b[72])^(a[39] & b[73])^(a[38] & b[74])^(a[37] & b[75])^(a[36] & b[76])^(a[35] & b[77])^(a[34] & b[78])^(a[33] & b[79])^(a[32] & b[80])^(a[31] & b[81])^(a[30] & b[82])^(a[29] & b[83])^(a[28] & b[84])^(a[27] & b[85])^(a[26] & b[86])^(a[25] & b[87])^(a[24] & b[88])^(a[23] & b[89])^(a[22] & b[90])^(a[21] & b[91])^(a[20] & b[92])^(a[19] & b[93])^(a[18] & b[94])^(a[17] & b[95])^(a[16] & b[96])^(a[15] & b[97])^(a[14] & b[98])^(a[13] & b[99])^(a[12] & b[100])^(a[11] & b[101])^(a[10] & b[102])^(a[9] & b[103])^(a[8] & b[104])^(a[7] & b[105])^(a[6] & b[106])^(a[5] & b[107])^(a[4] & b[108])^(a[3] & b[109])^(a[2] & b[110])^(a[1] & b[111])^(a[0] & b[112]);
assign y[113] = (a[113] & b[0])^(a[112] & b[1])^(a[111] & b[2])^(a[110] & b[3])^(a[109] & b[4])^(a[108] & b[5])^(a[107] & b[6])^(a[106] & b[7])^(a[105] & b[8])^(a[104] & b[9])^(a[103] & b[10])^(a[102] & b[11])^(a[101] & b[12])^(a[100] & b[13])^(a[99] & b[14])^(a[98] & b[15])^(a[97] & b[16])^(a[96] & b[17])^(a[95] & b[18])^(a[94] & b[19])^(a[93] & b[20])^(a[92] & b[21])^(a[91] & b[22])^(a[90] & b[23])^(a[89] & b[24])^(a[88] & b[25])^(a[87] & b[26])^(a[86] & b[27])^(a[85] & b[28])^(a[84] & b[29])^(a[83] & b[30])^(a[82] & b[31])^(a[81] & b[32])^(a[80] & b[33])^(a[79] & b[34])^(a[78] & b[35])^(a[77] & b[36])^(a[76] & b[37])^(a[75] & b[38])^(a[74] & b[39])^(a[73] & b[40])^(a[72] & b[41])^(a[71] & b[42])^(a[70] & b[43])^(a[69] & b[44])^(a[68] & b[45])^(a[67] & b[46])^(a[66] & b[47])^(a[65] & b[48])^(a[64] & b[49])^(a[63] & b[50])^(a[62] & b[51])^(a[61] & b[52])^(a[60] & b[53])^(a[59] & b[54])^(a[58] & b[55])^(a[57] & b[56])^(a[56] & b[57])^(a[55] & b[58])^(a[54] & b[59])^(a[53] & b[60])^(a[52] & b[61])^(a[51] & b[62])^(a[50] & b[63])^(a[49] & b[64])^(a[48] & b[65])^(a[47] & b[66])^(a[46] & b[67])^(a[45] & b[68])^(a[44] & b[69])^(a[43] & b[70])^(a[42] & b[71])^(a[41] & b[72])^(a[40] & b[73])^(a[39] & b[74])^(a[38] & b[75])^(a[37] & b[76])^(a[36] & b[77])^(a[35] & b[78])^(a[34] & b[79])^(a[33] & b[80])^(a[32] & b[81])^(a[31] & b[82])^(a[30] & b[83])^(a[29] & b[84])^(a[28] & b[85])^(a[27] & b[86])^(a[26] & b[87])^(a[25] & b[88])^(a[24] & b[89])^(a[23] & b[90])^(a[22] & b[91])^(a[21] & b[92])^(a[20] & b[93])^(a[19] & b[94])^(a[18] & b[95])^(a[17] & b[96])^(a[16] & b[97])^(a[15] & b[98])^(a[14] & b[99])^(a[13] & b[100])^(a[12] & b[101])^(a[11] & b[102])^(a[10] & b[103])^(a[9] & b[104])^(a[8] & b[105])^(a[7] & b[106])^(a[6] & b[107])^(a[5] & b[108])^(a[4] & b[109])^(a[3] & b[110])^(a[2] & b[111])^(a[1] & b[112])^(a[0] & b[113]);
assign y[114] = (a[114] & b[0])^(a[113] & b[1])^(a[112] & b[2])^(a[111] & b[3])^(a[110] & b[4])^(a[109] & b[5])^(a[108] & b[6])^(a[107] & b[7])^(a[106] & b[8])^(a[105] & b[9])^(a[104] & b[10])^(a[103] & b[11])^(a[102] & b[12])^(a[101] & b[13])^(a[100] & b[14])^(a[99] & b[15])^(a[98] & b[16])^(a[97] & b[17])^(a[96] & b[18])^(a[95] & b[19])^(a[94] & b[20])^(a[93] & b[21])^(a[92] & b[22])^(a[91] & b[23])^(a[90] & b[24])^(a[89] & b[25])^(a[88] & b[26])^(a[87] & b[27])^(a[86] & b[28])^(a[85] & b[29])^(a[84] & b[30])^(a[83] & b[31])^(a[82] & b[32])^(a[81] & b[33])^(a[80] & b[34])^(a[79] & b[35])^(a[78] & b[36])^(a[77] & b[37])^(a[76] & b[38])^(a[75] & b[39])^(a[74] & b[40])^(a[73] & b[41])^(a[72] & b[42])^(a[71] & b[43])^(a[70] & b[44])^(a[69] & b[45])^(a[68] & b[46])^(a[67] & b[47])^(a[66] & b[48])^(a[65] & b[49])^(a[64] & b[50])^(a[63] & b[51])^(a[62] & b[52])^(a[61] & b[53])^(a[60] & b[54])^(a[59] & b[55])^(a[58] & b[56])^(a[57] & b[57])^(a[56] & b[58])^(a[55] & b[59])^(a[54] & b[60])^(a[53] & b[61])^(a[52] & b[62])^(a[51] & b[63])^(a[50] & b[64])^(a[49] & b[65])^(a[48] & b[66])^(a[47] & b[67])^(a[46] & b[68])^(a[45] & b[69])^(a[44] & b[70])^(a[43] & b[71])^(a[42] & b[72])^(a[41] & b[73])^(a[40] & b[74])^(a[39] & b[75])^(a[38] & b[76])^(a[37] & b[77])^(a[36] & b[78])^(a[35] & b[79])^(a[34] & b[80])^(a[33] & b[81])^(a[32] & b[82])^(a[31] & b[83])^(a[30] & b[84])^(a[29] & b[85])^(a[28] & b[86])^(a[27] & b[87])^(a[26] & b[88])^(a[25] & b[89])^(a[24] & b[90])^(a[23] & b[91])^(a[22] & b[92])^(a[21] & b[93])^(a[20] & b[94])^(a[19] & b[95])^(a[18] & b[96])^(a[17] & b[97])^(a[16] & b[98])^(a[15] & b[99])^(a[14] & b[100])^(a[13] & b[101])^(a[12] & b[102])^(a[11] & b[103])^(a[10] & b[104])^(a[9] & b[105])^(a[8] & b[106])^(a[7] & b[107])^(a[6] & b[108])^(a[5] & b[109])^(a[4] & b[110])^(a[3] & b[111])^(a[2] & b[112])^(a[1] & b[113])^(a[0] & b[114]);
assign y[115] = (a[115] & b[0])^(a[114] & b[1])^(a[113] & b[2])^(a[112] & b[3])^(a[111] & b[4])^(a[110] & b[5])^(a[109] & b[6])^(a[108] & b[7])^(a[107] & b[8])^(a[106] & b[9])^(a[105] & b[10])^(a[104] & b[11])^(a[103] & b[12])^(a[102] & b[13])^(a[101] & b[14])^(a[100] & b[15])^(a[99] & b[16])^(a[98] & b[17])^(a[97] & b[18])^(a[96] & b[19])^(a[95] & b[20])^(a[94] & b[21])^(a[93] & b[22])^(a[92] & b[23])^(a[91] & b[24])^(a[90] & b[25])^(a[89] & b[26])^(a[88] & b[27])^(a[87] & b[28])^(a[86] & b[29])^(a[85] & b[30])^(a[84] & b[31])^(a[83] & b[32])^(a[82] & b[33])^(a[81] & b[34])^(a[80] & b[35])^(a[79] & b[36])^(a[78] & b[37])^(a[77] & b[38])^(a[76] & b[39])^(a[75] & b[40])^(a[74] & b[41])^(a[73] & b[42])^(a[72] & b[43])^(a[71] & b[44])^(a[70] & b[45])^(a[69] & b[46])^(a[68] & b[47])^(a[67] & b[48])^(a[66] & b[49])^(a[65] & b[50])^(a[64] & b[51])^(a[63] & b[52])^(a[62] & b[53])^(a[61] & b[54])^(a[60] & b[55])^(a[59] & b[56])^(a[58] & b[57])^(a[57] & b[58])^(a[56] & b[59])^(a[55] & b[60])^(a[54] & b[61])^(a[53] & b[62])^(a[52] & b[63])^(a[51] & b[64])^(a[50] & b[65])^(a[49] & b[66])^(a[48] & b[67])^(a[47] & b[68])^(a[46] & b[69])^(a[45] & b[70])^(a[44] & b[71])^(a[43] & b[72])^(a[42] & b[73])^(a[41] & b[74])^(a[40] & b[75])^(a[39] & b[76])^(a[38] & b[77])^(a[37] & b[78])^(a[36] & b[79])^(a[35] & b[80])^(a[34] & b[81])^(a[33] & b[82])^(a[32] & b[83])^(a[31] & b[84])^(a[30] & b[85])^(a[29] & b[86])^(a[28] & b[87])^(a[27] & b[88])^(a[26] & b[89])^(a[25] & b[90])^(a[24] & b[91])^(a[23] & b[92])^(a[22] & b[93])^(a[21] & b[94])^(a[20] & b[95])^(a[19] & b[96])^(a[18] & b[97])^(a[17] & b[98])^(a[16] & b[99])^(a[15] & b[100])^(a[14] & b[101])^(a[13] & b[102])^(a[12] & b[103])^(a[11] & b[104])^(a[10] & b[105])^(a[9] & b[106])^(a[8] & b[107])^(a[7] & b[108])^(a[6] & b[109])^(a[5] & b[110])^(a[4] & b[111])^(a[3] & b[112])^(a[2] & b[113])^(a[1] & b[114])^(a[0] & b[115]);
assign y[116] = (a[116] & b[0])^(a[115] & b[1])^(a[114] & b[2])^(a[113] & b[3])^(a[112] & b[4])^(a[111] & b[5])^(a[110] & b[6])^(a[109] & b[7])^(a[108] & b[8])^(a[107] & b[9])^(a[106] & b[10])^(a[105] & b[11])^(a[104] & b[12])^(a[103] & b[13])^(a[102] & b[14])^(a[101] & b[15])^(a[100] & b[16])^(a[99] & b[17])^(a[98] & b[18])^(a[97] & b[19])^(a[96] & b[20])^(a[95] & b[21])^(a[94] & b[22])^(a[93] & b[23])^(a[92] & b[24])^(a[91] & b[25])^(a[90] & b[26])^(a[89] & b[27])^(a[88] & b[28])^(a[87] & b[29])^(a[86] & b[30])^(a[85] & b[31])^(a[84] & b[32])^(a[83] & b[33])^(a[82] & b[34])^(a[81] & b[35])^(a[80] & b[36])^(a[79] & b[37])^(a[78] & b[38])^(a[77] & b[39])^(a[76] & b[40])^(a[75] & b[41])^(a[74] & b[42])^(a[73] & b[43])^(a[72] & b[44])^(a[71] & b[45])^(a[70] & b[46])^(a[69] & b[47])^(a[68] & b[48])^(a[67] & b[49])^(a[66] & b[50])^(a[65] & b[51])^(a[64] & b[52])^(a[63] & b[53])^(a[62] & b[54])^(a[61] & b[55])^(a[60] & b[56])^(a[59] & b[57])^(a[58] & b[58])^(a[57] & b[59])^(a[56] & b[60])^(a[55] & b[61])^(a[54] & b[62])^(a[53] & b[63])^(a[52] & b[64])^(a[51] & b[65])^(a[50] & b[66])^(a[49] & b[67])^(a[48] & b[68])^(a[47] & b[69])^(a[46] & b[70])^(a[45] & b[71])^(a[44] & b[72])^(a[43] & b[73])^(a[42] & b[74])^(a[41] & b[75])^(a[40] & b[76])^(a[39] & b[77])^(a[38] & b[78])^(a[37] & b[79])^(a[36] & b[80])^(a[35] & b[81])^(a[34] & b[82])^(a[33] & b[83])^(a[32] & b[84])^(a[31] & b[85])^(a[30] & b[86])^(a[29] & b[87])^(a[28] & b[88])^(a[27] & b[89])^(a[26] & b[90])^(a[25] & b[91])^(a[24] & b[92])^(a[23] & b[93])^(a[22] & b[94])^(a[21] & b[95])^(a[20] & b[96])^(a[19] & b[97])^(a[18] & b[98])^(a[17] & b[99])^(a[16] & b[100])^(a[15] & b[101])^(a[14] & b[102])^(a[13] & b[103])^(a[12] & b[104])^(a[11] & b[105])^(a[10] & b[106])^(a[9] & b[107])^(a[8] & b[108])^(a[7] & b[109])^(a[6] & b[110])^(a[5] & b[111])^(a[4] & b[112])^(a[3] & b[113])^(a[2] & b[114])^(a[1] & b[115])^(a[0] & b[116]);
assign y[117] = (a[117] & b[0])^(a[116] & b[1])^(a[115] & b[2])^(a[114] & b[3])^(a[113] & b[4])^(a[112] & b[5])^(a[111] & b[6])^(a[110] & b[7])^(a[109] & b[8])^(a[108] & b[9])^(a[107] & b[10])^(a[106] & b[11])^(a[105] & b[12])^(a[104] & b[13])^(a[103] & b[14])^(a[102] & b[15])^(a[101] & b[16])^(a[100] & b[17])^(a[99] & b[18])^(a[98] & b[19])^(a[97] & b[20])^(a[96] & b[21])^(a[95] & b[22])^(a[94] & b[23])^(a[93] & b[24])^(a[92] & b[25])^(a[91] & b[26])^(a[90] & b[27])^(a[89] & b[28])^(a[88] & b[29])^(a[87] & b[30])^(a[86] & b[31])^(a[85] & b[32])^(a[84] & b[33])^(a[83] & b[34])^(a[82] & b[35])^(a[81] & b[36])^(a[80] & b[37])^(a[79] & b[38])^(a[78] & b[39])^(a[77] & b[40])^(a[76] & b[41])^(a[75] & b[42])^(a[74] & b[43])^(a[73] & b[44])^(a[72] & b[45])^(a[71] & b[46])^(a[70] & b[47])^(a[69] & b[48])^(a[68] & b[49])^(a[67] & b[50])^(a[66] & b[51])^(a[65] & b[52])^(a[64] & b[53])^(a[63] & b[54])^(a[62] & b[55])^(a[61] & b[56])^(a[60] & b[57])^(a[59] & b[58])^(a[58] & b[59])^(a[57] & b[60])^(a[56] & b[61])^(a[55] & b[62])^(a[54] & b[63])^(a[53] & b[64])^(a[52] & b[65])^(a[51] & b[66])^(a[50] & b[67])^(a[49] & b[68])^(a[48] & b[69])^(a[47] & b[70])^(a[46] & b[71])^(a[45] & b[72])^(a[44] & b[73])^(a[43] & b[74])^(a[42] & b[75])^(a[41] & b[76])^(a[40] & b[77])^(a[39] & b[78])^(a[38] & b[79])^(a[37] & b[80])^(a[36] & b[81])^(a[35] & b[82])^(a[34] & b[83])^(a[33] & b[84])^(a[32] & b[85])^(a[31] & b[86])^(a[30] & b[87])^(a[29] & b[88])^(a[28] & b[89])^(a[27] & b[90])^(a[26] & b[91])^(a[25] & b[92])^(a[24] & b[93])^(a[23] & b[94])^(a[22] & b[95])^(a[21] & b[96])^(a[20] & b[97])^(a[19] & b[98])^(a[18] & b[99])^(a[17] & b[100])^(a[16] & b[101])^(a[15] & b[102])^(a[14] & b[103])^(a[13] & b[104])^(a[12] & b[105])^(a[11] & b[106])^(a[10] & b[107])^(a[9] & b[108])^(a[8] & b[109])^(a[7] & b[110])^(a[6] & b[111])^(a[5] & b[112])^(a[4] & b[113])^(a[3] & b[114])^(a[2] & b[115])^(a[1] & b[116])^(a[0] & b[117]);
assign y[118] = (a[118] & b[0])^(a[117] & b[1])^(a[116] & b[2])^(a[115] & b[3])^(a[114] & b[4])^(a[113] & b[5])^(a[112] & b[6])^(a[111] & b[7])^(a[110] & b[8])^(a[109] & b[9])^(a[108] & b[10])^(a[107] & b[11])^(a[106] & b[12])^(a[105] & b[13])^(a[104] & b[14])^(a[103] & b[15])^(a[102] & b[16])^(a[101] & b[17])^(a[100] & b[18])^(a[99] & b[19])^(a[98] & b[20])^(a[97] & b[21])^(a[96] & b[22])^(a[95] & b[23])^(a[94] & b[24])^(a[93] & b[25])^(a[92] & b[26])^(a[91] & b[27])^(a[90] & b[28])^(a[89] & b[29])^(a[88] & b[30])^(a[87] & b[31])^(a[86] & b[32])^(a[85] & b[33])^(a[84] & b[34])^(a[83] & b[35])^(a[82] & b[36])^(a[81] & b[37])^(a[80] & b[38])^(a[79] & b[39])^(a[78] & b[40])^(a[77] & b[41])^(a[76] & b[42])^(a[75] & b[43])^(a[74] & b[44])^(a[73] & b[45])^(a[72] & b[46])^(a[71] & b[47])^(a[70] & b[48])^(a[69] & b[49])^(a[68] & b[50])^(a[67] & b[51])^(a[66] & b[52])^(a[65] & b[53])^(a[64] & b[54])^(a[63] & b[55])^(a[62] & b[56])^(a[61] & b[57])^(a[60] & b[58])^(a[59] & b[59])^(a[58] & b[60])^(a[57] & b[61])^(a[56] & b[62])^(a[55] & b[63])^(a[54] & b[64])^(a[53] & b[65])^(a[52] & b[66])^(a[51] & b[67])^(a[50] & b[68])^(a[49] & b[69])^(a[48] & b[70])^(a[47] & b[71])^(a[46] & b[72])^(a[45] & b[73])^(a[44] & b[74])^(a[43] & b[75])^(a[42] & b[76])^(a[41] & b[77])^(a[40] & b[78])^(a[39] & b[79])^(a[38] & b[80])^(a[37] & b[81])^(a[36] & b[82])^(a[35] & b[83])^(a[34] & b[84])^(a[33] & b[85])^(a[32] & b[86])^(a[31] & b[87])^(a[30] & b[88])^(a[29] & b[89])^(a[28] & b[90])^(a[27] & b[91])^(a[26] & b[92])^(a[25] & b[93])^(a[24] & b[94])^(a[23] & b[95])^(a[22] & b[96])^(a[21] & b[97])^(a[20] & b[98])^(a[19] & b[99])^(a[18] & b[100])^(a[17] & b[101])^(a[16] & b[102])^(a[15] & b[103])^(a[14] & b[104])^(a[13] & b[105])^(a[12] & b[106])^(a[11] & b[107])^(a[10] & b[108])^(a[9] & b[109])^(a[8] & b[110])^(a[7] & b[111])^(a[6] & b[112])^(a[5] & b[113])^(a[4] & b[114])^(a[3] & b[115])^(a[2] & b[116])^(a[1] & b[117])^(a[0] & b[118]);
assign y[119] = (a[119] & b[0])^(a[118] & b[1])^(a[117] & b[2])^(a[116] & b[3])^(a[115] & b[4])^(a[114] & b[5])^(a[113] & b[6])^(a[112] & b[7])^(a[111] & b[8])^(a[110] & b[9])^(a[109] & b[10])^(a[108] & b[11])^(a[107] & b[12])^(a[106] & b[13])^(a[105] & b[14])^(a[104] & b[15])^(a[103] & b[16])^(a[102] & b[17])^(a[101] & b[18])^(a[100] & b[19])^(a[99] & b[20])^(a[98] & b[21])^(a[97] & b[22])^(a[96] & b[23])^(a[95] & b[24])^(a[94] & b[25])^(a[93] & b[26])^(a[92] & b[27])^(a[91] & b[28])^(a[90] & b[29])^(a[89] & b[30])^(a[88] & b[31])^(a[87] & b[32])^(a[86] & b[33])^(a[85] & b[34])^(a[84] & b[35])^(a[83] & b[36])^(a[82] & b[37])^(a[81] & b[38])^(a[80] & b[39])^(a[79] & b[40])^(a[78] & b[41])^(a[77] & b[42])^(a[76] & b[43])^(a[75] & b[44])^(a[74] & b[45])^(a[73] & b[46])^(a[72] & b[47])^(a[71] & b[48])^(a[70] & b[49])^(a[69] & b[50])^(a[68] & b[51])^(a[67] & b[52])^(a[66] & b[53])^(a[65] & b[54])^(a[64] & b[55])^(a[63] & b[56])^(a[62] & b[57])^(a[61] & b[58])^(a[60] & b[59])^(a[59] & b[60])^(a[58] & b[61])^(a[57] & b[62])^(a[56] & b[63])^(a[55] & b[64])^(a[54] & b[65])^(a[53] & b[66])^(a[52] & b[67])^(a[51] & b[68])^(a[50] & b[69])^(a[49] & b[70])^(a[48] & b[71])^(a[47] & b[72])^(a[46] & b[73])^(a[45] & b[74])^(a[44] & b[75])^(a[43] & b[76])^(a[42] & b[77])^(a[41] & b[78])^(a[40] & b[79])^(a[39] & b[80])^(a[38] & b[81])^(a[37] & b[82])^(a[36] & b[83])^(a[35] & b[84])^(a[34] & b[85])^(a[33] & b[86])^(a[32] & b[87])^(a[31] & b[88])^(a[30] & b[89])^(a[29] & b[90])^(a[28] & b[91])^(a[27] & b[92])^(a[26] & b[93])^(a[25] & b[94])^(a[24] & b[95])^(a[23] & b[96])^(a[22] & b[97])^(a[21] & b[98])^(a[20] & b[99])^(a[19] & b[100])^(a[18] & b[101])^(a[17] & b[102])^(a[16] & b[103])^(a[15] & b[104])^(a[14] & b[105])^(a[13] & b[106])^(a[12] & b[107])^(a[11] & b[108])^(a[10] & b[109])^(a[9] & b[110])^(a[8] & b[111])^(a[7] & b[112])^(a[6] & b[113])^(a[5] & b[114])^(a[4] & b[115])^(a[3] & b[116])^(a[2] & b[117])^(a[1] & b[118])^(a[0] & b[119]);
assign y[120] = (a[120] & b[0])^(a[119] & b[1])^(a[118] & b[2])^(a[117] & b[3])^(a[116] & b[4])^(a[115] & b[5])^(a[114] & b[6])^(a[113] & b[7])^(a[112] & b[8])^(a[111] & b[9])^(a[110] & b[10])^(a[109] & b[11])^(a[108] & b[12])^(a[107] & b[13])^(a[106] & b[14])^(a[105] & b[15])^(a[104] & b[16])^(a[103] & b[17])^(a[102] & b[18])^(a[101] & b[19])^(a[100] & b[20])^(a[99] & b[21])^(a[98] & b[22])^(a[97] & b[23])^(a[96] & b[24])^(a[95] & b[25])^(a[94] & b[26])^(a[93] & b[27])^(a[92] & b[28])^(a[91] & b[29])^(a[90] & b[30])^(a[89] & b[31])^(a[88] & b[32])^(a[87] & b[33])^(a[86] & b[34])^(a[85] & b[35])^(a[84] & b[36])^(a[83] & b[37])^(a[82] & b[38])^(a[81] & b[39])^(a[80] & b[40])^(a[79] & b[41])^(a[78] & b[42])^(a[77] & b[43])^(a[76] & b[44])^(a[75] & b[45])^(a[74] & b[46])^(a[73] & b[47])^(a[72] & b[48])^(a[71] & b[49])^(a[70] & b[50])^(a[69] & b[51])^(a[68] & b[52])^(a[67] & b[53])^(a[66] & b[54])^(a[65] & b[55])^(a[64] & b[56])^(a[63] & b[57])^(a[62] & b[58])^(a[61] & b[59])^(a[60] & b[60])^(a[59] & b[61])^(a[58] & b[62])^(a[57] & b[63])^(a[56] & b[64])^(a[55] & b[65])^(a[54] & b[66])^(a[53] & b[67])^(a[52] & b[68])^(a[51] & b[69])^(a[50] & b[70])^(a[49] & b[71])^(a[48] & b[72])^(a[47] & b[73])^(a[46] & b[74])^(a[45] & b[75])^(a[44] & b[76])^(a[43] & b[77])^(a[42] & b[78])^(a[41] & b[79])^(a[40] & b[80])^(a[39] & b[81])^(a[38] & b[82])^(a[37] & b[83])^(a[36] & b[84])^(a[35] & b[85])^(a[34] & b[86])^(a[33] & b[87])^(a[32] & b[88])^(a[31] & b[89])^(a[30] & b[90])^(a[29] & b[91])^(a[28] & b[92])^(a[27] & b[93])^(a[26] & b[94])^(a[25] & b[95])^(a[24] & b[96])^(a[23] & b[97])^(a[22] & b[98])^(a[21] & b[99])^(a[20] & b[100])^(a[19] & b[101])^(a[18] & b[102])^(a[17] & b[103])^(a[16] & b[104])^(a[15] & b[105])^(a[14] & b[106])^(a[13] & b[107])^(a[12] & b[108])^(a[11] & b[109])^(a[10] & b[110])^(a[9] & b[111])^(a[8] & b[112])^(a[7] & b[113])^(a[6] & b[114])^(a[5] & b[115])^(a[4] & b[116])^(a[3] & b[117])^(a[2] & b[118])^(a[1] & b[119])^(a[0] & b[120]);
assign y[121] = (a[121] & b[0])^(a[120] & b[1])^(a[119] & b[2])^(a[118] & b[3])^(a[117] & b[4])^(a[116] & b[5])^(a[115] & b[6])^(a[114] & b[7])^(a[113] & b[8])^(a[112] & b[9])^(a[111] & b[10])^(a[110] & b[11])^(a[109] & b[12])^(a[108] & b[13])^(a[107] & b[14])^(a[106] & b[15])^(a[105] & b[16])^(a[104] & b[17])^(a[103] & b[18])^(a[102] & b[19])^(a[101] & b[20])^(a[100] & b[21])^(a[99] & b[22])^(a[98] & b[23])^(a[97] & b[24])^(a[96] & b[25])^(a[95] & b[26])^(a[94] & b[27])^(a[93] & b[28])^(a[92] & b[29])^(a[91] & b[30])^(a[90] & b[31])^(a[89] & b[32])^(a[88] & b[33])^(a[87] & b[34])^(a[86] & b[35])^(a[85] & b[36])^(a[84] & b[37])^(a[83] & b[38])^(a[82] & b[39])^(a[81] & b[40])^(a[80] & b[41])^(a[79] & b[42])^(a[78] & b[43])^(a[77] & b[44])^(a[76] & b[45])^(a[75] & b[46])^(a[74] & b[47])^(a[73] & b[48])^(a[72] & b[49])^(a[71] & b[50])^(a[70] & b[51])^(a[69] & b[52])^(a[68] & b[53])^(a[67] & b[54])^(a[66] & b[55])^(a[65] & b[56])^(a[64] & b[57])^(a[63] & b[58])^(a[62] & b[59])^(a[61] & b[60])^(a[60] & b[61])^(a[59] & b[62])^(a[58] & b[63])^(a[57] & b[64])^(a[56] & b[65])^(a[55] & b[66])^(a[54] & b[67])^(a[53] & b[68])^(a[52] & b[69])^(a[51] & b[70])^(a[50] & b[71])^(a[49] & b[72])^(a[48] & b[73])^(a[47] & b[74])^(a[46] & b[75])^(a[45] & b[76])^(a[44] & b[77])^(a[43] & b[78])^(a[42] & b[79])^(a[41] & b[80])^(a[40] & b[81])^(a[39] & b[82])^(a[38] & b[83])^(a[37] & b[84])^(a[36] & b[85])^(a[35] & b[86])^(a[34] & b[87])^(a[33] & b[88])^(a[32] & b[89])^(a[31] & b[90])^(a[30] & b[91])^(a[29] & b[92])^(a[28] & b[93])^(a[27] & b[94])^(a[26] & b[95])^(a[25] & b[96])^(a[24] & b[97])^(a[23] & b[98])^(a[22] & b[99])^(a[21] & b[100])^(a[20] & b[101])^(a[19] & b[102])^(a[18] & b[103])^(a[17] & b[104])^(a[16] & b[105])^(a[15] & b[106])^(a[14] & b[107])^(a[13] & b[108])^(a[12] & b[109])^(a[11] & b[110])^(a[10] & b[111])^(a[9] & b[112])^(a[8] & b[113])^(a[7] & b[114])^(a[6] & b[115])^(a[5] & b[116])^(a[4] & b[117])^(a[3] & b[118])^(a[2] & b[119])^(a[1] & b[120])^(a[0] & b[121]);
assign y[122] = (a[122] & b[0])^(a[121] & b[1])^(a[120] & b[2])^(a[119] & b[3])^(a[118] & b[4])^(a[117] & b[5])^(a[116] & b[6])^(a[115] & b[7])^(a[114] & b[8])^(a[113] & b[9])^(a[112] & b[10])^(a[111] & b[11])^(a[110] & b[12])^(a[109] & b[13])^(a[108] & b[14])^(a[107] & b[15])^(a[106] & b[16])^(a[105] & b[17])^(a[104] & b[18])^(a[103] & b[19])^(a[102] & b[20])^(a[101] & b[21])^(a[100] & b[22])^(a[99] & b[23])^(a[98] & b[24])^(a[97] & b[25])^(a[96] & b[26])^(a[95] & b[27])^(a[94] & b[28])^(a[93] & b[29])^(a[92] & b[30])^(a[91] & b[31])^(a[90] & b[32])^(a[89] & b[33])^(a[88] & b[34])^(a[87] & b[35])^(a[86] & b[36])^(a[85] & b[37])^(a[84] & b[38])^(a[83] & b[39])^(a[82] & b[40])^(a[81] & b[41])^(a[80] & b[42])^(a[79] & b[43])^(a[78] & b[44])^(a[77] & b[45])^(a[76] & b[46])^(a[75] & b[47])^(a[74] & b[48])^(a[73] & b[49])^(a[72] & b[50])^(a[71] & b[51])^(a[70] & b[52])^(a[69] & b[53])^(a[68] & b[54])^(a[67] & b[55])^(a[66] & b[56])^(a[65] & b[57])^(a[64] & b[58])^(a[63] & b[59])^(a[62] & b[60])^(a[61] & b[61])^(a[60] & b[62])^(a[59] & b[63])^(a[58] & b[64])^(a[57] & b[65])^(a[56] & b[66])^(a[55] & b[67])^(a[54] & b[68])^(a[53] & b[69])^(a[52] & b[70])^(a[51] & b[71])^(a[50] & b[72])^(a[49] & b[73])^(a[48] & b[74])^(a[47] & b[75])^(a[46] & b[76])^(a[45] & b[77])^(a[44] & b[78])^(a[43] & b[79])^(a[42] & b[80])^(a[41] & b[81])^(a[40] & b[82])^(a[39] & b[83])^(a[38] & b[84])^(a[37] & b[85])^(a[36] & b[86])^(a[35] & b[87])^(a[34] & b[88])^(a[33] & b[89])^(a[32] & b[90])^(a[31] & b[91])^(a[30] & b[92])^(a[29] & b[93])^(a[28] & b[94])^(a[27] & b[95])^(a[26] & b[96])^(a[25] & b[97])^(a[24] & b[98])^(a[23] & b[99])^(a[22] & b[100])^(a[21] & b[101])^(a[20] & b[102])^(a[19] & b[103])^(a[18] & b[104])^(a[17] & b[105])^(a[16] & b[106])^(a[15] & b[107])^(a[14] & b[108])^(a[13] & b[109])^(a[12] & b[110])^(a[11] & b[111])^(a[10] & b[112])^(a[9] & b[113])^(a[8] & b[114])^(a[7] & b[115])^(a[6] & b[116])^(a[5] & b[117])^(a[4] & b[118])^(a[3] & b[119])^(a[2] & b[120])^(a[1] & b[121])^(a[0] & b[122]);
assign y[123] = (a[123] & b[0])^(a[122] & b[1])^(a[121] & b[2])^(a[120] & b[3])^(a[119] & b[4])^(a[118] & b[5])^(a[117] & b[6])^(a[116] & b[7])^(a[115] & b[8])^(a[114] & b[9])^(a[113] & b[10])^(a[112] & b[11])^(a[111] & b[12])^(a[110] & b[13])^(a[109] & b[14])^(a[108] & b[15])^(a[107] & b[16])^(a[106] & b[17])^(a[105] & b[18])^(a[104] & b[19])^(a[103] & b[20])^(a[102] & b[21])^(a[101] & b[22])^(a[100] & b[23])^(a[99] & b[24])^(a[98] & b[25])^(a[97] & b[26])^(a[96] & b[27])^(a[95] & b[28])^(a[94] & b[29])^(a[93] & b[30])^(a[92] & b[31])^(a[91] & b[32])^(a[90] & b[33])^(a[89] & b[34])^(a[88] & b[35])^(a[87] & b[36])^(a[86] & b[37])^(a[85] & b[38])^(a[84] & b[39])^(a[83] & b[40])^(a[82] & b[41])^(a[81] & b[42])^(a[80] & b[43])^(a[79] & b[44])^(a[78] & b[45])^(a[77] & b[46])^(a[76] & b[47])^(a[75] & b[48])^(a[74] & b[49])^(a[73] & b[50])^(a[72] & b[51])^(a[71] & b[52])^(a[70] & b[53])^(a[69] & b[54])^(a[68] & b[55])^(a[67] & b[56])^(a[66] & b[57])^(a[65] & b[58])^(a[64] & b[59])^(a[63] & b[60])^(a[62] & b[61])^(a[61] & b[62])^(a[60] & b[63])^(a[59] & b[64])^(a[58] & b[65])^(a[57] & b[66])^(a[56] & b[67])^(a[55] & b[68])^(a[54] & b[69])^(a[53] & b[70])^(a[52] & b[71])^(a[51] & b[72])^(a[50] & b[73])^(a[49] & b[74])^(a[48] & b[75])^(a[47] & b[76])^(a[46] & b[77])^(a[45] & b[78])^(a[44] & b[79])^(a[43] & b[80])^(a[42] & b[81])^(a[41] & b[82])^(a[40] & b[83])^(a[39] & b[84])^(a[38] & b[85])^(a[37] & b[86])^(a[36] & b[87])^(a[35] & b[88])^(a[34] & b[89])^(a[33] & b[90])^(a[32] & b[91])^(a[31] & b[92])^(a[30] & b[93])^(a[29] & b[94])^(a[28] & b[95])^(a[27] & b[96])^(a[26] & b[97])^(a[25] & b[98])^(a[24] & b[99])^(a[23] & b[100])^(a[22] & b[101])^(a[21] & b[102])^(a[20] & b[103])^(a[19] & b[104])^(a[18] & b[105])^(a[17] & b[106])^(a[16] & b[107])^(a[15] & b[108])^(a[14] & b[109])^(a[13] & b[110])^(a[12] & b[111])^(a[11] & b[112])^(a[10] & b[113])^(a[9] & b[114])^(a[8] & b[115])^(a[7] & b[116])^(a[6] & b[117])^(a[5] & b[118])^(a[4] & b[119])^(a[3] & b[120])^(a[2] & b[121])^(a[1] & b[122])^(a[0] & b[123]);
assign y[124] = (a[124] & b[0])^(a[123] & b[1])^(a[122] & b[2])^(a[121] & b[3])^(a[120] & b[4])^(a[119] & b[5])^(a[118] & b[6])^(a[117] & b[7])^(a[116] & b[8])^(a[115] & b[9])^(a[114] & b[10])^(a[113] & b[11])^(a[112] & b[12])^(a[111] & b[13])^(a[110] & b[14])^(a[109] & b[15])^(a[108] & b[16])^(a[107] & b[17])^(a[106] & b[18])^(a[105] & b[19])^(a[104] & b[20])^(a[103] & b[21])^(a[102] & b[22])^(a[101] & b[23])^(a[100] & b[24])^(a[99] & b[25])^(a[98] & b[26])^(a[97] & b[27])^(a[96] & b[28])^(a[95] & b[29])^(a[94] & b[30])^(a[93] & b[31])^(a[92] & b[32])^(a[91] & b[33])^(a[90] & b[34])^(a[89] & b[35])^(a[88] & b[36])^(a[87] & b[37])^(a[86] & b[38])^(a[85] & b[39])^(a[84] & b[40])^(a[83] & b[41])^(a[82] & b[42])^(a[81] & b[43])^(a[80] & b[44])^(a[79] & b[45])^(a[78] & b[46])^(a[77] & b[47])^(a[76] & b[48])^(a[75] & b[49])^(a[74] & b[50])^(a[73] & b[51])^(a[72] & b[52])^(a[71] & b[53])^(a[70] & b[54])^(a[69] & b[55])^(a[68] & b[56])^(a[67] & b[57])^(a[66] & b[58])^(a[65] & b[59])^(a[64] & b[60])^(a[63] & b[61])^(a[62] & b[62])^(a[61] & b[63])^(a[60] & b[64])^(a[59] & b[65])^(a[58] & b[66])^(a[57] & b[67])^(a[56] & b[68])^(a[55] & b[69])^(a[54] & b[70])^(a[53] & b[71])^(a[52] & b[72])^(a[51] & b[73])^(a[50] & b[74])^(a[49] & b[75])^(a[48] & b[76])^(a[47] & b[77])^(a[46] & b[78])^(a[45] & b[79])^(a[44] & b[80])^(a[43] & b[81])^(a[42] & b[82])^(a[41] & b[83])^(a[40] & b[84])^(a[39] & b[85])^(a[38] & b[86])^(a[37] & b[87])^(a[36] & b[88])^(a[35] & b[89])^(a[34] & b[90])^(a[33] & b[91])^(a[32] & b[92])^(a[31] & b[93])^(a[30] & b[94])^(a[29] & b[95])^(a[28] & b[96])^(a[27] & b[97])^(a[26] & b[98])^(a[25] & b[99])^(a[24] & b[100])^(a[23] & b[101])^(a[22] & b[102])^(a[21] & b[103])^(a[20] & b[104])^(a[19] & b[105])^(a[18] & b[106])^(a[17] & b[107])^(a[16] & b[108])^(a[15] & b[109])^(a[14] & b[110])^(a[13] & b[111])^(a[12] & b[112])^(a[11] & b[113])^(a[10] & b[114])^(a[9] & b[115])^(a[8] & b[116])^(a[7] & b[117])^(a[6] & b[118])^(a[5] & b[119])^(a[4] & b[120])^(a[3] & b[121])^(a[2] & b[122])^(a[1] & b[123])^(a[0] & b[124]);
assign y[125] = (a[125] & b[0])^(a[124] & b[1])^(a[123] & b[2])^(a[122] & b[3])^(a[121] & b[4])^(a[120] & b[5])^(a[119] & b[6])^(a[118] & b[7])^(a[117] & b[8])^(a[116] & b[9])^(a[115] & b[10])^(a[114] & b[11])^(a[113] & b[12])^(a[112] & b[13])^(a[111] & b[14])^(a[110] & b[15])^(a[109] & b[16])^(a[108] & b[17])^(a[107] & b[18])^(a[106] & b[19])^(a[105] & b[20])^(a[104] & b[21])^(a[103] & b[22])^(a[102] & b[23])^(a[101] & b[24])^(a[100] & b[25])^(a[99] & b[26])^(a[98] & b[27])^(a[97] & b[28])^(a[96] & b[29])^(a[95] & b[30])^(a[94] & b[31])^(a[93] & b[32])^(a[92] & b[33])^(a[91] & b[34])^(a[90] & b[35])^(a[89] & b[36])^(a[88] & b[37])^(a[87] & b[38])^(a[86] & b[39])^(a[85] & b[40])^(a[84] & b[41])^(a[83] & b[42])^(a[82] & b[43])^(a[81] & b[44])^(a[80] & b[45])^(a[79] & b[46])^(a[78] & b[47])^(a[77] & b[48])^(a[76] & b[49])^(a[75] & b[50])^(a[74] & b[51])^(a[73] & b[52])^(a[72] & b[53])^(a[71] & b[54])^(a[70] & b[55])^(a[69] & b[56])^(a[68] & b[57])^(a[67] & b[58])^(a[66] & b[59])^(a[65] & b[60])^(a[64] & b[61])^(a[63] & b[62])^(a[62] & b[63])^(a[61] & b[64])^(a[60] & b[65])^(a[59] & b[66])^(a[58] & b[67])^(a[57] & b[68])^(a[56] & b[69])^(a[55] & b[70])^(a[54] & b[71])^(a[53] & b[72])^(a[52] & b[73])^(a[51] & b[74])^(a[50] & b[75])^(a[49] & b[76])^(a[48] & b[77])^(a[47] & b[78])^(a[46] & b[79])^(a[45] & b[80])^(a[44] & b[81])^(a[43] & b[82])^(a[42] & b[83])^(a[41] & b[84])^(a[40] & b[85])^(a[39] & b[86])^(a[38] & b[87])^(a[37] & b[88])^(a[36] & b[89])^(a[35] & b[90])^(a[34] & b[91])^(a[33] & b[92])^(a[32] & b[93])^(a[31] & b[94])^(a[30] & b[95])^(a[29] & b[96])^(a[28] & b[97])^(a[27] & b[98])^(a[26] & b[99])^(a[25] & b[100])^(a[24] & b[101])^(a[23] & b[102])^(a[22] & b[103])^(a[21] & b[104])^(a[20] & b[105])^(a[19] & b[106])^(a[18] & b[107])^(a[17] & b[108])^(a[16] & b[109])^(a[15] & b[110])^(a[14] & b[111])^(a[13] & b[112])^(a[12] & b[113])^(a[11] & b[114])^(a[10] & b[115])^(a[9] & b[116])^(a[8] & b[117])^(a[7] & b[118])^(a[6] & b[119])^(a[5] & b[120])^(a[4] & b[121])^(a[3] & b[122])^(a[2] & b[123])^(a[1] & b[124])^(a[0] & b[125]);
assign y[126] = (a[126] & b[0])^(a[125] & b[1])^(a[124] & b[2])^(a[123] & b[3])^(a[122] & b[4])^(a[121] & b[5])^(a[120] & b[6])^(a[119] & b[7])^(a[118] & b[8])^(a[117] & b[9])^(a[116] & b[10])^(a[115] & b[11])^(a[114] & b[12])^(a[113] & b[13])^(a[112] & b[14])^(a[111] & b[15])^(a[110] & b[16])^(a[109] & b[17])^(a[108] & b[18])^(a[107] & b[19])^(a[106] & b[20])^(a[105] & b[21])^(a[104] & b[22])^(a[103] & b[23])^(a[102] & b[24])^(a[101] & b[25])^(a[100] & b[26])^(a[99] & b[27])^(a[98] & b[28])^(a[97] & b[29])^(a[96] & b[30])^(a[95] & b[31])^(a[94] & b[32])^(a[93] & b[33])^(a[92] & b[34])^(a[91] & b[35])^(a[90] & b[36])^(a[89] & b[37])^(a[88] & b[38])^(a[87] & b[39])^(a[86] & b[40])^(a[85] & b[41])^(a[84] & b[42])^(a[83] & b[43])^(a[82] & b[44])^(a[81] & b[45])^(a[80] & b[46])^(a[79] & b[47])^(a[78] & b[48])^(a[77] & b[49])^(a[76] & b[50])^(a[75] & b[51])^(a[74] & b[52])^(a[73] & b[53])^(a[72] & b[54])^(a[71] & b[55])^(a[70] & b[56])^(a[69] & b[57])^(a[68] & b[58])^(a[67] & b[59])^(a[66] & b[60])^(a[65] & b[61])^(a[64] & b[62])^(a[63] & b[63])^(a[62] & b[64])^(a[61] & b[65])^(a[60] & b[66])^(a[59] & b[67])^(a[58] & b[68])^(a[57] & b[69])^(a[56] & b[70])^(a[55] & b[71])^(a[54] & b[72])^(a[53] & b[73])^(a[52] & b[74])^(a[51] & b[75])^(a[50] & b[76])^(a[49] & b[77])^(a[48] & b[78])^(a[47] & b[79])^(a[46] & b[80])^(a[45] & b[81])^(a[44] & b[82])^(a[43] & b[83])^(a[42] & b[84])^(a[41] & b[85])^(a[40] & b[86])^(a[39] & b[87])^(a[38] & b[88])^(a[37] & b[89])^(a[36] & b[90])^(a[35] & b[91])^(a[34] & b[92])^(a[33] & b[93])^(a[32] & b[94])^(a[31] & b[95])^(a[30] & b[96])^(a[29] & b[97])^(a[28] & b[98])^(a[27] & b[99])^(a[26] & b[100])^(a[25] & b[101])^(a[24] & b[102])^(a[23] & b[103])^(a[22] & b[104])^(a[21] & b[105])^(a[20] & b[106])^(a[19] & b[107])^(a[18] & b[108])^(a[17] & b[109])^(a[16] & b[110])^(a[15] & b[111])^(a[14] & b[112])^(a[13] & b[113])^(a[12] & b[114])^(a[11] & b[115])^(a[10] & b[116])^(a[9] & b[117])^(a[8] & b[118])^(a[7] & b[119])^(a[6] & b[120])^(a[5] & b[121])^(a[4] & b[122])^(a[3] & b[123])^(a[2] & b[124])^(a[1] & b[125])^(a[0] & b[126]);
assign y[127] = (a[127] & b[0])^(a[126] & b[1])^(a[125] & b[2])^(a[124] & b[3])^(a[123] & b[4])^(a[122] & b[5])^(a[121] & b[6])^(a[120] & b[7])^(a[119] & b[8])^(a[118] & b[9])^(a[117] & b[10])^(a[116] & b[11])^(a[115] & b[12])^(a[114] & b[13])^(a[113] & b[14])^(a[112] & b[15])^(a[111] & b[16])^(a[110] & b[17])^(a[109] & b[18])^(a[108] & b[19])^(a[107] & b[20])^(a[106] & b[21])^(a[105] & b[22])^(a[104] & b[23])^(a[103] & b[24])^(a[102] & b[25])^(a[101] & b[26])^(a[100] & b[27])^(a[99] & b[28])^(a[98] & b[29])^(a[97] & b[30])^(a[96] & b[31])^(a[95] & b[32])^(a[94] & b[33])^(a[93] & b[34])^(a[92] & b[35])^(a[91] & b[36])^(a[90] & b[37])^(a[89] & b[38])^(a[88] & b[39])^(a[87] & b[40])^(a[86] & b[41])^(a[85] & b[42])^(a[84] & b[43])^(a[83] & b[44])^(a[82] & b[45])^(a[81] & b[46])^(a[80] & b[47])^(a[79] & b[48])^(a[78] & b[49])^(a[77] & b[50])^(a[76] & b[51])^(a[75] & b[52])^(a[74] & b[53])^(a[73] & b[54])^(a[72] & b[55])^(a[71] & b[56])^(a[70] & b[57])^(a[69] & b[58])^(a[68] & b[59])^(a[67] & b[60])^(a[66] & b[61])^(a[65] & b[62])^(a[64] & b[63])^(a[63] & b[64])^(a[62] & b[65])^(a[61] & b[66])^(a[60] & b[67])^(a[59] & b[68])^(a[58] & b[69])^(a[57] & b[70])^(a[56] & b[71])^(a[55] & b[72])^(a[54] & b[73])^(a[53] & b[74])^(a[52] & b[75])^(a[51] & b[76])^(a[50] & b[77])^(a[49] & b[78])^(a[48] & b[79])^(a[47] & b[80])^(a[46] & b[81])^(a[45] & b[82])^(a[44] & b[83])^(a[43] & b[84])^(a[42] & b[85])^(a[41] & b[86])^(a[40] & b[87])^(a[39] & b[88])^(a[38] & b[89])^(a[37] & b[90])^(a[36] & b[91])^(a[35] & b[92])^(a[34] & b[93])^(a[33] & b[94])^(a[32] & b[95])^(a[31] & b[96])^(a[30] & b[97])^(a[29] & b[98])^(a[28] & b[99])^(a[27] & b[100])^(a[26] & b[101])^(a[25] & b[102])^(a[24] & b[103])^(a[23] & b[104])^(a[22] & b[105])^(a[21] & b[106])^(a[20] & b[107])^(a[19] & b[108])^(a[18] & b[109])^(a[17] & b[110])^(a[16] & b[111])^(a[15] & b[112])^(a[14] & b[113])^(a[13] & b[114])^(a[12] & b[115])^(a[11] & b[116])^(a[10] & b[117])^(a[9] & b[118])^(a[8] & b[119])^(a[7] & b[120])^(a[6] & b[121])^(a[5] & b[122])^(a[4] & b[123])^(a[3] & b[124])^(a[2] & b[125])^(a[1] & b[126])^(a[0] & b[127]);
assign y[128] = (a[128] & b[0])^(a[127] & b[1])^(a[126] & b[2])^(a[125] & b[3])^(a[124] & b[4])^(a[123] & b[5])^(a[122] & b[6])^(a[121] & b[7])^(a[120] & b[8])^(a[119] & b[9])^(a[118] & b[10])^(a[117] & b[11])^(a[116] & b[12])^(a[115] & b[13])^(a[114] & b[14])^(a[113] & b[15])^(a[112] & b[16])^(a[111] & b[17])^(a[110] & b[18])^(a[109] & b[19])^(a[108] & b[20])^(a[107] & b[21])^(a[106] & b[22])^(a[105] & b[23])^(a[104] & b[24])^(a[103] & b[25])^(a[102] & b[26])^(a[101] & b[27])^(a[100] & b[28])^(a[99] & b[29])^(a[98] & b[30])^(a[97] & b[31])^(a[96] & b[32])^(a[95] & b[33])^(a[94] & b[34])^(a[93] & b[35])^(a[92] & b[36])^(a[91] & b[37])^(a[90] & b[38])^(a[89] & b[39])^(a[88] & b[40])^(a[87] & b[41])^(a[86] & b[42])^(a[85] & b[43])^(a[84] & b[44])^(a[83] & b[45])^(a[82] & b[46])^(a[81] & b[47])^(a[80] & b[48])^(a[79] & b[49])^(a[78] & b[50])^(a[77] & b[51])^(a[76] & b[52])^(a[75] & b[53])^(a[74] & b[54])^(a[73] & b[55])^(a[72] & b[56])^(a[71] & b[57])^(a[70] & b[58])^(a[69] & b[59])^(a[68] & b[60])^(a[67] & b[61])^(a[66] & b[62])^(a[65] & b[63])^(a[64] & b[64])^(a[63] & b[65])^(a[62] & b[66])^(a[61] & b[67])^(a[60] & b[68])^(a[59] & b[69])^(a[58] & b[70])^(a[57] & b[71])^(a[56] & b[72])^(a[55] & b[73])^(a[54] & b[74])^(a[53] & b[75])^(a[52] & b[76])^(a[51] & b[77])^(a[50] & b[78])^(a[49] & b[79])^(a[48] & b[80])^(a[47] & b[81])^(a[46] & b[82])^(a[45] & b[83])^(a[44] & b[84])^(a[43] & b[85])^(a[42] & b[86])^(a[41] & b[87])^(a[40] & b[88])^(a[39] & b[89])^(a[38] & b[90])^(a[37] & b[91])^(a[36] & b[92])^(a[35] & b[93])^(a[34] & b[94])^(a[33] & b[95])^(a[32] & b[96])^(a[31] & b[97])^(a[30] & b[98])^(a[29] & b[99])^(a[28] & b[100])^(a[27] & b[101])^(a[26] & b[102])^(a[25] & b[103])^(a[24] & b[104])^(a[23] & b[105])^(a[22] & b[106])^(a[21] & b[107])^(a[20] & b[108])^(a[19] & b[109])^(a[18] & b[110])^(a[17] & b[111])^(a[16] & b[112])^(a[15] & b[113])^(a[14] & b[114])^(a[13] & b[115])^(a[12] & b[116])^(a[11] & b[117])^(a[10] & b[118])^(a[9] & b[119])^(a[8] & b[120])^(a[7] & b[121])^(a[6] & b[122])^(a[5] & b[123])^(a[4] & b[124])^(a[3] & b[125])^(a[2] & b[126])^(a[1] & b[127])^(a[0] & b[128]);
assign y[129] = (a[129] & b[0])^(a[128] & b[1])^(a[127] & b[2])^(a[126] & b[3])^(a[125] & b[4])^(a[124] & b[5])^(a[123] & b[6])^(a[122] & b[7])^(a[121] & b[8])^(a[120] & b[9])^(a[119] & b[10])^(a[118] & b[11])^(a[117] & b[12])^(a[116] & b[13])^(a[115] & b[14])^(a[114] & b[15])^(a[113] & b[16])^(a[112] & b[17])^(a[111] & b[18])^(a[110] & b[19])^(a[109] & b[20])^(a[108] & b[21])^(a[107] & b[22])^(a[106] & b[23])^(a[105] & b[24])^(a[104] & b[25])^(a[103] & b[26])^(a[102] & b[27])^(a[101] & b[28])^(a[100] & b[29])^(a[99] & b[30])^(a[98] & b[31])^(a[97] & b[32])^(a[96] & b[33])^(a[95] & b[34])^(a[94] & b[35])^(a[93] & b[36])^(a[92] & b[37])^(a[91] & b[38])^(a[90] & b[39])^(a[89] & b[40])^(a[88] & b[41])^(a[87] & b[42])^(a[86] & b[43])^(a[85] & b[44])^(a[84] & b[45])^(a[83] & b[46])^(a[82] & b[47])^(a[81] & b[48])^(a[80] & b[49])^(a[79] & b[50])^(a[78] & b[51])^(a[77] & b[52])^(a[76] & b[53])^(a[75] & b[54])^(a[74] & b[55])^(a[73] & b[56])^(a[72] & b[57])^(a[71] & b[58])^(a[70] & b[59])^(a[69] & b[60])^(a[68] & b[61])^(a[67] & b[62])^(a[66] & b[63])^(a[65] & b[64])^(a[64] & b[65])^(a[63] & b[66])^(a[62] & b[67])^(a[61] & b[68])^(a[60] & b[69])^(a[59] & b[70])^(a[58] & b[71])^(a[57] & b[72])^(a[56] & b[73])^(a[55] & b[74])^(a[54] & b[75])^(a[53] & b[76])^(a[52] & b[77])^(a[51] & b[78])^(a[50] & b[79])^(a[49] & b[80])^(a[48] & b[81])^(a[47] & b[82])^(a[46] & b[83])^(a[45] & b[84])^(a[44] & b[85])^(a[43] & b[86])^(a[42] & b[87])^(a[41] & b[88])^(a[40] & b[89])^(a[39] & b[90])^(a[38] & b[91])^(a[37] & b[92])^(a[36] & b[93])^(a[35] & b[94])^(a[34] & b[95])^(a[33] & b[96])^(a[32] & b[97])^(a[31] & b[98])^(a[30] & b[99])^(a[29] & b[100])^(a[28] & b[101])^(a[27] & b[102])^(a[26] & b[103])^(a[25] & b[104])^(a[24] & b[105])^(a[23] & b[106])^(a[22] & b[107])^(a[21] & b[108])^(a[20] & b[109])^(a[19] & b[110])^(a[18] & b[111])^(a[17] & b[112])^(a[16] & b[113])^(a[15] & b[114])^(a[14] & b[115])^(a[13] & b[116])^(a[12] & b[117])^(a[11] & b[118])^(a[10] & b[119])^(a[9] & b[120])^(a[8] & b[121])^(a[7] & b[122])^(a[6] & b[123])^(a[5] & b[124])^(a[4] & b[125])^(a[3] & b[126])^(a[2] & b[127])^(a[1] & b[128])^(a[0] & b[129]);
assign y[130] = (a[130] & b[0])^(a[129] & b[1])^(a[128] & b[2])^(a[127] & b[3])^(a[126] & b[4])^(a[125] & b[5])^(a[124] & b[6])^(a[123] & b[7])^(a[122] & b[8])^(a[121] & b[9])^(a[120] & b[10])^(a[119] & b[11])^(a[118] & b[12])^(a[117] & b[13])^(a[116] & b[14])^(a[115] & b[15])^(a[114] & b[16])^(a[113] & b[17])^(a[112] & b[18])^(a[111] & b[19])^(a[110] & b[20])^(a[109] & b[21])^(a[108] & b[22])^(a[107] & b[23])^(a[106] & b[24])^(a[105] & b[25])^(a[104] & b[26])^(a[103] & b[27])^(a[102] & b[28])^(a[101] & b[29])^(a[100] & b[30])^(a[99] & b[31])^(a[98] & b[32])^(a[97] & b[33])^(a[96] & b[34])^(a[95] & b[35])^(a[94] & b[36])^(a[93] & b[37])^(a[92] & b[38])^(a[91] & b[39])^(a[90] & b[40])^(a[89] & b[41])^(a[88] & b[42])^(a[87] & b[43])^(a[86] & b[44])^(a[85] & b[45])^(a[84] & b[46])^(a[83] & b[47])^(a[82] & b[48])^(a[81] & b[49])^(a[80] & b[50])^(a[79] & b[51])^(a[78] & b[52])^(a[77] & b[53])^(a[76] & b[54])^(a[75] & b[55])^(a[74] & b[56])^(a[73] & b[57])^(a[72] & b[58])^(a[71] & b[59])^(a[70] & b[60])^(a[69] & b[61])^(a[68] & b[62])^(a[67] & b[63])^(a[66] & b[64])^(a[65] & b[65])^(a[64] & b[66])^(a[63] & b[67])^(a[62] & b[68])^(a[61] & b[69])^(a[60] & b[70])^(a[59] & b[71])^(a[58] & b[72])^(a[57] & b[73])^(a[56] & b[74])^(a[55] & b[75])^(a[54] & b[76])^(a[53] & b[77])^(a[52] & b[78])^(a[51] & b[79])^(a[50] & b[80])^(a[49] & b[81])^(a[48] & b[82])^(a[47] & b[83])^(a[46] & b[84])^(a[45] & b[85])^(a[44] & b[86])^(a[43] & b[87])^(a[42] & b[88])^(a[41] & b[89])^(a[40] & b[90])^(a[39] & b[91])^(a[38] & b[92])^(a[37] & b[93])^(a[36] & b[94])^(a[35] & b[95])^(a[34] & b[96])^(a[33] & b[97])^(a[32] & b[98])^(a[31] & b[99])^(a[30] & b[100])^(a[29] & b[101])^(a[28] & b[102])^(a[27] & b[103])^(a[26] & b[104])^(a[25] & b[105])^(a[24] & b[106])^(a[23] & b[107])^(a[22] & b[108])^(a[21] & b[109])^(a[20] & b[110])^(a[19] & b[111])^(a[18] & b[112])^(a[17] & b[113])^(a[16] & b[114])^(a[15] & b[115])^(a[14] & b[116])^(a[13] & b[117])^(a[12] & b[118])^(a[11] & b[119])^(a[10] & b[120])^(a[9] & b[121])^(a[8] & b[122])^(a[7] & b[123])^(a[6] & b[124])^(a[5] & b[125])^(a[4] & b[126])^(a[3] & b[127])^(a[2] & b[128])^(a[1] & b[129])^(a[0] & b[130]);
assign y[131] = (a[131] & b[0])^(a[130] & b[1])^(a[129] & b[2])^(a[128] & b[3])^(a[127] & b[4])^(a[126] & b[5])^(a[125] & b[6])^(a[124] & b[7])^(a[123] & b[8])^(a[122] & b[9])^(a[121] & b[10])^(a[120] & b[11])^(a[119] & b[12])^(a[118] & b[13])^(a[117] & b[14])^(a[116] & b[15])^(a[115] & b[16])^(a[114] & b[17])^(a[113] & b[18])^(a[112] & b[19])^(a[111] & b[20])^(a[110] & b[21])^(a[109] & b[22])^(a[108] & b[23])^(a[107] & b[24])^(a[106] & b[25])^(a[105] & b[26])^(a[104] & b[27])^(a[103] & b[28])^(a[102] & b[29])^(a[101] & b[30])^(a[100] & b[31])^(a[99] & b[32])^(a[98] & b[33])^(a[97] & b[34])^(a[96] & b[35])^(a[95] & b[36])^(a[94] & b[37])^(a[93] & b[38])^(a[92] & b[39])^(a[91] & b[40])^(a[90] & b[41])^(a[89] & b[42])^(a[88] & b[43])^(a[87] & b[44])^(a[86] & b[45])^(a[85] & b[46])^(a[84] & b[47])^(a[83] & b[48])^(a[82] & b[49])^(a[81] & b[50])^(a[80] & b[51])^(a[79] & b[52])^(a[78] & b[53])^(a[77] & b[54])^(a[76] & b[55])^(a[75] & b[56])^(a[74] & b[57])^(a[73] & b[58])^(a[72] & b[59])^(a[71] & b[60])^(a[70] & b[61])^(a[69] & b[62])^(a[68] & b[63])^(a[67] & b[64])^(a[66] & b[65])^(a[65] & b[66])^(a[64] & b[67])^(a[63] & b[68])^(a[62] & b[69])^(a[61] & b[70])^(a[60] & b[71])^(a[59] & b[72])^(a[58] & b[73])^(a[57] & b[74])^(a[56] & b[75])^(a[55] & b[76])^(a[54] & b[77])^(a[53] & b[78])^(a[52] & b[79])^(a[51] & b[80])^(a[50] & b[81])^(a[49] & b[82])^(a[48] & b[83])^(a[47] & b[84])^(a[46] & b[85])^(a[45] & b[86])^(a[44] & b[87])^(a[43] & b[88])^(a[42] & b[89])^(a[41] & b[90])^(a[40] & b[91])^(a[39] & b[92])^(a[38] & b[93])^(a[37] & b[94])^(a[36] & b[95])^(a[35] & b[96])^(a[34] & b[97])^(a[33] & b[98])^(a[32] & b[99])^(a[31] & b[100])^(a[30] & b[101])^(a[29] & b[102])^(a[28] & b[103])^(a[27] & b[104])^(a[26] & b[105])^(a[25] & b[106])^(a[24] & b[107])^(a[23] & b[108])^(a[22] & b[109])^(a[21] & b[110])^(a[20] & b[111])^(a[19] & b[112])^(a[18] & b[113])^(a[17] & b[114])^(a[16] & b[115])^(a[15] & b[116])^(a[14] & b[117])^(a[13] & b[118])^(a[12] & b[119])^(a[11] & b[120])^(a[10] & b[121])^(a[9] & b[122])^(a[8] & b[123])^(a[7] & b[124])^(a[6] & b[125])^(a[5] & b[126])^(a[4] & b[127])^(a[3] & b[128])^(a[2] & b[129])^(a[1] & b[130])^(a[0] & b[131]);
assign y[132] = (a[132] & b[0])^(a[131] & b[1])^(a[130] & b[2])^(a[129] & b[3])^(a[128] & b[4])^(a[127] & b[5])^(a[126] & b[6])^(a[125] & b[7])^(a[124] & b[8])^(a[123] & b[9])^(a[122] & b[10])^(a[121] & b[11])^(a[120] & b[12])^(a[119] & b[13])^(a[118] & b[14])^(a[117] & b[15])^(a[116] & b[16])^(a[115] & b[17])^(a[114] & b[18])^(a[113] & b[19])^(a[112] & b[20])^(a[111] & b[21])^(a[110] & b[22])^(a[109] & b[23])^(a[108] & b[24])^(a[107] & b[25])^(a[106] & b[26])^(a[105] & b[27])^(a[104] & b[28])^(a[103] & b[29])^(a[102] & b[30])^(a[101] & b[31])^(a[100] & b[32])^(a[99] & b[33])^(a[98] & b[34])^(a[97] & b[35])^(a[96] & b[36])^(a[95] & b[37])^(a[94] & b[38])^(a[93] & b[39])^(a[92] & b[40])^(a[91] & b[41])^(a[90] & b[42])^(a[89] & b[43])^(a[88] & b[44])^(a[87] & b[45])^(a[86] & b[46])^(a[85] & b[47])^(a[84] & b[48])^(a[83] & b[49])^(a[82] & b[50])^(a[81] & b[51])^(a[80] & b[52])^(a[79] & b[53])^(a[78] & b[54])^(a[77] & b[55])^(a[76] & b[56])^(a[75] & b[57])^(a[74] & b[58])^(a[73] & b[59])^(a[72] & b[60])^(a[71] & b[61])^(a[70] & b[62])^(a[69] & b[63])^(a[68] & b[64])^(a[67] & b[65])^(a[66] & b[66])^(a[65] & b[67])^(a[64] & b[68])^(a[63] & b[69])^(a[62] & b[70])^(a[61] & b[71])^(a[60] & b[72])^(a[59] & b[73])^(a[58] & b[74])^(a[57] & b[75])^(a[56] & b[76])^(a[55] & b[77])^(a[54] & b[78])^(a[53] & b[79])^(a[52] & b[80])^(a[51] & b[81])^(a[50] & b[82])^(a[49] & b[83])^(a[48] & b[84])^(a[47] & b[85])^(a[46] & b[86])^(a[45] & b[87])^(a[44] & b[88])^(a[43] & b[89])^(a[42] & b[90])^(a[41] & b[91])^(a[40] & b[92])^(a[39] & b[93])^(a[38] & b[94])^(a[37] & b[95])^(a[36] & b[96])^(a[35] & b[97])^(a[34] & b[98])^(a[33] & b[99])^(a[32] & b[100])^(a[31] & b[101])^(a[30] & b[102])^(a[29] & b[103])^(a[28] & b[104])^(a[27] & b[105])^(a[26] & b[106])^(a[25] & b[107])^(a[24] & b[108])^(a[23] & b[109])^(a[22] & b[110])^(a[21] & b[111])^(a[20] & b[112])^(a[19] & b[113])^(a[18] & b[114])^(a[17] & b[115])^(a[16] & b[116])^(a[15] & b[117])^(a[14] & b[118])^(a[13] & b[119])^(a[12] & b[120])^(a[11] & b[121])^(a[10] & b[122])^(a[9] & b[123])^(a[8] & b[124])^(a[7] & b[125])^(a[6] & b[126])^(a[5] & b[127])^(a[4] & b[128])^(a[3] & b[129])^(a[2] & b[130])^(a[1] & b[131])^(a[0] & b[132]);
assign y[133] = (a[133] & b[0])^(a[132] & b[1])^(a[131] & b[2])^(a[130] & b[3])^(a[129] & b[4])^(a[128] & b[5])^(a[127] & b[6])^(a[126] & b[7])^(a[125] & b[8])^(a[124] & b[9])^(a[123] & b[10])^(a[122] & b[11])^(a[121] & b[12])^(a[120] & b[13])^(a[119] & b[14])^(a[118] & b[15])^(a[117] & b[16])^(a[116] & b[17])^(a[115] & b[18])^(a[114] & b[19])^(a[113] & b[20])^(a[112] & b[21])^(a[111] & b[22])^(a[110] & b[23])^(a[109] & b[24])^(a[108] & b[25])^(a[107] & b[26])^(a[106] & b[27])^(a[105] & b[28])^(a[104] & b[29])^(a[103] & b[30])^(a[102] & b[31])^(a[101] & b[32])^(a[100] & b[33])^(a[99] & b[34])^(a[98] & b[35])^(a[97] & b[36])^(a[96] & b[37])^(a[95] & b[38])^(a[94] & b[39])^(a[93] & b[40])^(a[92] & b[41])^(a[91] & b[42])^(a[90] & b[43])^(a[89] & b[44])^(a[88] & b[45])^(a[87] & b[46])^(a[86] & b[47])^(a[85] & b[48])^(a[84] & b[49])^(a[83] & b[50])^(a[82] & b[51])^(a[81] & b[52])^(a[80] & b[53])^(a[79] & b[54])^(a[78] & b[55])^(a[77] & b[56])^(a[76] & b[57])^(a[75] & b[58])^(a[74] & b[59])^(a[73] & b[60])^(a[72] & b[61])^(a[71] & b[62])^(a[70] & b[63])^(a[69] & b[64])^(a[68] & b[65])^(a[67] & b[66])^(a[66] & b[67])^(a[65] & b[68])^(a[64] & b[69])^(a[63] & b[70])^(a[62] & b[71])^(a[61] & b[72])^(a[60] & b[73])^(a[59] & b[74])^(a[58] & b[75])^(a[57] & b[76])^(a[56] & b[77])^(a[55] & b[78])^(a[54] & b[79])^(a[53] & b[80])^(a[52] & b[81])^(a[51] & b[82])^(a[50] & b[83])^(a[49] & b[84])^(a[48] & b[85])^(a[47] & b[86])^(a[46] & b[87])^(a[45] & b[88])^(a[44] & b[89])^(a[43] & b[90])^(a[42] & b[91])^(a[41] & b[92])^(a[40] & b[93])^(a[39] & b[94])^(a[38] & b[95])^(a[37] & b[96])^(a[36] & b[97])^(a[35] & b[98])^(a[34] & b[99])^(a[33] & b[100])^(a[32] & b[101])^(a[31] & b[102])^(a[30] & b[103])^(a[29] & b[104])^(a[28] & b[105])^(a[27] & b[106])^(a[26] & b[107])^(a[25] & b[108])^(a[24] & b[109])^(a[23] & b[110])^(a[22] & b[111])^(a[21] & b[112])^(a[20] & b[113])^(a[19] & b[114])^(a[18] & b[115])^(a[17] & b[116])^(a[16] & b[117])^(a[15] & b[118])^(a[14] & b[119])^(a[13] & b[120])^(a[12] & b[121])^(a[11] & b[122])^(a[10] & b[123])^(a[9] & b[124])^(a[8] & b[125])^(a[7] & b[126])^(a[6] & b[127])^(a[5] & b[128])^(a[4] & b[129])^(a[3] & b[130])^(a[2] & b[131])^(a[1] & b[132])^(a[0] & b[133]);
assign y[134] = (a[134] & b[0])^(a[133] & b[1])^(a[132] & b[2])^(a[131] & b[3])^(a[130] & b[4])^(a[129] & b[5])^(a[128] & b[6])^(a[127] & b[7])^(a[126] & b[8])^(a[125] & b[9])^(a[124] & b[10])^(a[123] & b[11])^(a[122] & b[12])^(a[121] & b[13])^(a[120] & b[14])^(a[119] & b[15])^(a[118] & b[16])^(a[117] & b[17])^(a[116] & b[18])^(a[115] & b[19])^(a[114] & b[20])^(a[113] & b[21])^(a[112] & b[22])^(a[111] & b[23])^(a[110] & b[24])^(a[109] & b[25])^(a[108] & b[26])^(a[107] & b[27])^(a[106] & b[28])^(a[105] & b[29])^(a[104] & b[30])^(a[103] & b[31])^(a[102] & b[32])^(a[101] & b[33])^(a[100] & b[34])^(a[99] & b[35])^(a[98] & b[36])^(a[97] & b[37])^(a[96] & b[38])^(a[95] & b[39])^(a[94] & b[40])^(a[93] & b[41])^(a[92] & b[42])^(a[91] & b[43])^(a[90] & b[44])^(a[89] & b[45])^(a[88] & b[46])^(a[87] & b[47])^(a[86] & b[48])^(a[85] & b[49])^(a[84] & b[50])^(a[83] & b[51])^(a[82] & b[52])^(a[81] & b[53])^(a[80] & b[54])^(a[79] & b[55])^(a[78] & b[56])^(a[77] & b[57])^(a[76] & b[58])^(a[75] & b[59])^(a[74] & b[60])^(a[73] & b[61])^(a[72] & b[62])^(a[71] & b[63])^(a[70] & b[64])^(a[69] & b[65])^(a[68] & b[66])^(a[67] & b[67])^(a[66] & b[68])^(a[65] & b[69])^(a[64] & b[70])^(a[63] & b[71])^(a[62] & b[72])^(a[61] & b[73])^(a[60] & b[74])^(a[59] & b[75])^(a[58] & b[76])^(a[57] & b[77])^(a[56] & b[78])^(a[55] & b[79])^(a[54] & b[80])^(a[53] & b[81])^(a[52] & b[82])^(a[51] & b[83])^(a[50] & b[84])^(a[49] & b[85])^(a[48] & b[86])^(a[47] & b[87])^(a[46] & b[88])^(a[45] & b[89])^(a[44] & b[90])^(a[43] & b[91])^(a[42] & b[92])^(a[41] & b[93])^(a[40] & b[94])^(a[39] & b[95])^(a[38] & b[96])^(a[37] & b[97])^(a[36] & b[98])^(a[35] & b[99])^(a[34] & b[100])^(a[33] & b[101])^(a[32] & b[102])^(a[31] & b[103])^(a[30] & b[104])^(a[29] & b[105])^(a[28] & b[106])^(a[27] & b[107])^(a[26] & b[108])^(a[25] & b[109])^(a[24] & b[110])^(a[23] & b[111])^(a[22] & b[112])^(a[21] & b[113])^(a[20] & b[114])^(a[19] & b[115])^(a[18] & b[116])^(a[17] & b[117])^(a[16] & b[118])^(a[15] & b[119])^(a[14] & b[120])^(a[13] & b[121])^(a[12] & b[122])^(a[11] & b[123])^(a[10] & b[124])^(a[9] & b[125])^(a[8] & b[126])^(a[7] & b[127])^(a[6] & b[128])^(a[5] & b[129])^(a[4] & b[130])^(a[3] & b[131])^(a[2] & b[132])^(a[1] & b[133])^(a[0] & b[134]);
assign y[135] = (a[135] & b[0])^(a[134] & b[1])^(a[133] & b[2])^(a[132] & b[3])^(a[131] & b[4])^(a[130] & b[5])^(a[129] & b[6])^(a[128] & b[7])^(a[127] & b[8])^(a[126] & b[9])^(a[125] & b[10])^(a[124] & b[11])^(a[123] & b[12])^(a[122] & b[13])^(a[121] & b[14])^(a[120] & b[15])^(a[119] & b[16])^(a[118] & b[17])^(a[117] & b[18])^(a[116] & b[19])^(a[115] & b[20])^(a[114] & b[21])^(a[113] & b[22])^(a[112] & b[23])^(a[111] & b[24])^(a[110] & b[25])^(a[109] & b[26])^(a[108] & b[27])^(a[107] & b[28])^(a[106] & b[29])^(a[105] & b[30])^(a[104] & b[31])^(a[103] & b[32])^(a[102] & b[33])^(a[101] & b[34])^(a[100] & b[35])^(a[99] & b[36])^(a[98] & b[37])^(a[97] & b[38])^(a[96] & b[39])^(a[95] & b[40])^(a[94] & b[41])^(a[93] & b[42])^(a[92] & b[43])^(a[91] & b[44])^(a[90] & b[45])^(a[89] & b[46])^(a[88] & b[47])^(a[87] & b[48])^(a[86] & b[49])^(a[85] & b[50])^(a[84] & b[51])^(a[83] & b[52])^(a[82] & b[53])^(a[81] & b[54])^(a[80] & b[55])^(a[79] & b[56])^(a[78] & b[57])^(a[77] & b[58])^(a[76] & b[59])^(a[75] & b[60])^(a[74] & b[61])^(a[73] & b[62])^(a[72] & b[63])^(a[71] & b[64])^(a[70] & b[65])^(a[69] & b[66])^(a[68] & b[67])^(a[67] & b[68])^(a[66] & b[69])^(a[65] & b[70])^(a[64] & b[71])^(a[63] & b[72])^(a[62] & b[73])^(a[61] & b[74])^(a[60] & b[75])^(a[59] & b[76])^(a[58] & b[77])^(a[57] & b[78])^(a[56] & b[79])^(a[55] & b[80])^(a[54] & b[81])^(a[53] & b[82])^(a[52] & b[83])^(a[51] & b[84])^(a[50] & b[85])^(a[49] & b[86])^(a[48] & b[87])^(a[47] & b[88])^(a[46] & b[89])^(a[45] & b[90])^(a[44] & b[91])^(a[43] & b[92])^(a[42] & b[93])^(a[41] & b[94])^(a[40] & b[95])^(a[39] & b[96])^(a[38] & b[97])^(a[37] & b[98])^(a[36] & b[99])^(a[35] & b[100])^(a[34] & b[101])^(a[33] & b[102])^(a[32] & b[103])^(a[31] & b[104])^(a[30] & b[105])^(a[29] & b[106])^(a[28] & b[107])^(a[27] & b[108])^(a[26] & b[109])^(a[25] & b[110])^(a[24] & b[111])^(a[23] & b[112])^(a[22] & b[113])^(a[21] & b[114])^(a[20] & b[115])^(a[19] & b[116])^(a[18] & b[117])^(a[17] & b[118])^(a[16] & b[119])^(a[15] & b[120])^(a[14] & b[121])^(a[13] & b[122])^(a[12] & b[123])^(a[11] & b[124])^(a[10] & b[125])^(a[9] & b[126])^(a[8] & b[127])^(a[7] & b[128])^(a[6] & b[129])^(a[5] & b[130])^(a[4] & b[131])^(a[3] & b[132])^(a[2] & b[133])^(a[1] & b[134])^(a[0] & b[135]);
assign y[136] = (a[136] & b[0])^(a[135] & b[1])^(a[134] & b[2])^(a[133] & b[3])^(a[132] & b[4])^(a[131] & b[5])^(a[130] & b[6])^(a[129] & b[7])^(a[128] & b[8])^(a[127] & b[9])^(a[126] & b[10])^(a[125] & b[11])^(a[124] & b[12])^(a[123] & b[13])^(a[122] & b[14])^(a[121] & b[15])^(a[120] & b[16])^(a[119] & b[17])^(a[118] & b[18])^(a[117] & b[19])^(a[116] & b[20])^(a[115] & b[21])^(a[114] & b[22])^(a[113] & b[23])^(a[112] & b[24])^(a[111] & b[25])^(a[110] & b[26])^(a[109] & b[27])^(a[108] & b[28])^(a[107] & b[29])^(a[106] & b[30])^(a[105] & b[31])^(a[104] & b[32])^(a[103] & b[33])^(a[102] & b[34])^(a[101] & b[35])^(a[100] & b[36])^(a[99] & b[37])^(a[98] & b[38])^(a[97] & b[39])^(a[96] & b[40])^(a[95] & b[41])^(a[94] & b[42])^(a[93] & b[43])^(a[92] & b[44])^(a[91] & b[45])^(a[90] & b[46])^(a[89] & b[47])^(a[88] & b[48])^(a[87] & b[49])^(a[86] & b[50])^(a[85] & b[51])^(a[84] & b[52])^(a[83] & b[53])^(a[82] & b[54])^(a[81] & b[55])^(a[80] & b[56])^(a[79] & b[57])^(a[78] & b[58])^(a[77] & b[59])^(a[76] & b[60])^(a[75] & b[61])^(a[74] & b[62])^(a[73] & b[63])^(a[72] & b[64])^(a[71] & b[65])^(a[70] & b[66])^(a[69] & b[67])^(a[68] & b[68])^(a[67] & b[69])^(a[66] & b[70])^(a[65] & b[71])^(a[64] & b[72])^(a[63] & b[73])^(a[62] & b[74])^(a[61] & b[75])^(a[60] & b[76])^(a[59] & b[77])^(a[58] & b[78])^(a[57] & b[79])^(a[56] & b[80])^(a[55] & b[81])^(a[54] & b[82])^(a[53] & b[83])^(a[52] & b[84])^(a[51] & b[85])^(a[50] & b[86])^(a[49] & b[87])^(a[48] & b[88])^(a[47] & b[89])^(a[46] & b[90])^(a[45] & b[91])^(a[44] & b[92])^(a[43] & b[93])^(a[42] & b[94])^(a[41] & b[95])^(a[40] & b[96])^(a[39] & b[97])^(a[38] & b[98])^(a[37] & b[99])^(a[36] & b[100])^(a[35] & b[101])^(a[34] & b[102])^(a[33] & b[103])^(a[32] & b[104])^(a[31] & b[105])^(a[30] & b[106])^(a[29] & b[107])^(a[28] & b[108])^(a[27] & b[109])^(a[26] & b[110])^(a[25] & b[111])^(a[24] & b[112])^(a[23] & b[113])^(a[22] & b[114])^(a[21] & b[115])^(a[20] & b[116])^(a[19] & b[117])^(a[18] & b[118])^(a[17] & b[119])^(a[16] & b[120])^(a[15] & b[121])^(a[14] & b[122])^(a[13] & b[123])^(a[12] & b[124])^(a[11] & b[125])^(a[10] & b[126])^(a[9] & b[127])^(a[8] & b[128])^(a[7] & b[129])^(a[6] & b[130])^(a[5] & b[131])^(a[4] & b[132])^(a[3] & b[133])^(a[2] & b[134])^(a[1] & b[135])^(a[0] & b[136]);
assign y[137] = (a[137] & b[0])^(a[136] & b[1])^(a[135] & b[2])^(a[134] & b[3])^(a[133] & b[4])^(a[132] & b[5])^(a[131] & b[6])^(a[130] & b[7])^(a[129] & b[8])^(a[128] & b[9])^(a[127] & b[10])^(a[126] & b[11])^(a[125] & b[12])^(a[124] & b[13])^(a[123] & b[14])^(a[122] & b[15])^(a[121] & b[16])^(a[120] & b[17])^(a[119] & b[18])^(a[118] & b[19])^(a[117] & b[20])^(a[116] & b[21])^(a[115] & b[22])^(a[114] & b[23])^(a[113] & b[24])^(a[112] & b[25])^(a[111] & b[26])^(a[110] & b[27])^(a[109] & b[28])^(a[108] & b[29])^(a[107] & b[30])^(a[106] & b[31])^(a[105] & b[32])^(a[104] & b[33])^(a[103] & b[34])^(a[102] & b[35])^(a[101] & b[36])^(a[100] & b[37])^(a[99] & b[38])^(a[98] & b[39])^(a[97] & b[40])^(a[96] & b[41])^(a[95] & b[42])^(a[94] & b[43])^(a[93] & b[44])^(a[92] & b[45])^(a[91] & b[46])^(a[90] & b[47])^(a[89] & b[48])^(a[88] & b[49])^(a[87] & b[50])^(a[86] & b[51])^(a[85] & b[52])^(a[84] & b[53])^(a[83] & b[54])^(a[82] & b[55])^(a[81] & b[56])^(a[80] & b[57])^(a[79] & b[58])^(a[78] & b[59])^(a[77] & b[60])^(a[76] & b[61])^(a[75] & b[62])^(a[74] & b[63])^(a[73] & b[64])^(a[72] & b[65])^(a[71] & b[66])^(a[70] & b[67])^(a[69] & b[68])^(a[68] & b[69])^(a[67] & b[70])^(a[66] & b[71])^(a[65] & b[72])^(a[64] & b[73])^(a[63] & b[74])^(a[62] & b[75])^(a[61] & b[76])^(a[60] & b[77])^(a[59] & b[78])^(a[58] & b[79])^(a[57] & b[80])^(a[56] & b[81])^(a[55] & b[82])^(a[54] & b[83])^(a[53] & b[84])^(a[52] & b[85])^(a[51] & b[86])^(a[50] & b[87])^(a[49] & b[88])^(a[48] & b[89])^(a[47] & b[90])^(a[46] & b[91])^(a[45] & b[92])^(a[44] & b[93])^(a[43] & b[94])^(a[42] & b[95])^(a[41] & b[96])^(a[40] & b[97])^(a[39] & b[98])^(a[38] & b[99])^(a[37] & b[100])^(a[36] & b[101])^(a[35] & b[102])^(a[34] & b[103])^(a[33] & b[104])^(a[32] & b[105])^(a[31] & b[106])^(a[30] & b[107])^(a[29] & b[108])^(a[28] & b[109])^(a[27] & b[110])^(a[26] & b[111])^(a[25] & b[112])^(a[24] & b[113])^(a[23] & b[114])^(a[22] & b[115])^(a[21] & b[116])^(a[20] & b[117])^(a[19] & b[118])^(a[18] & b[119])^(a[17] & b[120])^(a[16] & b[121])^(a[15] & b[122])^(a[14] & b[123])^(a[13] & b[124])^(a[12] & b[125])^(a[11] & b[126])^(a[10] & b[127])^(a[9] & b[128])^(a[8] & b[129])^(a[7] & b[130])^(a[6] & b[131])^(a[5] & b[132])^(a[4] & b[133])^(a[3] & b[134])^(a[2] & b[135])^(a[1] & b[136])^(a[0] & b[137]);
assign y[138] = (a[138] & b[0])^(a[137] & b[1])^(a[136] & b[2])^(a[135] & b[3])^(a[134] & b[4])^(a[133] & b[5])^(a[132] & b[6])^(a[131] & b[7])^(a[130] & b[8])^(a[129] & b[9])^(a[128] & b[10])^(a[127] & b[11])^(a[126] & b[12])^(a[125] & b[13])^(a[124] & b[14])^(a[123] & b[15])^(a[122] & b[16])^(a[121] & b[17])^(a[120] & b[18])^(a[119] & b[19])^(a[118] & b[20])^(a[117] & b[21])^(a[116] & b[22])^(a[115] & b[23])^(a[114] & b[24])^(a[113] & b[25])^(a[112] & b[26])^(a[111] & b[27])^(a[110] & b[28])^(a[109] & b[29])^(a[108] & b[30])^(a[107] & b[31])^(a[106] & b[32])^(a[105] & b[33])^(a[104] & b[34])^(a[103] & b[35])^(a[102] & b[36])^(a[101] & b[37])^(a[100] & b[38])^(a[99] & b[39])^(a[98] & b[40])^(a[97] & b[41])^(a[96] & b[42])^(a[95] & b[43])^(a[94] & b[44])^(a[93] & b[45])^(a[92] & b[46])^(a[91] & b[47])^(a[90] & b[48])^(a[89] & b[49])^(a[88] & b[50])^(a[87] & b[51])^(a[86] & b[52])^(a[85] & b[53])^(a[84] & b[54])^(a[83] & b[55])^(a[82] & b[56])^(a[81] & b[57])^(a[80] & b[58])^(a[79] & b[59])^(a[78] & b[60])^(a[77] & b[61])^(a[76] & b[62])^(a[75] & b[63])^(a[74] & b[64])^(a[73] & b[65])^(a[72] & b[66])^(a[71] & b[67])^(a[70] & b[68])^(a[69] & b[69])^(a[68] & b[70])^(a[67] & b[71])^(a[66] & b[72])^(a[65] & b[73])^(a[64] & b[74])^(a[63] & b[75])^(a[62] & b[76])^(a[61] & b[77])^(a[60] & b[78])^(a[59] & b[79])^(a[58] & b[80])^(a[57] & b[81])^(a[56] & b[82])^(a[55] & b[83])^(a[54] & b[84])^(a[53] & b[85])^(a[52] & b[86])^(a[51] & b[87])^(a[50] & b[88])^(a[49] & b[89])^(a[48] & b[90])^(a[47] & b[91])^(a[46] & b[92])^(a[45] & b[93])^(a[44] & b[94])^(a[43] & b[95])^(a[42] & b[96])^(a[41] & b[97])^(a[40] & b[98])^(a[39] & b[99])^(a[38] & b[100])^(a[37] & b[101])^(a[36] & b[102])^(a[35] & b[103])^(a[34] & b[104])^(a[33] & b[105])^(a[32] & b[106])^(a[31] & b[107])^(a[30] & b[108])^(a[29] & b[109])^(a[28] & b[110])^(a[27] & b[111])^(a[26] & b[112])^(a[25] & b[113])^(a[24] & b[114])^(a[23] & b[115])^(a[22] & b[116])^(a[21] & b[117])^(a[20] & b[118])^(a[19] & b[119])^(a[18] & b[120])^(a[17] & b[121])^(a[16] & b[122])^(a[15] & b[123])^(a[14] & b[124])^(a[13] & b[125])^(a[12] & b[126])^(a[11] & b[127])^(a[10] & b[128])^(a[9] & b[129])^(a[8] & b[130])^(a[7] & b[131])^(a[6] & b[132])^(a[5] & b[133])^(a[4] & b[134])^(a[3] & b[135])^(a[2] & b[136])^(a[1] & b[137])^(a[0] & b[138]);
assign y[139] = (a[139] & b[0])^(a[138] & b[1])^(a[137] & b[2])^(a[136] & b[3])^(a[135] & b[4])^(a[134] & b[5])^(a[133] & b[6])^(a[132] & b[7])^(a[131] & b[8])^(a[130] & b[9])^(a[129] & b[10])^(a[128] & b[11])^(a[127] & b[12])^(a[126] & b[13])^(a[125] & b[14])^(a[124] & b[15])^(a[123] & b[16])^(a[122] & b[17])^(a[121] & b[18])^(a[120] & b[19])^(a[119] & b[20])^(a[118] & b[21])^(a[117] & b[22])^(a[116] & b[23])^(a[115] & b[24])^(a[114] & b[25])^(a[113] & b[26])^(a[112] & b[27])^(a[111] & b[28])^(a[110] & b[29])^(a[109] & b[30])^(a[108] & b[31])^(a[107] & b[32])^(a[106] & b[33])^(a[105] & b[34])^(a[104] & b[35])^(a[103] & b[36])^(a[102] & b[37])^(a[101] & b[38])^(a[100] & b[39])^(a[99] & b[40])^(a[98] & b[41])^(a[97] & b[42])^(a[96] & b[43])^(a[95] & b[44])^(a[94] & b[45])^(a[93] & b[46])^(a[92] & b[47])^(a[91] & b[48])^(a[90] & b[49])^(a[89] & b[50])^(a[88] & b[51])^(a[87] & b[52])^(a[86] & b[53])^(a[85] & b[54])^(a[84] & b[55])^(a[83] & b[56])^(a[82] & b[57])^(a[81] & b[58])^(a[80] & b[59])^(a[79] & b[60])^(a[78] & b[61])^(a[77] & b[62])^(a[76] & b[63])^(a[75] & b[64])^(a[74] & b[65])^(a[73] & b[66])^(a[72] & b[67])^(a[71] & b[68])^(a[70] & b[69])^(a[69] & b[70])^(a[68] & b[71])^(a[67] & b[72])^(a[66] & b[73])^(a[65] & b[74])^(a[64] & b[75])^(a[63] & b[76])^(a[62] & b[77])^(a[61] & b[78])^(a[60] & b[79])^(a[59] & b[80])^(a[58] & b[81])^(a[57] & b[82])^(a[56] & b[83])^(a[55] & b[84])^(a[54] & b[85])^(a[53] & b[86])^(a[52] & b[87])^(a[51] & b[88])^(a[50] & b[89])^(a[49] & b[90])^(a[48] & b[91])^(a[47] & b[92])^(a[46] & b[93])^(a[45] & b[94])^(a[44] & b[95])^(a[43] & b[96])^(a[42] & b[97])^(a[41] & b[98])^(a[40] & b[99])^(a[39] & b[100])^(a[38] & b[101])^(a[37] & b[102])^(a[36] & b[103])^(a[35] & b[104])^(a[34] & b[105])^(a[33] & b[106])^(a[32] & b[107])^(a[31] & b[108])^(a[30] & b[109])^(a[29] & b[110])^(a[28] & b[111])^(a[27] & b[112])^(a[26] & b[113])^(a[25] & b[114])^(a[24] & b[115])^(a[23] & b[116])^(a[22] & b[117])^(a[21] & b[118])^(a[20] & b[119])^(a[19] & b[120])^(a[18] & b[121])^(a[17] & b[122])^(a[16] & b[123])^(a[15] & b[124])^(a[14] & b[125])^(a[13] & b[126])^(a[12] & b[127])^(a[11] & b[128])^(a[10] & b[129])^(a[9] & b[130])^(a[8] & b[131])^(a[7] & b[132])^(a[6] & b[133])^(a[5] & b[134])^(a[4] & b[135])^(a[3] & b[136])^(a[2] & b[137])^(a[1] & b[138])^(a[0] & b[139]);
assign y[140] = (a[140] & b[0])^(a[139] & b[1])^(a[138] & b[2])^(a[137] & b[3])^(a[136] & b[4])^(a[135] & b[5])^(a[134] & b[6])^(a[133] & b[7])^(a[132] & b[8])^(a[131] & b[9])^(a[130] & b[10])^(a[129] & b[11])^(a[128] & b[12])^(a[127] & b[13])^(a[126] & b[14])^(a[125] & b[15])^(a[124] & b[16])^(a[123] & b[17])^(a[122] & b[18])^(a[121] & b[19])^(a[120] & b[20])^(a[119] & b[21])^(a[118] & b[22])^(a[117] & b[23])^(a[116] & b[24])^(a[115] & b[25])^(a[114] & b[26])^(a[113] & b[27])^(a[112] & b[28])^(a[111] & b[29])^(a[110] & b[30])^(a[109] & b[31])^(a[108] & b[32])^(a[107] & b[33])^(a[106] & b[34])^(a[105] & b[35])^(a[104] & b[36])^(a[103] & b[37])^(a[102] & b[38])^(a[101] & b[39])^(a[100] & b[40])^(a[99] & b[41])^(a[98] & b[42])^(a[97] & b[43])^(a[96] & b[44])^(a[95] & b[45])^(a[94] & b[46])^(a[93] & b[47])^(a[92] & b[48])^(a[91] & b[49])^(a[90] & b[50])^(a[89] & b[51])^(a[88] & b[52])^(a[87] & b[53])^(a[86] & b[54])^(a[85] & b[55])^(a[84] & b[56])^(a[83] & b[57])^(a[82] & b[58])^(a[81] & b[59])^(a[80] & b[60])^(a[79] & b[61])^(a[78] & b[62])^(a[77] & b[63])^(a[76] & b[64])^(a[75] & b[65])^(a[74] & b[66])^(a[73] & b[67])^(a[72] & b[68])^(a[71] & b[69])^(a[70] & b[70])^(a[69] & b[71])^(a[68] & b[72])^(a[67] & b[73])^(a[66] & b[74])^(a[65] & b[75])^(a[64] & b[76])^(a[63] & b[77])^(a[62] & b[78])^(a[61] & b[79])^(a[60] & b[80])^(a[59] & b[81])^(a[58] & b[82])^(a[57] & b[83])^(a[56] & b[84])^(a[55] & b[85])^(a[54] & b[86])^(a[53] & b[87])^(a[52] & b[88])^(a[51] & b[89])^(a[50] & b[90])^(a[49] & b[91])^(a[48] & b[92])^(a[47] & b[93])^(a[46] & b[94])^(a[45] & b[95])^(a[44] & b[96])^(a[43] & b[97])^(a[42] & b[98])^(a[41] & b[99])^(a[40] & b[100])^(a[39] & b[101])^(a[38] & b[102])^(a[37] & b[103])^(a[36] & b[104])^(a[35] & b[105])^(a[34] & b[106])^(a[33] & b[107])^(a[32] & b[108])^(a[31] & b[109])^(a[30] & b[110])^(a[29] & b[111])^(a[28] & b[112])^(a[27] & b[113])^(a[26] & b[114])^(a[25] & b[115])^(a[24] & b[116])^(a[23] & b[117])^(a[22] & b[118])^(a[21] & b[119])^(a[20] & b[120])^(a[19] & b[121])^(a[18] & b[122])^(a[17] & b[123])^(a[16] & b[124])^(a[15] & b[125])^(a[14] & b[126])^(a[13] & b[127])^(a[12] & b[128])^(a[11] & b[129])^(a[10] & b[130])^(a[9] & b[131])^(a[8] & b[132])^(a[7] & b[133])^(a[6] & b[134])^(a[5] & b[135])^(a[4] & b[136])^(a[3] & b[137])^(a[2] & b[138])^(a[1] & b[139])^(a[0] & b[140]);
assign y[141] = (a[141] & b[0])^(a[140] & b[1])^(a[139] & b[2])^(a[138] & b[3])^(a[137] & b[4])^(a[136] & b[5])^(a[135] & b[6])^(a[134] & b[7])^(a[133] & b[8])^(a[132] & b[9])^(a[131] & b[10])^(a[130] & b[11])^(a[129] & b[12])^(a[128] & b[13])^(a[127] & b[14])^(a[126] & b[15])^(a[125] & b[16])^(a[124] & b[17])^(a[123] & b[18])^(a[122] & b[19])^(a[121] & b[20])^(a[120] & b[21])^(a[119] & b[22])^(a[118] & b[23])^(a[117] & b[24])^(a[116] & b[25])^(a[115] & b[26])^(a[114] & b[27])^(a[113] & b[28])^(a[112] & b[29])^(a[111] & b[30])^(a[110] & b[31])^(a[109] & b[32])^(a[108] & b[33])^(a[107] & b[34])^(a[106] & b[35])^(a[105] & b[36])^(a[104] & b[37])^(a[103] & b[38])^(a[102] & b[39])^(a[101] & b[40])^(a[100] & b[41])^(a[99] & b[42])^(a[98] & b[43])^(a[97] & b[44])^(a[96] & b[45])^(a[95] & b[46])^(a[94] & b[47])^(a[93] & b[48])^(a[92] & b[49])^(a[91] & b[50])^(a[90] & b[51])^(a[89] & b[52])^(a[88] & b[53])^(a[87] & b[54])^(a[86] & b[55])^(a[85] & b[56])^(a[84] & b[57])^(a[83] & b[58])^(a[82] & b[59])^(a[81] & b[60])^(a[80] & b[61])^(a[79] & b[62])^(a[78] & b[63])^(a[77] & b[64])^(a[76] & b[65])^(a[75] & b[66])^(a[74] & b[67])^(a[73] & b[68])^(a[72] & b[69])^(a[71] & b[70])^(a[70] & b[71])^(a[69] & b[72])^(a[68] & b[73])^(a[67] & b[74])^(a[66] & b[75])^(a[65] & b[76])^(a[64] & b[77])^(a[63] & b[78])^(a[62] & b[79])^(a[61] & b[80])^(a[60] & b[81])^(a[59] & b[82])^(a[58] & b[83])^(a[57] & b[84])^(a[56] & b[85])^(a[55] & b[86])^(a[54] & b[87])^(a[53] & b[88])^(a[52] & b[89])^(a[51] & b[90])^(a[50] & b[91])^(a[49] & b[92])^(a[48] & b[93])^(a[47] & b[94])^(a[46] & b[95])^(a[45] & b[96])^(a[44] & b[97])^(a[43] & b[98])^(a[42] & b[99])^(a[41] & b[100])^(a[40] & b[101])^(a[39] & b[102])^(a[38] & b[103])^(a[37] & b[104])^(a[36] & b[105])^(a[35] & b[106])^(a[34] & b[107])^(a[33] & b[108])^(a[32] & b[109])^(a[31] & b[110])^(a[30] & b[111])^(a[29] & b[112])^(a[28] & b[113])^(a[27] & b[114])^(a[26] & b[115])^(a[25] & b[116])^(a[24] & b[117])^(a[23] & b[118])^(a[22] & b[119])^(a[21] & b[120])^(a[20] & b[121])^(a[19] & b[122])^(a[18] & b[123])^(a[17] & b[124])^(a[16] & b[125])^(a[15] & b[126])^(a[14] & b[127])^(a[13] & b[128])^(a[12] & b[129])^(a[11] & b[130])^(a[10] & b[131])^(a[9] & b[132])^(a[8] & b[133])^(a[7] & b[134])^(a[6] & b[135])^(a[5] & b[136])^(a[4] & b[137])^(a[3] & b[138])^(a[2] & b[139])^(a[1] & b[140])^(a[0] & b[141]);
assign y[142] = (a[142] & b[0])^(a[141] & b[1])^(a[140] & b[2])^(a[139] & b[3])^(a[138] & b[4])^(a[137] & b[5])^(a[136] & b[6])^(a[135] & b[7])^(a[134] & b[8])^(a[133] & b[9])^(a[132] & b[10])^(a[131] & b[11])^(a[130] & b[12])^(a[129] & b[13])^(a[128] & b[14])^(a[127] & b[15])^(a[126] & b[16])^(a[125] & b[17])^(a[124] & b[18])^(a[123] & b[19])^(a[122] & b[20])^(a[121] & b[21])^(a[120] & b[22])^(a[119] & b[23])^(a[118] & b[24])^(a[117] & b[25])^(a[116] & b[26])^(a[115] & b[27])^(a[114] & b[28])^(a[113] & b[29])^(a[112] & b[30])^(a[111] & b[31])^(a[110] & b[32])^(a[109] & b[33])^(a[108] & b[34])^(a[107] & b[35])^(a[106] & b[36])^(a[105] & b[37])^(a[104] & b[38])^(a[103] & b[39])^(a[102] & b[40])^(a[101] & b[41])^(a[100] & b[42])^(a[99] & b[43])^(a[98] & b[44])^(a[97] & b[45])^(a[96] & b[46])^(a[95] & b[47])^(a[94] & b[48])^(a[93] & b[49])^(a[92] & b[50])^(a[91] & b[51])^(a[90] & b[52])^(a[89] & b[53])^(a[88] & b[54])^(a[87] & b[55])^(a[86] & b[56])^(a[85] & b[57])^(a[84] & b[58])^(a[83] & b[59])^(a[82] & b[60])^(a[81] & b[61])^(a[80] & b[62])^(a[79] & b[63])^(a[78] & b[64])^(a[77] & b[65])^(a[76] & b[66])^(a[75] & b[67])^(a[74] & b[68])^(a[73] & b[69])^(a[72] & b[70])^(a[71] & b[71])^(a[70] & b[72])^(a[69] & b[73])^(a[68] & b[74])^(a[67] & b[75])^(a[66] & b[76])^(a[65] & b[77])^(a[64] & b[78])^(a[63] & b[79])^(a[62] & b[80])^(a[61] & b[81])^(a[60] & b[82])^(a[59] & b[83])^(a[58] & b[84])^(a[57] & b[85])^(a[56] & b[86])^(a[55] & b[87])^(a[54] & b[88])^(a[53] & b[89])^(a[52] & b[90])^(a[51] & b[91])^(a[50] & b[92])^(a[49] & b[93])^(a[48] & b[94])^(a[47] & b[95])^(a[46] & b[96])^(a[45] & b[97])^(a[44] & b[98])^(a[43] & b[99])^(a[42] & b[100])^(a[41] & b[101])^(a[40] & b[102])^(a[39] & b[103])^(a[38] & b[104])^(a[37] & b[105])^(a[36] & b[106])^(a[35] & b[107])^(a[34] & b[108])^(a[33] & b[109])^(a[32] & b[110])^(a[31] & b[111])^(a[30] & b[112])^(a[29] & b[113])^(a[28] & b[114])^(a[27] & b[115])^(a[26] & b[116])^(a[25] & b[117])^(a[24] & b[118])^(a[23] & b[119])^(a[22] & b[120])^(a[21] & b[121])^(a[20] & b[122])^(a[19] & b[123])^(a[18] & b[124])^(a[17] & b[125])^(a[16] & b[126])^(a[15] & b[127])^(a[14] & b[128])^(a[13] & b[129])^(a[12] & b[130])^(a[11] & b[131])^(a[10] & b[132])^(a[9] & b[133])^(a[8] & b[134])^(a[7] & b[135])^(a[6] & b[136])^(a[5] & b[137])^(a[4] & b[138])^(a[3] & b[139])^(a[2] & b[140])^(a[1] & b[141])^(a[0] & b[142]);
assign y[143] = (a[143] & b[0])^(a[142] & b[1])^(a[141] & b[2])^(a[140] & b[3])^(a[139] & b[4])^(a[138] & b[5])^(a[137] & b[6])^(a[136] & b[7])^(a[135] & b[8])^(a[134] & b[9])^(a[133] & b[10])^(a[132] & b[11])^(a[131] & b[12])^(a[130] & b[13])^(a[129] & b[14])^(a[128] & b[15])^(a[127] & b[16])^(a[126] & b[17])^(a[125] & b[18])^(a[124] & b[19])^(a[123] & b[20])^(a[122] & b[21])^(a[121] & b[22])^(a[120] & b[23])^(a[119] & b[24])^(a[118] & b[25])^(a[117] & b[26])^(a[116] & b[27])^(a[115] & b[28])^(a[114] & b[29])^(a[113] & b[30])^(a[112] & b[31])^(a[111] & b[32])^(a[110] & b[33])^(a[109] & b[34])^(a[108] & b[35])^(a[107] & b[36])^(a[106] & b[37])^(a[105] & b[38])^(a[104] & b[39])^(a[103] & b[40])^(a[102] & b[41])^(a[101] & b[42])^(a[100] & b[43])^(a[99] & b[44])^(a[98] & b[45])^(a[97] & b[46])^(a[96] & b[47])^(a[95] & b[48])^(a[94] & b[49])^(a[93] & b[50])^(a[92] & b[51])^(a[91] & b[52])^(a[90] & b[53])^(a[89] & b[54])^(a[88] & b[55])^(a[87] & b[56])^(a[86] & b[57])^(a[85] & b[58])^(a[84] & b[59])^(a[83] & b[60])^(a[82] & b[61])^(a[81] & b[62])^(a[80] & b[63])^(a[79] & b[64])^(a[78] & b[65])^(a[77] & b[66])^(a[76] & b[67])^(a[75] & b[68])^(a[74] & b[69])^(a[73] & b[70])^(a[72] & b[71])^(a[71] & b[72])^(a[70] & b[73])^(a[69] & b[74])^(a[68] & b[75])^(a[67] & b[76])^(a[66] & b[77])^(a[65] & b[78])^(a[64] & b[79])^(a[63] & b[80])^(a[62] & b[81])^(a[61] & b[82])^(a[60] & b[83])^(a[59] & b[84])^(a[58] & b[85])^(a[57] & b[86])^(a[56] & b[87])^(a[55] & b[88])^(a[54] & b[89])^(a[53] & b[90])^(a[52] & b[91])^(a[51] & b[92])^(a[50] & b[93])^(a[49] & b[94])^(a[48] & b[95])^(a[47] & b[96])^(a[46] & b[97])^(a[45] & b[98])^(a[44] & b[99])^(a[43] & b[100])^(a[42] & b[101])^(a[41] & b[102])^(a[40] & b[103])^(a[39] & b[104])^(a[38] & b[105])^(a[37] & b[106])^(a[36] & b[107])^(a[35] & b[108])^(a[34] & b[109])^(a[33] & b[110])^(a[32] & b[111])^(a[31] & b[112])^(a[30] & b[113])^(a[29] & b[114])^(a[28] & b[115])^(a[27] & b[116])^(a[26] & b[117])^(a[25] & b[118])^(a[24] & b[119])^(a[23] & b[120])^(a[22] & b[121])^(a[21] & b[122])^(a[20] & b[123])^(a[19] & b[124])^(a[18] & b[125])^(a[17] & b[126])^(a[16] & b[127])^(a[15] & b[128])^(a[14] & b[129])^(a[13] & b[130])^(a[12] & b[131])^(a[11] & b[132])^(a[10] & b[133])^(a[9] & b[134])^(a[8] & b[135])^(a[7] & b[136])^(a[6] & b[137])^(a[5] & b[138])^(a[4] & b[139])^(a[3] & b[140])^(a[2] & b[141])^(a[1] & b[142])^(a[0] & b[143]);
assign y[144] = (a[144] & b[0])^(a[143] & b[1])^(a[142] & b[2])^(a[141] & b[3])^(a[140] & b[4])^(a[139] & b[5])^(a[138] & b[6])^(a[137] & b[7])^(a[136] & b[8])^(a[135] & b[9])^(a[134] & b[10])^(a[133] & b[11])^(a[132] & b[12])^(a[131] & b[13])^(a[130] & b[14])^(a[129] & b[15])^(a[128] & b[16])^(a[127] & b[17])^(a[126] & b[18])^(a[125] & b[19])^(a[124] & b[20])^(a[123] & b[21])^(a[122] & b[22])^(a[121] & b[23])^(a[120] & b[24])^(a[119] & b[25])^(a[118] & b[26])^(a[117] & b[27])^(a[116] & b[28])^(a[115] & b[29])^(a[114] & b[30])^(a[113] & b[31])^(a[112] & b[32])^(a[111] & b[33])^(a[110] & b[34])^(a[109] & b[35])^(a[108] & b[36])^(a[107] & b[37])^(a[106] & b[38])^(a[105] & b[39])^(a[104] & b[40])^(a[103] & b[41])^(a[102] & b[42])^(a[101] & b[43])^(a[100] & b[44])^(a[99] & b[45])^(a[98] & b[46])^(a[97] & b[47])^(a[96] & b[48])^(a[95] & b[49])^(a[94] & b[50])^(a[93] & b[51])^(a[92] & b[52])^(a[91] & b[53])^(a[90] & b[54])^(a[89] & b[55])^(a[88] & b[56])^(a[87] & b[57])^(a[86] & b[58])^(a[85] & b[59])^(a[84] & b[60])^(a[83] & b[61])^(a[82] & b[62])^(a[81] & b[63])^(a[80] & b[64])^(a[79] & b[65])^(a[78] & b[66])^(a[77] & b[67])^(a[76] & b[68])^(a[75] & b[69])^(a[74] & b[70])^(a[73] & b[71])^(a[72] & b[72])^(a[71] & b[73])^(a[70] & b[74])^(a[69] & b[75])^(a[68] & b[76])^(a[67] & b[77])^(a[66] & b[78])^(a[65] & b[79])^(a[64] & b[80])^(a[63] & b[81])^(a[62] & b[82])^(a[61] & b[83])^(a[60] & b[84])^(a[59] & b[85])^(a[58] & b[86])^(a[57] & b[87])^(a[56] & b[88])^(a[55] & b[89])^(a[54] & b[90])^(a[53] & b[91])^(a[52] & b[92])^(a[51] & b[93])^(a[50] & b[94])^(a[49] & b[95])^(a[48] & b[96])^(a[47] & b[97])^(a[46] & b[98])^(a[45] & b[99])^(a[44] & b[100])^(a[43] & b[101])^(a[42] & b[102])^(a[41] & b[103])^(a[40] & b[104])^(a[39] & b[105])^(a[38] & b[106])^(a[37] & b[107])^(a[36] & b[108])^(a[35] & b[109])^(a[34] & b[110])^(a[33] & b[111])^(a[32] & b[112])^(a[31] & b[113])^(a[30] & b[114])^(a[29] & b[115])^(a[28] & b[116])^(a[27] & b[117])^(a[26] & b[118])^(a[25] & b[119])^(a[24] & b[120])^(a[23] & b[121])^(a[22] & b[122])^(a[21] & b[123])^(a[20] & b[124])^(a[19] & b[125])^(a[18] & b[126])^(a[17] & b[127])^(a[16] & b[128])^(a[15] & b[129])^(a[14] & b[130])^(a[13] & b[131])^(a[12] & b[132])^(a[11] & b[133])^(a[10] & b[134])^(a[9] & b[135])^(a[8] & b[136])^(a[7] & b[137])^(a[6] & b[138])^(a[5] & b[139])^(a[4] & b[140])^(a[3] & b[141])^(a[2] & b[142])^(a[1] & b[143])^(a[0] & b[144]);
assign y[145] = (a[145] & b[0])^(a[144] & b[1])^(a[143] & b[2])^(a[142] & b[3])^(a[141] & b[4])^(a[140] & b[5])^(a[139] & b[6])^(a[138] & b[7])^(a[137] & b[8])^(a[136] & b[9])^(a[135] & b[10])^(a[134] & b[11])^(a[133] & b[12])^(a[132] & b[13])^(a[131] & b[14])^(a[130] & b[15])^(a[129] & b[16])^(a[128] & b[17])^(a[127] & b[18])^(a[126] & b[19])^(a[125] & b[20])^(a[124] & b[21])^(a[123] & b[22])^(a[122] & b[23])^(a[121] & b[24])^(a[120] & b[25])^(a[119] & b[26])^(a[118] & b[27])^(a[117] & b[28])^(a[116] & b[29])^(a[115] & b[30])^(a[114] & b[31])^(a[113] & b[32])^(a[112] & b[33])^(a[111] & b[34])^(a[110] & b[35])^(a[109] & b[36])^(a[108] & b[37])^(a[107] & b[38])^(a[106] & b[39])^(a[105] & b[40])^(a[104] & b[41])^(a[103] & b[42])^(a[102] & b[43])^(a[101] & b[44])^(a[100] & b[45])^(a[99] & b[46])^(a[98] & b[47])^(a[97] & b[48])^(a[96] & b[49])^(a[95] & b[50])^(a[94] & b[51])^(a[93] & b[52])^(a[92] & b[53])^(a[91] & b[54])^(a[90] & b[55])^(a[89] & b[56])^(a[88] & b[57])^(a[87] & b[58])^(a[86] & b[59])^(a[85] & b[60])^(a[84] & b[61])^(a[83] & b[62])^(a[82] & b[63])^(a[81] & b[64])^(a[80] & b[65])^(a[79] & b[66])^(a[78] & b[67])^(a[77] & b[68])^(a[76] & b[69])^(a[75] & b[70])^(a[74] & b[71])^(a[73] & b[72])^(a[72] & b[73])^(a[71] & b[74])^(a[70] & b[75])^(a[69] & b[76])^(a[68] & b[77])^(a[67] & b[78])^(a[66] & b[79])^(a[65] & b[80])^(a[64] & b[81])^(a[63] & b[82])^(a[62] & b[83])^(a[61] & b[84])^(a[60] & b[85])^(a[59] & b[86])^(a[58] & b[87])^(a[57] & b[88])^(a[56] & b[89])^(a[55] & b[90])^(a[54] & b[91])^(a[53] & b[92])^(a[52] & b[93])^(a[51] & b[94])^(a[50] & b[95])^(a[49] & b[96])^(a[48] & b[97])^(a[47] & b[98])^(a[46] & b[99])^(a[45] & b[100])^(a[44] & b[101])^(a[43] & b[102])^(a[42] & b[103])^(a[41] & b[104])^(a[40] & b[105])^(a[39] & b[106])^(a[38] & b[107])^(a[37] & b[108])^(a[36] & b[109])^(a[35] & b[110])^(a[34] & b[111])^(a[33] & b[112])^(a[32] & b[113])^(a[31] & b[114])^(a[30] & b[115])^(a[29] & b[116])^(a[28] & b[117])^(a[27] & b[118])^(a[26] & b[119])^(a[25] & b[120])^(a[24] & b[121])^(a[23] & b[122])^(a[22] & b[123])^(a[21] & b[124])^(a[20] & b[125])^(a[19] & b[126])^(a[18] & b[127])^(a[17] & b[128])^(a[16] & b[129])^(a[15] & b[130])^(a[14] & b[131])^(a[13] & b[132])^(a[12] & b[133])^(a[11] & b[134])^(a[10] & b[135])^(a[9] & b[136])^(a[8] & b[137])^(a[7] & b[138])^(a[6] & b[139])^(a[5] & b[140])^(a[4] & b[141])^(a[3] & b[142])^(a[2] & b[143])^(a[1] & b[144])^(a[0] & b[145]);
assign y[146] = (a[146] & b[0])^(a[145] & b[1])^(a[144] & b[2])^(a[143] & b[3])^(a[142] & b[4])^(a[141] & b[5])^(a[140] & b[6])^(a[139] & b[7])^(a[138] & b[8])^(a[137] & b[9])^(a[136] & b[10])^(a[135] & b[11])^(a[134] & b[12])^(a[133] & b[13])^(a[132] & b[14])^(a[131] & b[15])^(a[130] & b[16])^(a[129] & b[17])^(a[128] & b[18])^(a[127] & b[19])^(a[126] & b[20])^(a[125] & b[21])^(a[124] & b[22])^(a[123] & b[23])^(a[122] & b[24])^(a[121] & b[25])^(a[120] & b[26])^(a[119] & b[27])^(a[118] & b[28])^(a[117] & b[29])^(a[116] & b[30])^(a[115] & b[31])^(a[114] & b[32])^(a[113] & b[33])^(a[112] & b[34])^(a[111] & b[35])^(a[110] & b[36])^(a[109] & b[37])^(a[108] & b[38])^(a[107] & b[39])^(a[106] & b[40])^(a[105] & b[41])^(a[104] & b[42])^(a[103] & b[43])^(a[102] & b[44])^(a[101] & b[45])^(a[100] & b[46])^(a[99] & b[47])^(a[98] & b[48])^(a[97] & b[49])^(a[96] & b[50])^(a[95] & b[51])^(a[94] & b[52])^(a[93] & b[53])^(a[92] & b[54])^(a[91] & b[55])^(a[90] & b[56])^(a[89] & b[57])^(a[88] & b[58])^(a[87] & b[59])^(a[86] & b[60])^(a[85] & b[61])^(a[84] & b[62])^(a[83] & b[63])^(a[82] & b[64])^(a[81] & b[65])^(a[80] & b[66])^(a[79] & b[67])^(a[78] & b[68])^(a[77] & b[69])^(a[76] & b[70])^(a[75] & b[71])^(a[74] & b[72])^(a[73] & b[73])^(a[72] & b[74])^(a[71] & b[75])^(a[70] & b[76])^(a[69] & b[77])^(a[68] & b[78])^(a[67] & b[79])^(a[66] & b[80])^(a[65] & b[81])^(a[64] & b[82])^(a[63] & b[83])^(a[62] & b[84])^(a[61] & b[85])^(a[60] & b[86])^(a[59] & b[87])^(a[58] & b[88])^(a[57] & b[89])^(a[56] & b[90])^(a[55] & b[91])^(a[54] & b[92])^(a[53] & b[93])^(a[52] & b[94])^(a[51] & b[95])^(a[50] & b[96])^(a[49] & b[97])^(a[48] & b[98])^(a[47] & b[99])^(a[46] & b[100])^(a[45] & b[101])^(a[44] & b[102])^(a[43] & b[103])^(a[42] & b[104])^(a[41] & b[105])^(a[40] & b[106])^(a[39] & b[107])^(a[38] & b[108])^(a[37] & b[109])^(a[36] & b[110])^(a[35] & b[111])^(a[34] & b[112])^(a[33] & b[113])^(a[32] & b[114])^(a[31] & b[115])^(a[30] & b[116])^(a[29] & b[117])^(a[28] & b[118])^(a[27] & b[119])^(a[26] & b[120])^(a[25] & b[121])^(a[24] & b[122])^(a[23] & b[123])^(a[22] & b[124])^(a[21] & b[125])^(a[20] & b[126])^(a[19] & b[127])^(a[18] & b[128])^(a[17] & b[129])^(a[16] & b[130])^(a[15] & b[131])^(a[14] & b[132])^(a[13] & b[133])^(a[12] & b[134])^(a[11] & b[135])^(a[10] & b[136])^(a[9] & b[137])^(a[8] & b[138])^(a[7] & b[139])^(a[6] & b[140])^(a[5] & b[141])^(a[4] & b[142])^(a[3] & b[143])^(a[2] & b[144])^(a[1] & b[145])^(a[0] & b[146]);
assign y[147] = (a[147] & b[0])^(a[146] & b[1])^(a[145] & b[2])^(a[144] & b[3])^(a[143] & b[4])^(a[142] & b[5])^(a[141] & b[6])^(a[140] & b[7])^(a[139] & b[8])^(a[138] & b[9])^(a[137] & b[10])^(a[136] & b[11])^(a[135] & b[12])^(a[134] & b[13])^(a[133] & b[14])^(a[132] & b[15])^(a[131] & b[16])^(a[130] & b[17])^(a[129] & b[18])^(a[128] & b[19])^(a[127] & b[20])^(a[126] & b[21])^(a[125] & b[22])^(a[124] & b[23])^(a[123] & b[24])^(a[122] & b[25])^(a[121] & b[26])^(a[120] & b[27])^(a[119] & b[28])^(a[118] & b[29])^(a[117] & b[30])^(a[116] & b[31])^(a[115] & b[32])^(a[114] & b[33])^(a[113] & b[34])^(a[112] & b[35])^(a[111] & b[36])^(a[110] & b[37])^(a[109] & b[38])^(a[108] & b[39])^(a[107] & b[40])^(a[106] & b[41])^(a[105] & b[42])^(a[104] & b[43])^(a[103] & b[44])^(a[102] & b[45])^(a[101] & b[46])^(a[100] & b[47])^(a[99] & b[48])^(a[98] & b[49])^(a[97] & b[50])^(a[96] & b[51])^(a[95] & b[52])^(a[94] & b[53])^(a[93] & b[54])^(a[92] & b[55])^(a[91] & b[56])^(a[90] & b[57])^(a[89] & b[58])^(a[88] & b[59])^(a[87] & b[60])^(a[86] & b[61])^(a[85] & b[62])^(a[84] & b[63])^(a[83] & b[64])^(a[82] & b[65])^(a[81] & b[66])^(a[80] & b[67])^(a[79] & b[68])^(a[78] & b[69])^(a[77] & b[70])^(a[76] & b[71])^(a[75] & b[72])^(a[74] & b[73])^(a[73] & b[74])^(a[72] & b[75])^(a[71] & b[76])^(a[70] & b[77])^(a[69] & b[78])^(a[68] & b[79])^(a[67] & b[80])^(a[66] & b[81])^(a[65] & b[82])^(a[64] & b[83])^(a[63] & b[84])^(a[62] & b[85])^(a[61] & b[86])^(a[60] & b[87])^(a[59] & b[88])^(a[58] & b[89])^(a[57] & b[90])^(a[56] & b[91])^(a[55] & b[92])^(a[54] & b[93])^(a[53] & b[94])^(a[52] & b[95])^(a[51] & b[96])^(a[50] & b[97])^(a[49] & b[98])^(a[48] & b[99])^(a[47] & b[100])^(a[46] & b[101])^(a[45] & b[102])^(a[44] & b[103])^(a[43] & b[104])^(a[42] & b[105])^(a[41] & b[106])^(a[40] & b[107])^(a[39] & b[108])^(a[38] & b[109])^(a[37] & b[110])^(a[36] & b[111])^(a[35] & b[112])^(a[34] & b[113])^(a[33] & b[114])^(a[32] & b[115])^(a[31] & b[116])^(a[30] & b[117])^(a[29] & b[118])^(a[28] & b[119])^(a[27] & b[120])^(a[26] & b[121])^(a[25] & b[122])^(a[24] & b[123])^(a[23] & b[124])^(a[22] & b[125])^(a[21] & b[126])^(a[20] & b[127])^(a[19] & b[128])^(a[18] & b[129])^(a[17] & b[130])^(a[16] & b[131])^(a[15] & b[132])^(a[14] & b[133])^(a[13] & b[134])^(a[12] & b[135])^(a[11] & b[136])^(a[10] & b[137])^(a[9] & b[138])^(a[8] & b[139])^(a[7] & b[140])^(a[6] & b[141])^(a[5] & b[142])^(a[4] & b[143])^(a[3] & b[144])^(a[2] & b[145])^(a[1] & b[146])^(a[0] & b[147]);
assign y[148] = (a[148] & b[0])^(a[147] & b[1])^(a[146] & b[2])^(a[145] & b[3])^(a[144] & b[4])^(a[143] & b[5])^(a[142] & b[6])^(a[141] & b[7])^(a[140] & b[8])^(a[139] & b[9])^(a[138] & b[10])^(a[137] & b[11])^(a[136] & b[12])^(a[135] & b[13])^(a[134] & b[14])^(a[133] & b[15])^(a[132] & b[16])^(a[131] & b[17])^(a[130] & b[18])^(a[129] & b[19])^(a[128] & b[20])^(a[127] & b[21])^(a[126] & b[22])^(a[125] & b[23])^(a[124] & b[24])^(a[123] & b[25])^(a[122] & b[26])^(a[121] & b[27])^(a[120] & b[28])^(a[119] & b[29])^(a[118] & b[30])^(a[117] & b[31])^(a[116] & b[32])^(a[115] & b[33])^(a[114] & b[34])^(a[113] & b[35])^(a[112] & b[36])^(a[111] & b[37])^(a[110] & b[38])^(a[109] & b[39])^(a[108] & b[40])^(a[107] & b[41])^(a[106] & b[42])^(a[105] & b[43])^(a[104] & b[44])^(a[103] & b[45])^(a[102] & b[46])^(a[101] & b[47])^(a[100] & b[48])^(a[99] & b[49])^(a[98] & b[50])^(a[97] & b[51])^(a[96] & b[52])^(a[95] & b[53])^(a[94] & b[54])^(a[93] & b[55])^(a[92] & b[56])^(a[91] & b[57])^(a[90] & b[58])^(a[89] & b[59])^(a[88] & b[60])^(a[87] & b[61])^(a[86] & b[62])^(a[85] & b[63])^(a[84] & b[64])^(a[83] & b[65])^(a[82] & b[66])^(a[81] & b[67])^(a[80] & b[68])^(a[79] & b[69])^(a[78] & b[70])^(a[77] & b[71])^(a[76] & b[72])^(a[75] & b[73])^(a[74] & b[74])^(a[73] & b[75])^(a[72] & b[76])^(a[71] & b[77])^(a[70] & b[78])^(a[69] & b[79])^(a[68] & b[80])^(a[67] & b[81])^(a[66] & b[82])^(a[65] & b[83])^(a[64] & b[84])^(a[63] & b[85])^(a[62] & b[86])^(a[61] & b[87])^(a[60] & b[88])^(a[59] & b[89])^(a[58] & b[90])^(a[57] & b[91])^(a[56] & b[92])^(a[55] & b[93])^(a[54] & b[94])^(a[53] & b[95])^(a[52] & b[96])^(a[51] & b[97])^(a[50] & b[98])^(a[49] & b[99])^(a[48] & b[100])^(a[47] & b[101])^(a[46] & b[102])^(a[45] & b[103])^(a[44] & b[104])^(a[43] & b[105])^(a[42] & b[106])^(a[41] & b[107])^(a[40] & b[108])^(a[39] & b[109])^(a[38] & b[110])^(a[37] & b[111])^(a[36] & b[112])^(a[35] & b[113])^(a[34] & b[114])^(a[33] & b[115])^(a[32] & b[116])^(a[31] & b[117])^(a[30] & b[118])^(a[29] & b[119])^(a[28] & b[120])^(a[27] & b[121])^(a[26] & b[122])^(a[25] & b[123])^(a[24] & b[124])^(a[23] & b[125])^(a[22] & b[126])^(a[21] & b[127])^(a[20] & b[128])^(a[19] & b[129])^(a[18] & b[130])^(a[17] & b[131])^(a[16] & b[132])^(a[15] & b[133])^(a[14] & b[134])^(a[13] & b[135])^(a[12] & b[136])^(a[11] & b[137])^(a[10] & b[138])^(a[9] & b[139])^(a[8] & b[140])^(a[7] & b[141])^(a[6] & b[142])^(a[5] & b[143])^(a[4] & b[144])^(a[3] & b[145])^(a[2] & b[146])^(a[1] & b[147])^(a[0] & b[148]);
assign y[149] = (a[149] & b[0])^(a[148] & b[1])^(a[147] & b[2])^(a[146] & b[3])^(a[145] & b[4])^(a[144] & b[5])^(a[143] & b[6])^(a[142] & b[7])^(a[141] & b[8])^(a[140] & b[9])^(a[139] & b[10])^(a[138] & b[11])^(a[137] & b[12])^(a[136] & b[13])^(a[135] & b[14])^(a[134] & b[15])^(a[133] & b[16])^(a[132] & b[17])^(a[131] & b[18])^(a[130] & b[19])^(a[129] & b[20])^(a[128] & b[21])^(a[127] & b[22])^(a[126] & b[23])^(a[125] & b[24])^(a[124] & b[25])^(a[123] & b[26])^(a[122] & b[27])^(a[121] & b[28])^(a[120] & b[29])^(a[119] & b[30])^(a[118] & b[31])^(a[117] & b[32])^(a[116] & b[33])^(a[115] & b[34])^(a[114] & b[35])^(a[113] & b[36])^(a[112] & b[37])^(a[111] & b[38])^(a[110] & b[39])^(a[109] & b[40])^(a[108] & b[41])^(a[107] & b[42])^(a[106] & b[43])^(a[105] & b[44])^(a[104] & b[45])^(a[103] & b[46])^(a[102] & b[47])^(a[101] & b[48])^(a[100] & b[49])^(a[99] & b[50])^(a[98] & b[51])^(a[97] & b[52])^(a[96] & b[53])^(a[95] & b[54])^(a[94] & b[55])^(a[93] & b[56])^(a[92] & b[57])^(a[91] & b[58])^(a[90] & b[59])^(a[89] & b[60])^(a[88] & b[61])^(a[87] & b[62])^(a[86] & b[63])^(a[85] & b[64])^(a[84] & b[65])^(a[83] & b[66])^(a[82] & b[67])^(a[81] & b[68])^(a[80] & b[69])^(a[79] & b[70])^(a[78] & b[71])^(a[77] & b[72])^(a[76] & b[73])^(a[75] & b[74])^(a[74] & b[75])^(a[73] & b[76])^(a[72] & b[77])^(a[71] & b[78])^(a[70] & b[79])^(a[69] & b[80])^(a[68] & b[81])^(a[67] & b[82])^(a[66] & b[83])^(a[65] & b[84])^(a[64] & b[85])^(a[63] & b[86])^(a[62] & b[87])^(a[61] & b[88])^(a[60] & b[89])^(a[59] & b[90])^(a[58] & b[91])^(a[57] & b[92])^(a[56] & b[93])^(a[55] & b[94])^(a[54] & b[95])^(a[53] & b[96])^(a[52] & b[97])^(a[51] & b[98])^(a[50] & b[99])^(a[49] & b[100])^(a[48] & b[101])^(a[47] & b[102])^(a[46] & b[103])^(a[45] & b[104])^(a[44] & b[105])^(a[43] & b[106])^(a[42] & b[107])^(a[41] & b[108])^(a[40] & b[109])^(a[39] & b[110])^(a[38] & b[111])^(a[37] & b[112])^(a[36] & b[113])^(a[35] & b[114])^(a[34] & b[115])^(a[33] & b[116])^(a[32] & b[117])^(a[31] & b[118])^(a[30] & b[119])^(a[29] & b[120])^(a[28] & b[121])^(a[27] & b[122])^(a[26] & b[123])^(a[25] & b[124])^(a[24] & b[125])^(a[23] & b[126])^(a[22] & b[127])^(a[21] & b[128])^(a[20] & b[129])^(a[19] & b[130])^(a[18] & b[131])^(a[17] & b[132])^(a[16] & b[133])^(a[15] & b[134])^(a[14] & b[135])^(a[13] & b[136])^(a[12] & b[137])^(a[11] & b[138])^(a[10] & b[139])^(a[9] & b[140])^(a[8] & b[141])^(a[7] & b[142])^(a[6] & b[143])^(a[5] & b[144])^(a[4] & b[145])^(a[3] & b[146])^(a[2] & b[147])^(a[1] & b[148])^(a[0] & b[149]);
assign y[150] = (a[150] & b[0])^(a[149] & b[1])^(a[148] & b[2])^(a[147] & b[3])^(a[146] & b[4])^(a[145] & b[5])^(a[144] & b[6])^(a[143] & b[7])^(a[142] & b[8])^(a[141] & b[9])^(a[140] & b[10])^(a[139] & b[11])^(a[138] & b[12])^(a[137] & b[13])^(a[136] & b[14])^(a[135] & b[15])^(a[134] & b[16])^(a[133] & b[17])^(a[132] & b[18])^(a[131] & b[19])^(a[130] & b[20])^(a[129] & b[21])^(a[128] & b[22])^(a[127] & b[23])^(a[126] & b[24])^(a[125] & b[25])^(a[124] & b[26])^(a[123] & b[27])^(a[122] & b[28])^(a[121] & b[29])^(a[120] & b[30])^(a[119] & b[31])^(a[118] & b[32])^(a[117] & b[33])^(a[116] & b[34])^(a[115] & b[35])^(a[114] & b[36])^(a[113] & b[37])^(a[112] & b[38])^(a[111] & b[39])^(a[110] & b[40])^(a[109] & b[41])^(a[108] & b[42])^(a[107] & b[43])^(a[106] & b[44])^(a[105] & b[45])^(a[104] & b[46])^(a[103] & b[47])^(a[102] & b[48])^(a[101] & b[49])^(a[100] & b[50])^(a[99] & b[51])^(a[98] & b[52])^(a[97] & b[53])^(a[96] & b[54])^(a[95] & b[55])^(a[94] & b[56])^(a[93] & b[57])^(a[92] & b[58])^(a[91] & b[59])^(a[90] & b[60])^(a[89] & b[61])^(a[88] & b[62])^(a[87] & b[63])^(a[86] & b[64])^(a[85] & b[65])^(a[84] & b[66])^(a[83] & b[67])^(a[82] & b[68])^(a[81] & b[69])^(a[80] & b[70])^(a[79] & b[71])^(a[78] & b[72])^(a[77] & b[73])^(a[76] & b[74])^(a[75] & b[75])^(a[74] & b[76])^(a[73] & b[77])^(a[72] & b[78])^(a[71] & b[79])^(a[70] & b[80])^(a[69] & b[81])^(a[68] & b[82])^(a[67] & b[83])^(a[66] & b[84])^(a[65] & b[85])^(a[64] & b[86])^(a[63] & b[87])^(a[62] & b[88])^(a[61] & b[89])^(a[60] & b[90])^(a[59] & b[91])^(a[58] & b[92])^(a[57] & b[93])^(a[56] & b[94])^(a[55] & b[95])^(a[54] & b[96])^(a[53] & b[97])^(a[52] & b[98])^(a[51] & b[99])^(a[50] & b[100])^(a[49] & b[101])^(a[48] & b[102])^(a[47] & b[103])^(a[46] & b[104])^(a[45] & b[105])^(a[44] & b[106])^(a[43] & b[107])^(a[42] & b[108])^(a[41] & b[109])^(a[40] & b[110])^(a[39] & b[111])^(a[38] & b[112])^(a[37] & b[113])^(a[36] & b[114])^(a[35] & b[115])^(a[34] & b[116])^(a[33] & b[117])^(a[32] & b[118])^(a[31] & b[119])^(a[30] & b[120])^(a[29] & b[121])^(a[28] & b[122])^(a[27] & b[123])^(a[26] & b[124])^(a[25] & b[125])^(a[24] & b[126])^(a[23] & b[127])^(a[22] & b[128])^(a[21] & b[129])^(a[20] & b[130])^(a[19] & b[131])^(a[18] & b[132])^(a[17] & b[133])^(a[16] & b[134])^(a[15] & b[135])^(a[14] & b[136])^(a[13] & b[137])^(a[12] & b[138])^(a[11] & b[139])^(a[10] & b[140])^(a[9] & b[141])^(a[8] & b[142])^(a[7] & b[143])^(a[6] & b[144])^(a[5] & b[145])^(a[4] & b[146])^(a[3] & b[147])^(a[2] & b[148])^(a[1] & b[149])^(a[0] & b[150]);
assign y[151] = (a[151] & b[0])^(a[150] & b[1])^(a[149] & b[2])^(a[148] & b[3])^(a[147] & b[4])^(a[146] & b[5])^(a[145] & b[6])^(a[144] & b[7])^(a[143] & b[8])^(a[142] & b[9])^(a[141] & b[10])^(a[140] & b[11])^(a[139] & b[12])^(a[138] & b[13])^(a[137] & b[14])^(a[136] & b[15])^(a[135] & b[16])^(a[134] & b[17])^(a[133] & b[18])^(a[132] & b[19])^(a[131] & b[20])^(a[130] & b[21])^(a[129] & b[22])^(a[128] & b[23])^(a[127] & b[24])^(a[126] & b[25])^(a[125] & b[26])^(a[124] & b[27])^(a[123] & b[28])^(a[122] & b[29])^(a[121] & b[30])^(a[120] & b[31])^(a[119] & b[32])^(a[118] & b[33])^(a[117] & b[34])^(a[116] & b[35])^(a[115] & b[36])^(a[114] & b[37])^(a[113] & b[38])^(a[112] & b[39])^(a[111] & b[40])^(a[110] & b[41])^(a[109] & b[42])^(a[108] & b[43])^(a[107] & b[44])^(a[106] & b[45])^(a[105] & b[46])^(a[104] & b[47])^(a[103] & b[48])^(a[102] & b[49])^(a[101] & b[50])^(a[100] & b[51])^(a[99] & b[52])^(a[98] & b[53])^(a[97] & b[54])^(a[96] & b[55])^(a[95] & b[56])^(a[94] & b[57])^(a[93] & b[58])^(a[92] & b[59])^(a[91] & b[60])^(a[90] & b[61])^(a[89] & b[62])^(a[88] & b[63])^(a[87] & b[64])^(a[86] & b[65])^(a[85] & b[66])^(a[84] & b[67])^(a[83] & b[68])^(a[82] & b[69])^(a[81] & b[70])^(a[80] & b[71])^(a[79] & b[72])^(a[78] & b[73])^(a[77] & b[74])^(a[76] & b[75])^(a[75] & b[76])^(a[74] & b[77])^(a[73] & b[78])^(a[72] & b[79])^(a[71] & b[80])^(a[70] & b[81])^(a[69] & b[82])^(a[68] & b[83])^(a[67] & b[84])^(a[66] & b[85])^(a[65] & b[86])^(a[64] & b[87])^(a[63] & b[88])^(a[62] & b[89])^(a[61] & b[90])^(a[60] & b[91])^(a[59] & b[92])^(a[58] & b[93])^(a[57] & b[94])^(a[56] & b[95])^(a[55] & b[96])^(a[54] & b[97])^(a[53] & b[98])^(a[52] & b[99])^(a[51] & b[100])^(a[50] & b[101])^(a[49] & b[102])^(a[48] & b[103])^(a[47] & b[104])^(a[46] & b[105])^(a[45] & b[106])^(a[44] & b[107])^(a[43] & b[108])^(a[42] & b[109])^(a[41] & b[110])^(a[40] & b[111])^(a[39] & b[112])^(a[38] & b[113])^(a[37] & b[114])^(a[36] & b[115])^(a[35] & b[116])^(a[34] & b[117])^(a[33] & b[118])^(a[32] & b[119])^(a[31] & b[120])^(a[30] & b[121])^(a[29] & b[122])^(a[28] & b[123])^(a[27] & b[124])^(a[26] & b[125])^(a[25] & b[126])^(a[24] & b[127])^(a[23] & b[128])^(a[22] & b[129])^(a[21] & b[130])^(a[20] & b[131])^(a[19] & b[132])^(a[18] & b[133])^(a[17] & b[134])^(a[16] & b[135])^(a[15] & b[136])^(a[14] & b[137])^(a[13] & b[138])^(a[12] & b[139])^(a[11] & b[140])^(a[10] & b[141])^(a[9] & b[142])^(a[8] & b[143])^(a[7] & b[144])^(a[6] & b[145])^(a[5] & b[146])^(a[4] & b[147])^(a[3] & b[148])^(a[2] & b[149])^(a[1] & b[150])^(a[0] & b[151]);
assign y[152] = (a[152] & b[0])^(a[151] & b[1])^(a[150] & b[2])^(a[149] & b[3])^(a[148] & b[4])^(a[147] & b[5])^(a[146] & b[6])^(a[145] & b[7])^(a[144] & b[8])^(a[143] & b[9])^(a[142] & b[10])^(a[141] & b[11])^(a[140] & b[12])^(a[139] & b[13])^(a[138] & b[14])^(a[137] & b[15])^(a[136] & b[16])^(a[135] & b[17])^(a[134] & b[18])^(a[133] & b[19])^(a[132] & b[20])^(a[131] & b[21])^(a[130] & b[22])^(a[129] & b[23])^(a[128] & b[24])^(a[127] & b[25])^(a[126] & b[26])^(a[125] & b[27])^(a[124] & b[28])^(a[123] & b[29])^(a[122] & b[30])^(a[121] & b[31])^(a[120] & b[32])^(a[119] & b[33])^(a[118] & b[34])^(a[117] & b[35])^(a[116] & b[36])^(a[115] & b[37])^(a[114] & b[38])^(a[113] & b[39])^(a[112] & b[40])^(a[111] & b[41])^(a[110] & b[42])^(a[109] & b[43])^(a[108] & b[44])^(a[107] & b[45])^(a[106] & b[46])^(a[105] & b[47])^(a[104] & b[48])^(a[103] & b[49])^(a[102] & b[50])^(a[101] & b[51])^(a[100] & b[52])^(a[99] & b[53])^(a[98] & b[54])^(a[97] & b[55])^(a[96] & b[56])^(a[95] & b[57])^(a[94] & b[58])^(a[93] & b[59])^(a[92] & b[60])^(a[91] & b[61])^(a[90] & b[62])^(a[89] & b[63])^(a[88] & b[64])^(a[87] & b[65])^(a[86] & b[66])^(a[85] & b[67])^(a[84] & b[68])^(a[83] & b[69])^(a[82] & b[70])^(a[81] & b[71])^(a[80] & b[72])^(a[79] & b[73])^(a[78] & b[74])^(a[77] & b[75])^(a[76] & b[76])^(a[75] & b[77])^(a[74] & b[78])^(a[73] & b[79])^(a[72] & b[80])^(a[71] & b[81])^(a[70] & b[82])^(a[69] & b[83])^(a[68] & b[84])^(a[67] & b[85])^(a[66] & b[86])^(a[65] & b[87])^(a[64] & b[88])^(a[63] & b[89])^(a[62] & b[90])^(a[61] & b[91])^(a[60] & b[92])^(a[59] & b[93])^(a[58] & b[94])^(a[57] & b[95])^(a[56] & b[96])^(a[55] & b[97])^(a[54] & b[98])^(a[53] & b[99])^(a[52] & b[100])^(a[51] & b[101])^(a[50] & b[102])^(a[49] & b[103])^(a[48] & b[104])^(a[47] & b[105])^(a[46] & b[106])^(a[45] & b[107])^(a[44] & b[108])^(a[43] & b[109])^(a[42] & b[110])^(a[41] & b[111])^(a[40] & b[112])^(a[39] & b[113])^(a[38] & b[114])^(a[37] & b[115])^(a[36] & b[116])^(a[35] & b[117])^(a[34] & b[118])^(a[33] & b[119])^(a[32] & b[120])^(a[31] & b[121])^(a[30] & b[122])^(a[29] & b[123])^(a[28] & b[124])^(a[27] & b[125])^(a[26] & b[126])^(a[25] & b[127])^(a[24] & b[128])^(a[23] & b[129])^(a[22] & b[130])^(a[21] & b[131])^(a[20] & b[132])^(a[19] & b[133])^(a[18] & b[134])^(a[17] & b[135])^(a[16] & b[136])^(a[15] & b[137])^(a[14] & b[138])^(a[13] & b[139])^(a[12] & b[140])^(a[11] & b[141])^(a[10] & b[142])^(a[9] & b[143])^(a[8] & b[144])^(a[7] & b[145])^(a[6] & b[146])^(a[5] & b[147])^(a[4] & b[148])^(a[3] & b[149])^(a[2] & b[150])^(a[1] & b[151])^(a[0] & b[152]);
assign y[153] = (a[153] & b[0])^(a[152] & b[1])^(a[151] & b[2])^(a[150] & b[3])^(a[149] & b[4])^(a[148] & b[5])^(a[147] & b[6])^(a[146] & b[7])^(a[145] & b[8])^(a[144] & b[9])^(a[143] & b[10])^(a[142] & b[11])^(a[141] & b[12])^(a[140] & b[13])^(a[139] & b[14])^(a[138] & b[15])^(a[137] & b[16])^(a[136] & b[17])^(a[135] & b[18])^(a[134] & b[19])^(a[133] & b[20])^(a[132] & b[21])^(a[131] & b[22])^(a[130] & b[23])^(a[129] & b[24])^(a[128] & b[25])^(a[127] & b[26])^(a[126] & b[27])^(a[125] & b[28])^(a[124] & b[29])^(a[123] & b[30])^(a[122] & b[31])^(a[121] & b[32])^(a[120] & b[33])^(a[119] & b[34])^(a[118] & b[35])^(a[117] & b[36])^(a[116] & b[37])^(a[115] & b[38])^(a[114] & b[39])^(a[113] & b[40])^(a[112] & b[41])^(a[111] & b[42])^(a[110] & b[43])^(a[109] & b[44])^(a[108] & b[45])^(a[107] & b[46])^(a[106] & b[47])^(a[105] & b[48])^(a[104] & b[49])^(a[103] & b[50])^(a[102] & b[51])^(a[101] & b[52])^(a[100] & b[53])^(a[99] & b[54])^(a[98] & b[55])^(a[97] & b[56])^(a[96] & b[57])^(a[95] & b[58])^(a[94] & b[59])^(a[93] & b[60])^(a[92] & b[61])^(a[91] & b[62])^(a[90] & b[63])^(a[89] & b[64])^(a[88] & b[65])^(a[87] & b[66])^(a[86] & b[67])^(a[85] & b[68])^(a[84] & b[69])^(a[83] & b[70])^(a[82] & b[71])^(a[81] & b[72])^(a[80] & b[73])^(a[79] & b[74])^(a[78] & b[75])^(a[77] & b[76])^(a[76] & b[77])^(a[75] & b[78])^(a[74] & b[79])^(a[73] & b[80])^(a[72] & b[81])^(a[71] & b[82])^(a[70] & b[83])^(a[69] & b[84])^(a[68] & b[85])^(a[67] & b[86])^(a[66] & b[87])^(a[65] & b[88])^(a[64] & b[89])^(a[63] & b[90])^(a[62] & b[91])^(a[61] & b[92])^(a[60] & b[93])^(a[59] & b[94])^(a[58] & b[95])^(a[57] & b[96])^(a[56] & b[97])^(a[55] & b[98])^(a[54] & b[99])^(a[53] & b[100])^(a[52] & b[101])^(a[51] & b[102])^(a[50] & b[103])^(a[49] & b[104])^(a[48] & b[105])^(a[47] & b[106])^(a[46] & b[107])^(a[45] & b[108])^(a[44] & b[109])^(a[43] & b[110])^(a[42] & b[111])^(a[41] & b[112])^(a[40] & b[113])^(a[39] & b[114])^(a[38] & b[115])^(a[37] & b[116])^(a[36] & b[117])^(a[35] & b[118])^(a[34] & b[119])^(a[33] & b[120])^(a[32] & b[121])^(a[31] & b[122])^(a[30] & b[123])^(a[29] & b[124])^(a[28] & b[125])^(a[27] & b[126])^(a[26] & b[127])^(a[25] & b[128])^(a[24] & b[129])^(a[23] & b[130])^(a[22] & b[131])^(a[21] & b[132])^(a[20] & b[133])^(a[19] & b[134])^(a[18] & b[135])^(a[17] & b[136])^(a[16] & b[137])^(a[15] & b[138])^(a[14] & b[139])^(a[13] & b[140])^(a[12] & b[141])^(a[11] & b[142])^(a[10] & b[143])^(a[9] & b[144])^(a[8] & b[145])^(a[7] & b[146])^(a[6] & b[147])^(a[5] & b[148])^(a[4] & b[149])^(a[3] & b[150])^(a[2] & b[151])^(a[1] & b[152])^(a[0] & b[153]);
assign y[154] = (a[154] & b[0])^(a[153] & b[1])^(a[152] & b[2])^(a[151] & b[3])^(a[150] & b[4])^(a[149] & b[5])^(a[148] & b[6])^(a[147] & b[7])^(a[146] & b[8])^(a[145] & b[9])^(a[144] & b[10])^(a[143] & b[11])^(a[142] & b[12])^(a[141] & b[13])^(a[140] & b[14])^(a[139] & b[15])^(a[138] & b[16])^(a[137] & b[17])^(a[136] & b[18])^(a[135] & b[19])^(a[134] & b[20])^(a[133] & b[21])^(a[132] & b[22])^(a[131] & b[23])^(a[130] & b[24])^(a[129] & b[25])^(a[128] & b[26])^(a[127] & b[27])^(a[126] & b[28])^(a[125] & b[29])^(a[124] & b[30])^(a[123] & b[31])^(a[122] & b[32])^(a[121] & b[33])^(a[120] & b[34])^(a[119] & b[35])^(a[118] & b[36])^(a[117] & b[37])^(a[116] & b[38])^(a[115] & b[39])^(a[114] & b[40])^(a[113] & b[41])^(a[112] & b[42])^(a[111] & b[43])^(a[110] & b[44])^(a[109] & b[45])^(a[108] & b[46])^(a[107] & b[47])^(a[106] & b[48])^(a[105] & b[49])^(a[104] & b[50])^(a[103] & b[51])^(a[102] & b[52])^(a[101] & b[53])^(a[100] & b[54])^(a[99] & b[55])^(a[98] & b[56])^(a[97] & b[57])^(a[96] & b[58])^(a[95] & b[59])^(a[94] & b[60])^(a[93] & b[61])^(a[92] & b[62])^(a[91] & b[63])^(a[90] & b[64])^(a[89] & b[65])^(a[88] & b[66])^(a[87] & b[67])^(a[86] & b[68])^(a[85] & b[69])^(a[84] & b[70])^(a[83] & b[71])^(a[82] & b[72])^(a[81] & b[73])^(a[80] & b[74])^(a[79] & b[75])^(a[78] & b[76])^(a[77] & b[77])^(a[76] & b[78])^(a[75] & b[79])^(a[74] & b[80])^(a[73] & b[81])^(a[72] & b[82])^(a[71] & b[83])^(a[70] & b[84])^(a[69] & b[85])^(a[68] & b[86])^(a[67] & b[87])^(a[66] & b[88])^(a[65] & b[89])^(a[64] & b[90])^(a[63] & b[91])^(a[62] & b[92])^(a[61] & b[93])^(a[60] & b[94])^(a[59] & b[95])^(a[58] & b[96])^(a[57] & b[97])^(a[56] & b[98])^(a[55] & b[99])^(a[54] & b[100])^(a[53] & b[101])^(a[52] & b[102])^(a[51] & b[103])^(a[50] & b[104])^(a[49] & b[105])^(a[48] & b[106])^(a[47] & b[107])^(a[46] & b[108])^(a[45] & b[109])^(a[44] & b[110])^(a[43] & b[111])^(a[42] & b[112])^(a[41] & b[113])^(a[40] & b[114])^(a[39] & b[115])^(a[38] & b[116])^(a[37] & b[117])^(a[36] & b[118])^(a[35] & b[119])^(a[34] & b[120])^(a[33] & b[121])^(a[32] & b[122])^(a[31] & b[123])^(a[30] & b[124])^(a[29] & b[125])^(a[28] & b[126])^(a[27] & b[127])^(a[26] & b[128])^(a[25] & b[129])^(a[24] & b[130])^(a[23] & b[131])^(a[22] & b[132])^(a[21] & b[133])^(a[20] & b[134])^(a[19] & b[135])^(a[18] & b[136])^(a[17] & b[137])^(a[16] & b[138])^(a[15] & b[139])^(a[14] & b[140])^(a[13] & b[141])^(a[12] & b[142])^(a[11] & b[143])^(a[10] & b[144])^(a[9] & b[145])^(a[8] & b[146])^(a[7] & b[147])^(a[6] & b[148])^(a[5] & b[149])^(a[4] & b[150])^(a[3] & b[151])^(a[2] & b[152])^(a[1] & b[153])^(a[0] & b[154]);
assign y[155] = (a[155] & b[0])^(a[154] & b[1])^(a[153] & b[2])^(a[152] & b[3])^(a[151] & b[4])^(a[150] & b[5])^(a[149] & b[6])^(a[148] & b[7])^(a[147] & b[8])^(a[146] & b[9])^(a[145] & b[10])^(a[144] & b[11])^(a[143] & b[12])^(a[142] & b[13])^(a[141] & b[14])^(a[140] & b[15])^(a[139] & b[16])^(a[138] & b[17])^(a[137] & b[18])^(a[136] & b[19])^(a[135] & b[20])^(a[134] & b[21])^(a[133] & b[22])^(a[132] & b[23])^(a[131] & b[24])^(a[130] & b[25])^(a[129] & b[26])^(a[128] & b[27])^(a[127] & b[28])^(a[126] & b[29])^(a[125] & b[30])^(a[124] & b[31])^(a[123] & b[32])^(a[122] & b[33])^(a[121] & b[34])^(a[120] & b[35])^(a[119] & b[36])^(a[118] & b[37])^(a[117] & b[38])^(a[116] & b[39])^(a[115] & b[40])^(a[114] & b[41])^(a[113] & b[42])^(a[112] & b[43])^(a[111] & b[44])^(a[110] & b[45])^(a[109] & b[46])^(a[108] & b[47])^(a[107] & b[48])^(a[106] & b[49])^(a[105] & b[50])^(a[104] & b[51])^(a[103] & b[52])^(a[102] & b[53])^(a[101] & b[54])^(a[100] & b[55])^(a[99] & b[56])^(a[98] & b[57])^(a[97] & b[58])^(a[96] & b[59])^(a[95] & b[60])^(a[94] & b[61])^(a[93] & b[62])^(a[92] & b[63])^(a[91] & b[64])^(a[90] & b[65])^(a[89] & b[66])^(a[88] & b[67])^(a[87] & b[68])^(a[86] & b[69])^(a[85] & b[70])^(a[84] & b[71])^(a[83] & b[72])^(a[82] & b[73])^(a[81] & b[74])^(a[80] & b[75])^(a[79] & b[76])^(a[78] & b[77])^(a[77] & b[78])^(a[76] & b[79])^(a[75] & b[80])^(a[74] & b[81])^(a[73] & b[82])^(a[72] & b[83])^(a[71] & b[84])^(a[70] & b[85])^(a[69] & b[86])^(a[68] & b[87])^(a[67] & b[88])^(a[66] & b[89])^(a[65] & b[90])^(a[64] & b[91])^(a[63] & b[92])^(a[62] & b[93])^(a[61] & b[94])^(a[60] & b[95])^(a[59] & b[96])^(a[58] & b[97])^(a[57] & b[98])^(a[56] & b[99])^(a[55] & b[100])^(a[54] & b[101])^(a[53] & b[102])^(a[52] & b[103])^(a[51] & b[104])^(a[50] & b[105])^(a[49] & b[106])^(a[48] & b[107])^(a[47] & b[108])^(a[46] & b[109])^(a[45] & b[110])^(a[44] & b[111])^(a[43] & b[112])^(a[42] & b[113])^(a[41] & b[114])^(a[40] & b[115])^(a[39] & b[116])^(a[38] & b[117])^(a[37] & b[118])^(a[36] & b[119])^(a[35] & b[120])^(a[34] & b[121])^(a[33] & b[122])^(a[32] & b[123])^(a[31] & b[124])^(a[30] & b[125])^(a[29] & b[126])^(a[28] & b[127])^(a[27] & b[128])^(a[26] & b[129])^(a[25] & b[130])^(a[24] & b[131])^(a[23] & b[132])^(a[22] & b[133])^(a[21] & b[134])^(a[20] & b[135])^(a[19] & b[136])^(a[18] & b[137])^(a[17] & b[138])^(a[16] & b[139])^(a[15] & b[140])^(a[14] & b[141])^(a[13] & b[142])^(a[12] & b[143])^(a[11] & b[144])^(a[10] & b[145])^(a[9] & b[146])^(a[8] & b[147])^(a[7] & b[148])^(a[6] & b[149])^(a[5] & b[150])^(a[4] & b[151])^(a[3] & b[152])^(a[2] & b[153])^(a[1] & b[154])^(a[0] & b[155]);
assign y[156] = (a[156] & b[0])^(a[155] & b[1])^(a[154] & b[2])^(a[153] & b[3])^(a[152] & b[4])^(a[151] & b[5])^(a[150] & b[6])^(a[149] & b[7])^(a[148] & b[8])^(a[147] & b[9])^(a[146] & b[10])^(a[145] & b[11])^(a[144] & b[12])^(a[143] & b[13])^(a[142] & b[14])^(a[141] & b[15])^(a[140] & b[16])^(a[139] & b[17])^(a[138] & b[18])^(a[137] & b[19])^(a[136] & b[20])^(a[135] & b[21])^(a[134] & b[22])^(a[133] & b[23])^(a[132] & b[24])^(a[131] & b[25])^(a[130] & b[26])^(a[129] & b[27])^(a[128] & b[28])^(a[127] & b[29])^(a[126] & b[30])^(a[125] & b[31])^(a[124] & b[32])^(a[123] & b[33])^(a[122] & b[34])^(a[121] & b[35])^(a[120] & b[36])^(a[119] & b[37])^(a[118] & b[38])^(a[117] & b[39])^(a[116] & b[40])^(a[115] & b[41])^(a[114] & b[42])^(a[113] & b[43])^(a[112] & b[44])^(a[111] & b[45])^(a[110] & b[46])^(a[109] & b[47])^(a[108] & b[48])^(a[107] & b[49])^(a[106] & b[50])^(a[105] & b[51])^(a[104] & b[52])^(a[103] & b[53])^(a[102] & b[54])^(a[101] & b[55])^(a[100] & b[56])^(a[99] & b[57])^(a[98] & b[58])^(a[97] & b[59])^(a[96] & b[60])^(a[95] & b[61])^(a[94] & b[62])^(a[93] & b[63])^(a[92] & b[64])^(a[91] & b[65])^(a[90] & b[66])^(a[89] & b[67])^(a[88] & b[68])^(a[87] & b[69])^(a[86] & b[70])^(a[85] & b[71])^(a[84] & b[72])^(a[83] & b[73])^(a[82] & b[74])^(a[81] & b[75])^(a[80] & b[76])^(a[79] & b[77])^(a[78] & b[78])^(a[77] & b[79])^(a[76] & b[80])^(a[75] & b[81])^(a[74] & b[82])^(a[73] & b[83])^(a[72] & b[84])^(a[71] & b[85])^(a[70] & b[86])^(a[69] & b[87])^(a[68] & b[88])^(a[67] & b[89])^(a[66] & b[90])^(a[65] & b[91])^(a[64] & b[92])^(a[63] & b[93])^(a[62] & b[94])^(a[61] & b[95])^(a[60] & b[96])^(a[59] & b[97])^(a[58] & b[98])^(a[57] & b[99])^(a[56] & b[100])^(a[55] & b[101])^(a[54] & b[102])^(a[53] & b[103])^(a[52] & b[104])^(a[51] & b[105])^(a[50] & b[106])^(a[49] & b[107])^(a[48] & b[108])^(a[47] & b[109])^(a[46] & b[110])^(a[45] & b[111])^(a[44] & b[112])^(a[43] & b[113])^(a[42] & b[114])^(a[41] & b[115])^(a[40] & b[116])^(a[39] & b[117])^(a[38] & b[118])^(a[37] & b[119])^(a[36] & b[120])^(a[35] & b[121])^(a[34] & b[122])^(a[33] & b[123])^(a[32] & b[124])^(a[31] & b[125])^(a[30] & b[126])^(a[29] & b[127])^(a[28] & b[128])^(a[27] & b[129])^(a[26] & b[130])^(a[25] & b[131])^(a[24] & b[132])^(a[23] & b[133])^(a[22] & b[134])^(a[21] & b[135])^(a[20] & b[136])^(a[19] & b[137])^(a[18] & b[138])^(a[17] & b[139])^(a[16] & b[140])^(a[15] & b[141])^(a[14] & b[142])^(a[13] & b[143])^(a[12] & b[144])^(a[11] & b[145])^(a[10] & b[146])^(a[9] & b[147])^(a[8] & b[148])^(a[7] & b[149])^(a[6] & b[150])^(a[5] & b[151])^(a[4] & b[152])^(a[3] & b[153])^(a[2] & b[154])^(a[1] & b[155])^(a[0] & b[156]);
assign y[157] = (a[157] & b[0])^(a[156] & b[1])^(a[155] & b[2])^(a[154] & b[3])^(a[153] & b[4])^(a[152] & b[5])^(a[151] & b[6])^(a[150] & b[7])^(a[149] & b[8])^(a[148] & b[9])^(a[147] & b[10])^(a[146] & b[11])^(a[145] & b[12])^(a[144] & b[13])^(a[143] & b[14])^(a[142] & b[15])^(a[141] & b[16])^(a[140] & b[17])^(a[139] & b[18])^(a[138] & b[19])^(a[137] & b[20])^(a[136] & b[21])^(a[135] & b[22])^(a[134] & b[23])^(a[133] & b[24])^(a[132] & b[25])^(a[131] & b[26])^(a[130] & b[27])^(a[129] & b[28])^(a[128] & b[29])^(a[127] & b[30])^(a[126] & b[31])^(a[125] & b[32])^(a[124] & b[33])^(a[123] & b[34])^(a[122] & b[35])^(a[121] & b[36])^(a[120] & b[37])^(a[119] & b[38])^(a[118] & b[39])^(a[117] & b[40])^(a[116] & b[41])^(a[115] & b[42])^(a[114] & b[43])^(a[113] & b[44])^(a[112] & b[45])^(a[111] & b[46])^(a[110] & b[47])^(a[109] & b[48])^(a[108] & b[49])^(a[107] & b[50])^(a[106] & b[51])^(a[105] & b[52])^(a[104] & b[53])^(a[103] & b[54])^(a[102] & b[55])^(a[101] & b[56])^(a[100] & b[57])^(a[99] & b[58])^(a[98] & b[59])^(a[97] & b[60])^(a[96] & b[61])^(a[95] & b[62])^(a[94] & b[63])^(a[93] & b[64])^(a[92] & b[65])^(a[91] & b[66])^(a[90] & b[67])^(a[89] & b[68])^(a[88] & b[69])^(a[87] & b[70])^(a[86] & b[71])^(a[85] & b[72])^(a[84] & b[73])^(a[83] & b[74])^(a[82] & b[75])^(a[81] & b[76])^(a[80] & b[77])^(a[79] & b[78])^(a[78] & b[79])^(a[77] & b[80])^(a[76] & b[81])^(a[75] & b[82])^(a[74] & b[83])^(a[73] & b[84])^(a[72] & b[85])^(a[71] & b[86])^(a[70] & b[87])^(a[69] & b[88])^(a[68] & b[89])^(a[67] & b[90])^(a[66] & b[91])^(a[65] & b[92])^(a[64] & b[93])^(a[63] & b[94])^(a[62] & b[95])^(a[61] & b[96])^(a[60] & b[97])^(a[59] & b[98])^(a[58] & b[99])^(a[57] & b[100])^(a[56] & b[101])^(a[55] & b[102])^(a[54] & b[103])^(a[53] & b[104])^(a[52] & b[105])^(a[51] & b[106])^(a[50] & b[107])^(a[49] & b[108])^(a[48] & b[109])^(a[47] & b[110])^(a[46] & b[111])^(a[45] & b[112])^(a[44] & b[113])^(a[43] & b[114])^(a[42] & b[115])^(a[41] & b[116])^(a[40] & b[117])^(a[39] & b[118])^(a[38] & b[119])^(a[37] & b[120])^(a[36] & b[121])^(a[35] & b[122])^(a[34] & b[123])^(a[33] & b[124])^(a[32] & b[125])^(a[31] & b[126])^(a[30] & b[127])^(a[29] & b[128])^(a[28] & b[129])^(a[27] & b[130])^(a[26] & b[131])^(a[25] & b[132])^(a[24] & b[133])^(a[23] & b[134])^(a[22] & b[135])^(a[21] & b[136])^(a[20] & b[137])^(a[19] & b[138])^(a[18] & b[139])^(a[17] & b[140])^(a[16] & b[141])^(a[15] & b[142])^(a[14] & b[143])^(a[13] & b[144])^(a[12] & b[145])^(a[11] & b[146])^(a[10] & b[147])^(a[9] & b[148])^(a[8] & b[149])^(a[7] & b[150])^(a[6] & b[151])^(a[5] & b[152])^(a[4] & b[153])^(a[3] & b[154])^(a[2] & b[155])^(a[1] & b[156])^(a[0] & b[157]);
assign y[158] = (a[158] & b[0])^(a[157] & b[1])^(a[156] & b[2])^(a[155] & b[3])^(a[154] & b[4])^(a[153] & b[5])^(a[152] & b[6])^(a[151] & b[7])^(a[150] & b[8])^(a[149] & b[9])^(a[148] & b[10])^(a[147] & b[11])^(a[146] & b[12])^(a[145] & b[13])^(a[144] & b[14])^(a[143] & b[15])^(a[142] & b[16])^(a[141] & b[17])^(a[140] & b[18])^(a[139] & b[19])^(a[138] & b[20])^(a[137] & b[21])^(a[136] & b[22])^(a[135] & b[23])^(a[134] & b[24])^(a[133] & b[25])^(a[132] & b[26])^(a[131] & b[27])^(a[130] & b[28])^(a[129] & b[29])^(a[128] & b[30])^(a[127] & b[31])^(a[126] & b[32])^(a[125] & b[33])^(a[124] & b[34])^(a[123] & b[35])^(a[122] & b[36])^(a[121] & b[37])^(a[120] & b[38])^(a[119] & b[39])^(a[118] & b[40])^(a[117] & b[41])^(a[116] & b[42])^(a[115] & b[43])^(a[114] & b[44])^(a[113] & b[45])^(a[112] & b[46])^(a[111] & b[47])^(a[110] & b[48])^(a[109] & b[49])^(a[108] & b[50])^(a[107] & b[51])^(a[106] & b[52])^(a[105] & b[53])^(a[104] & b[54])^(a[103] & b[55])^(a[102] & b[56])^(a[101] & b[57])^(a[100] & b[58])^(a[99] & b[59])^(a[98] & b[60])^(a[97] & b[61])^(a[96] & b[62])^(a[95] & b[63])^(a[94] & b[64])^(a[93] & b[65])^(a[92] & b[66])^(a[91] & b[67])^(a[90] & b[68])^(a[89] & b[69])^(a[88] & b[70])^(a[87] & b[71])^(a[86] & b[72])^(a[85] & b[73])^(a[84] & b[74])^(a[83] & b[75])^(a[82] & b[76])^(a[81] & b[77])^(a[80] & b[78])^(a[79] & b[79])^(a[78] & b[80])^(a[77] & b[81])^(a[76] & b[82])^(a[75] & b[83])^(a[74] & b[84])^(a[73] & b[85])^(a[72] & b[86])^(a[71] & b[87])^(a[70] & b[88])^(a[69] & b[89])^(a[68] & b[90])^(a[67] & b[91])^(a[66] & b[92])^(a[65] & b[93])^(a[64] & b[94])^(a[63] & b[95])^(a[62] & b[96])^(a[61] & b[97])^(a[60] & b[98])^(a[59] & b[99])^(a[58] & b[100])^(a[57] & b[101])^(a[56] & b[102])^(a[55] & b[103])^(a[54] & b[104])^(a[53] & b[105])^(a[52] & b[106])^(a[51] & b[107])^(a[50] & b[108])^(a[49] & b[109])^(a[48] & b[110])^(a[47] & b[111])^(a[46] & b[112])^(a[45] & b[113])^(a[44] & b[114])^(a[43] & b[115])^(a[42] & b[116])^(a[41] & b[117])^(a[40] & b[118])^(a[39] & b[119])^(a[38] & b[120])^(a[37] & b[121])^(a[36] & b[122])^(a[35] & b[123])^(a[34] & b[124])^(a[33] & b[125])^(a[32] & b[126])^(a[31] & b[127])^(a[30] & b[128])^(a[29] & b[129])^(a[28] & b[130])^(a[27] & b[131])^(a[26] & b[132])^(a[25] & b[133])^(a[24] & b[134])^(a[23] & b[135])^(a[22] & b[136])^(a[21] & b[137])^(a[20] & b[138])^(a[19] & b[139])^(a[18] & b[140])^(a[17] & b[141])^(a[16] & b[142])^(a[15] & b[143])^(a[14] & b[144])^(a[13] & b[145])^(a[12] & b[146])^(a[11] & b[147])^(a[10] & b[148])^(a[9] & b[149])^(a[8] & b[150])^(a[7] & b[151])^(a[6] & b[152])^(a[5] & b[153])^(a[4] & b[154])^(a[3] & b[155])^(a[2] & b[156])^(a[1] & b[157])^(a[0] & b[158]);
assign y[159] = (a[159] & b[0])^(a[158] & b[1])^(a[157] & b[2])^(a[156] & b[3])^(a[155] & b[4])^(a[154] & b[5])^(a[153] & b[6])^(a[152] & b[7])^(a[151] & b[8])^(a[150] & b[9])^(a[149] & b[10])^(a[148] & b[11])^(a[147] & b[12])^(a[146] & b[13])^(a[145] & b[14])^(a[144] & b[15])^(a[143] & b[16])^(a[142] & b[17])^(a[141] & b[18])^(a[140] & b[19])^(a[139] & b[20])^(a[138] & b[21])^(a[137] & b[22])^(a[136] & b[23])^(a[135] & b[24])^(a[134] & b[25])^(a[133] & b[26])^(a[132] & b[27])^(a[131] & b[28])^(a[130] & b[29])^(a[129] & b[30])^(a[128] & b[31])^(a[127] & b[32])^(a[126] & b[33])^(a[125] & b[34])^(a[124] & b[35])^(a[123] & b[36])^(a[122] & b[37])^(a[121] & b[38])^(a[120] & b[39])^(a[119] & b[40])^(a[118] & b[41])^(a[117] & b[42])^(a[116] & b[43])^(a[115] & b[44])^(a[114] & b[45])^(a[113] & b[46])^(a[112] & b[47])^(a[111] & b[48])^(a[110] & b[49])^(a[109] & b[50])^(a[108] & b[51])^(a[107] & b[52])^(a[106] & b[53])^(a[105] & b[54])^(a[104] & b[55])^(a[103] & b[56])^(a[102] & b[57])^(a[101] & b[58])^(a[100] & b[59])^(a[99] & b[60])^(a[98] & b[61])^(a[97] & b[62])^(a[96] & b[63])^(a[95] & b[64])^(a[94] & b[65])^(a[93] & b[66])^(a[92] & b[67])^(a[91] & b[68])^(a[90] & b[69])^(a[89] & b[70])^(a[88] & b[71])^(a[87] & b[72])^(a[86] & b[73])^(a[85] & b[74])^(a[84] & b[75])^(a[83] & b[76])^(a[82] & b[77])^(a[81] & b[78])^(a[80] & b[79])^(a[79] & b[80])^(a[78] & b[81])^(a[77] & b[82])^(a[76] & b[83])^(a[75] & b[84])^(a[74] & b[85])^(a[73] & b[86])^(a[72] & b[87])^(a[71] & b[88])^(a[70] & b[89])^(a[69] & b[90])^(a[68] & b[91])^(a[67] & b[92])^(a[66] & b[93])^(a[65] & b[94])^(a[64] & b[95])^(a[63] & b[96])^(a[62] & b[97])^(a[61] & b[98])^(a[60] & b[99])^(a[59] & b[100])^(a[58] & b[101])^(a[57] & b[102])^(a[56] & b[103])^(a[55] & b[104])^(a[54] & b[105])^(a[53] & b[106])^(a[52] & b[107])^(a[51] & b[108])^(a[50] & b[109])^(a[49] & b[110])^(a[48] & b[111])^(a[47] & b[112])^(a[46] & b[113])^(a[45] & b[114])^(a[44] & b[115])^(a[43] & b[116])^(a[42] & b[117])^(a[41] & b[118])^(a[40] & b[119])^(a[39] & b[120])^(a[38] & b[121])^(a[37] & b[122])^(a[36] & b[123])^(a[35] & b[124])^(a[34] & b[125])^(a[33] & b[126])^(a[32] & b[127])^(a[31] & b[128])^(a[30] & b[129])^(a[29] & b[130])^(a[28] & b[131])^(a[27] & b[132])^(a[26] & b[133])^(a[25] & b[134])^(a[24] & b[135])^(a[23] & b[136])^(a[22] & b[137])^(a[21] & b[138])^(a[20] & b[139])^(a[19] & b[140])^(a[18] & b[141])^(a[17] & b[142])^(a[16] & b[143])^(a[15] & b[144])^(a[14] & b[145])^(a[13] & b[146])^(a[12] & b[147])^(a[11] & b[148])^(a[10] & b[149])^(a[9] & b[150])^(a[8] & b[151])^(a[7] & b[152])^(a[6] & b[153])^(a[5] & b[154])^(a[4] & b[155])^(a[3] & b[156])^(a[2] & b[157])^(a[1] & b[158])^(a[0] & b[159]);
assign y[160] = (a[160] & b[0])^(a[159] & b[1])^(a[158] & b[2])^(a[157] & b[3])^(a[156] & b[4])^(a[155] & b[5])^(a[154] & b[6])^(a[153] & b[7])^(a[152] & b[8])^(a[151] & b[9])^(a[150] & b[10])^(a[149] & b[11])^(a[148] & b[12])^(a[147] & b[13])^(a[146] & b[14])^(a[145] & b[15])^(a[144] & b[16])^(a[143] & b[17])^(a[142] & b[18])^(a[141] & b[19])^(a[140] & b[20])^(a[139] & b[21])^(a[138] & b[22])^(a[137] & b[23])^(a[136] & b[24])^(a[135] & b[25])^(a[134] & b[26])^(a[133] & b[27])^(a[132] & b[28])^(a[131] & b[29])^(a[130] & b[30])^(a[129] & b[31])^(a[128] & b[32])^(a[127] & b[33])^(a[126] & b[34])^(a[125] & b[35])^(a[124] & b[36])^(a[123] & b[37])^(a[122] & b[38])^(a[121] & b[39])^(a[120] & b[40])^(a[119] & b[41])^(a[118] & b[42])^(a[117] & b[43])^(a[116] & b[44])^(a[115] & b[45])^(a[114] & b[46])^(a[113] & b[47])^(a[112] & b[48])^(a[111] & b[49])^(a[110] & b[50])^(a[109] & b[51])^(a[108] & b[52])^(a[107] & b[53])^(a[106] & b[54])^(a[105] & b[55])^(a[104] & b[56])^(a[103] & b[57])^(a[102] & b[58])^(a[101] & b[59])^(a[100] & b[60])^(a[99] & b[61])^(a[98] & b[62])^(a[97] & b[63])^(a[96] & b[64])^(a[95] & b[65])^(a[94] & b[66])^(a[93] & b[67])^(a[92] & b[68])^(a[91] & b[69])^(a[90] & b[70])^(a[89] & b[71])^(a[88] & b[72])^(a[87] & b[73])^(a[86] & b[74])^(a[85] & b[75])^(a[84] & b[76])^(a[83] & b[77])^(a[82] & b[78])^(a[81] & b[79])^(a[80] & b[80])^(a[79] & b[81])^(a[78] & b[82])^(a[77] & b[83])^(a[76] & b[84])^(a[75] & b[85])^(a[74] & b[86])^(a[73] & b[87])^(a[72] & b[88])^(a[71] & b[89])^(a[70] & b[90])^(a[69] & b[91])^(a[68] & b[92])^(a[67] & b[93])^(a[66] & b[94])^(a[65] & b[95])^(a[64] & b[96])^(a[63] & b[97])^(a[62] & b[98])^(a[61] & b[99])^(a[60] & b[100])^(a[59] & b[101])^(a[58] & b[102])^(a[57] & b[103])^(a[56] & b[104])^(a[55] & b[105])^(a[54] & b[106])^(a[53] & b[107])^(a[52] & b[108])^(a[51] & b[109])^(a[50] & b[110])^(a[49] & b[111])^(a[48] & b[112])^(a[47] & b[113])^(a[46] & b[114])^(a[45] & b[115])^(a[44] & b[116])^(a[43] & b[117])^(a[42] & b[118])^(a[41] & b[119])^(a[40] & b[120])^(a[39] & b[121])^(a[38] & b[122])^(a[37] & b[123])^(a[36] & b[124])^(a[35] & b[125])^(a[34] & b[126])^(a[33] & b[127])^(a[32] & b[128])^(a[31] & b[129])^(a[30] & b[130])^(a[29] & b[131])^(a[28] & b[132])^(a[27] & b[133])^(a[26] & b[134])^(a[25] & b[135])^(a[24] & b[136])^(a[23] & b[137])^(a[22] & b[138])^(a[21] & b[139])^(a[20] & b[140])^(a[19] & b[141])^(a[18] & b[142])^(a[17] & b[143])^(a[16] & b[144])^(a[15] & b[145])^(a[14] & b[146])^(a[13] & b[147])^(a[12] & b[148])^(a[11] & b[149])^(a[10] & b[150])^(a[9] & b[151])^(a[8] & b[152])^(a[7] & b[153])^(a[6] & b[154])^(a[5] & b[155])^(a[4] & b[156])^(a[3] & b[157])^(a[2] & b[158])^(a[1] & b[159])^(a[0] & b[160]);
assign y[161] = (a[161] & b[0])^(a[160] & b[1])^(a[159] & b[2])^(a[158] & b[3])^(a[157] & b[4])^(a[156] & b[5])^(a[155] & b[6])^(a[154] & b[7])^(a[153] & b[8])^(a[152] & b[9])^(a[151] & b[10])^(a[150] & b[11])^(a[149] & b[12])^(a[148] & b[13])^(a[147] & b[14])^(a[146] & b[15])^(a[145] & b[16])^(a[144] & b[17])^(a[143] & b[18])^(a[142] & b[19])^(a[141] & b[20])^(a[140] & b[21])^(a[139] & b[22])^(a[138] & b[23])^(a[137] & b[24])^(a[136] & b[25])^(a[135] & b[26])^(a[134] & b[27])^(a[133] & b[28])^(a[132] & b[29])^(a[131] & b[30])^(a[130] & b[31])^(a[129] & b[32])^(a[128] & b[33])^(a[127] & b[34])^(a[126] & b[35])^(a[125] & b[36])^(a[124] & b[37])^(a[123] & b[38])^(a[122] & b[39])^(a[121] & b[40])^(a[120] & b[41])^(a[119] & b[42])^(a[118] & b[43])^(a[117] & b[44])^(a[116] & b[45])^(a[115] & b[46])^(a[114] & b[47])^(a[113] & b[48])^(a[112] & b[49])^(a[111] & b[50])^(a[110] & b[51])^(a[109] & b[52])^(a[108] & b[53])^(a[107] & b[54])^(a[106] & b[55])^(a[105] & b[56])^(a[104] & b[57])^(a[103] & b[58])^(a[102] & b[59])^(a[101] & b[60])^(a[100] & b[61])^(a[99] & b[62])^(a[98] & b[63])^(a[97] & b[64])^(a[96] & b[65])^(a[95] & b[66])^(a[94] & b[67])^(a[93] & b[68])^(a[92] & b[69])^(a[91] & b[70])^(a[90] & b[71])^(a[89] & b[72])^(a[88] & b[73])^(a[87] & b[74])^(a[86] & b[75])^(a[85] & b[76])^(a[84] & b[77])^(a[83] & b[78])^(a[82] & b[79])^(a[81] & b[80])^(a[80] & b[81])^(a[79] & b[82])^(a[78] & b[83])^(a[77] & b[84])^(a[76] & b[85])^(a[75] & b[86])^(a[74] & b[87])^(a[73] & b[88])^(a[72] & b[89])^(a[71] & b[90])^(a[70] & b[91])^(a[69] & b[92])^(a[68] & b[93])^(a[67] & b[94])^(a[66] & b[95])^(a[65] & b[96])^(a[64] & b[97])^(a[63] & b[98])^(a[62] & b[99])^(a[61] & b[100])^(a[60] & b[101])^(a[59] & b[102])^(a[58] & b[103])^(a[57] & b[104])^(a[56] & b[105])^(a[55] & b[106])^(a[54] & b[107])^(a[53] & b[108])^(a[52] & b[109])^(a[51] & b[110])^(a[50] & b[111])^(a[49] & b[112])^(a[48] & b[113])^(a[47] & b[114])^(a[46] & b[115])^(a[45] & b[116])^(a[44] & b[117])^(a[43] & b[118])^(a[42] & b[119])^(a[41] & b[120])^(a[40] & b[121])^(a[39] & b[122])^(a[38] & b[123])^(a[37] & b[124])^(a[36] & b[125])^(a[35] & b[126])^(a[34] & b[127])^(a[33] & b[128])^(a[32] & b[129])^(a[31] & b[130])^(a[30] & b[131])^(a[29] & b[132])^(a[28] & b[133])^(a[27] & b[134])^(a[26] & b[135])^(a[25] & b[136])^(a[24] & b[137])^(a[23] & b[138])^(a[22] & b[139])^(a[21] & b[140])^(a[20] & b[141])^(a[19] & b[142])^(a[18] & b[143])^(a[17] & b[144])^(a[16] & b[145])^(a[15] & b[146])^(a[14] & b[147])^(a[13] & b[148])^(a[12] & b[149])^(a[11] & b[150])^(a[10] & b[151])^(a[9] & b[152])^(a[8] & b[153])^(a[7] & b[154])^(a[6] & b[155])^(a[5] & b[156])^(a[4] & b[157])^(a[3] & b[158])^(a[2] & b[159])^(a[1] & b[160])^(a[0] & b[161]);
assign y[162] = (a[162] & b[0])^(a[161] & b[1])^(a[160] & b[2])^(a[159] & b[3])^(a[158] & b[4])^(a[157] & b[5])^(a[156] & b[6])^(a[155] & b[7])^(a[154] & b[8])^(a[153] & b[9])^(a[152] & b[10])^(a[151] & b[11])^(a[150] & b[12])^(a[149] & b[13])^(a[148] & b[14])^(a[147] & b[15])^(a[146] & b[16])^(a[145] & b[17])^(a[144] & b[18])^(a[143] & b[19])^(a[142] & b[20])^(a[141] & b[21])^(a[140] & b[22])^(a[139] & b[23])^(a[138] & b[24])^(a[137] & b[25])^(a[136] & b[26])^(a[135] & b[27])^(a[134] & b[28])^(a[133] & b[29])^(a[132] & b[30])^(a[131] & b[31])^(a[130] & b[32])^(a[129] & b[33])^(a[128] & b[34])^(a[127] & b[35])^(a[126] & b[36])^(a[125] & b[37])^(a[124] & b[38])^(a[123] & b[39])^(a[122] & b[40])^(a[121] & b[41])^(a[120] & b[42])^(a[119] & b[43])^(a[118] & b[44])^(a[117] & b[45])^(a[116] & b[46])^(a[115] & b[47])^(a[114] & b[48])^(a[113] & b[49])^(a[112] & b[50])^(a[111] & b[51])^(a[110] & b[52])^(a[109] & b[53])^(a[108] & b[54])^(a[107] & b[55])^(a[106] & b[56])^(a[105] & b[57])^(a[104] & b[58])^(a[103] & b[59])^(a[102] & b[60])^(a[101] & b[61])^(a[100] & b[62])^(a[99] & b[63])^(a[98] & b[64])^(a[97] & b[65])^(a[96] & b[66])^(a[95] & b[67])^(a[94] & b[68])^(a[93] & b[69])^(a[92] & b[70])^(a[91] & b[71])^(a[90] & b[72])^(a[89] & b[73])^(a[88] & b[74])^(a[87] & b[75])^(a[86] & b[76])^(a[85] & b[77])^(a[84] & b[78])^(a[83] & b[79])^(a[82] & b[80])^(a[81] & b[81])^(a[80] & b[82])^(a[79] & b[83])^(a[78] & b[84])^(a[77] & b[85])^(a[76] & b[86])^(a[75] & b[87])^(a[74] & b[88])^(a[73] & b[89])^(a[72] & b[90])^(a[71] & b[91])^(a[70] & b[92])^(a[69] & b[93])^(a[68] & b[94])^(a[67] & b[95])^(a[66] & b[96])^(a[65] & b[97])^(a[64] & b[98])^(a[63] & b[99])^(a[62] & b[100])^(a[61] & b[101])^(a[60] & b[102])^(a[59] & b[103])^(a[58] & b[104])^(a[57] & b[105])^(a[56] & b[106])^(a[55] & b[107])^(a[54] & b[108])^(a[53] & b[109])^(a[52] & b[110])^(a[51] & b[111])^(a[50] & b[112])^(a[49] & b[113])^(a[48] & b[114])^(a[47] & b[115])^(a[46] & b[116])^(a[45] & b[117])^(a[44] & b[118])^(a[43] & b[119])^(a[42] & b[120])^(a[41] & b[121])^(a[40] & b[122])^(a[39] & b[123])^(a[38] & b[124])^(a[37] & b[125])^(a[36] & b[126])^(a[35] & b[127])^(a[34] & b[128])^(a[33] & b[129])^(a[32] & b[130])^(a[31] & b[131])^(a[30] & b[132])^(a[29] & b[133])^(a[28] & b[134])^(a[27] & b[135])^(a[26] & b[136])^(a[25] & b[137])^(a[24] & b[138])^(a[23] & b[139])^(a[22] & b[140])^(a[21] & b[141])^(a[20] & b[142])^(a[19] & b[143])^(a[18] & b[144])^(a[17] & b[145])^(a[16] & b[146])^(a[15] & b[147])^(a[14] & b[148])^(a[13] & b[149])^(a[12] & b[150])^(a[11] & b[151])^(a[10] & b[152])^(a[9] & b[153])^(a[8] & b[154])^(a[7] & b[155])^(a[6] & b[156])^(a[5] & b[157])^(a[4] & b[158])^(a[3] & b[159])^(a[2] & b[160])^(a[1] & b[161])^(a[0] & b[162]);
assign y[163] = (a[162] & b[1])^(a[161] & b[2])^(a[160] & b[3])^(a[159] & b[4])^(a[158] & b[5])^(a[157] & b[6])^(a[156] & b[7])^(a[155] & b[8])^(a[154] & b[9])^(a[153] & b[10])^(a[152] & b[11])^(a[151] & b[12])^(a[150] & b[13])^(a[149] & b[14])^(a[148] & b[15])^(a[147] & b[16])^(a[146] & b[17])^(a[145] & b[18])^(a[144] & b[19])^(a[143] & b[20])^(a[142] & b[21])^(a[141] & b[22])^(a[140] & b[23])^(a[139] & b[24])^(a[138] & b[25])^(a[137] & b[26])^(a[136] & b[27])^(a[135] & b[28])^(a[134] & b[29])^(a[133] & b[30])^(a[132] & b[31])^(a[131] & b[32])^(a[130] & b[33])^(a[129] & b[34])^(a[128] & b[35])^(a[127] & b[36])^(a[126] & b[37])^(a[125] & b[38])^(a[124] & b[39])^(a[123] & b[40])^(a[122] & b[41])^(a[121] & b[42])^(a[120] & b[43])^(a[119] & b[44])^(a[118] & b[45])^(a[117] & b[46])^(a[116] & b[47])^(a[115] & b[48])^(a[114] & b[49])^(a[113] & b[50])^(a[112] & b[51])^(a[111] & b[52])^(a[110] & b[53])^(a[109] & b[54])^(a[108] & b[55])^(a[107] & b[56])^(a[106] & b[57])^(a[105] & b[58])^(a[104] & b[59])^(a[103] & b[60])^(a[102] & b[61])^(a[101] & b[62])^(a[100] & b[63])^(a[99] & b[64])^(a[98] & b[65])^(a[97] & b[66])^(a[96] & b[67])^(a[95] & b[68])^(a[94] & b[69])^(a[93] & b[70])^(a[92] & b[71])^(a[91] & b[72])^(a[90] & b[73])^(a[89] & b[74])^(a[88] & b[75])^(a[87] & b[76])^(a[86] & b[77])^(a[85] & b[78])^(a[84] & b[79])^(a[83] & b[80])^(a[82] & b[81])^(a[81] & b[82])^(a[80] & b[83])^(a[79] & b[84])^(a[78] & b[85])^(a[77] & b[86])^(a[76] & b[87])^(a[75] & b[88])^(a[74] & b[89])^(a[73] & b[90])^(a[72] & b[91])^(a[71] & b[92])^(a[70] & b[93])^(a[69] & b[94])^(a[68] & b[95])^(a[67] & b[96])^(a[66] & b[97])^(a[65] & b[98])^(a[64] & b[99])^(a[63] & b[100])^(a[62] & b[101])^(a[61] & b[102])^(a[60] & b[103])^(a[59] & b[104])^(a[58] & b[105])^(a[57] & b[106])^(a[56] & b[107])^(a[55] & b[108])^(a[54] & b[109])^(a[53] & b[110])^(a[52] & b[111])^(a[51] & b[112])^(a[50] & b[113])^(a[49] & b[114])^(a[48] & b[115])^(a[47] & b[116])^(a[46] & b[117])^(a[45] & b[118])^(a[44] & b[119])^(a[43] & b[120])^(a[42] & b[121])^(a[41] & b[122])^(a[40] & b[123])^(a[39] & b[124])^(a[38] & b[125])^(a[37] & b[126])^(a[36] & b[127])^(a[35] & b[128])^(a[34] & b[129])^(a[33] & b[130])^(a[32] & b[131])^(a[31] & b[132])^(a[30] & b[133])^(a[29] & b[134])^(a[28] & b[135])^(a[27] & b[136])^(a[26] & b[137])^(a[25] & b[138])^(a[24] & b[139])^(a[23] & b[140])^(a[22] & b[141])^(a[21] & b[142])^(a[20] & b[143])^(a[19] & b[144])^(a[18] & b[145])^(a[17] & b[146])^(a[16] & b[147])^(a[15] & b[148])^(a[14] & b[149])^(a[13] & b[150])^(a[12] & b[151])^(a[11] & b[152])^(a[10] & b[153])^(a[9] & b[154])^(a[8] & b[155])^(a[7] & b[156])^(a[6] & b[157])^(a[5] & b[158])^(a[4] & b[159])^(a[3] & b[160])^(a[2] & b[161])^(a[1] & b[162]);
assign y[164] = (a[162] & b[2])^(a[161] & b[3])^(a[160] & b[4])^(a[159] & b[5])^(a[158] & b[6])^(a[157] & b[7])^(a[156] & b[8])^(a[155] & b[9])^(a[154] & b[10])^(a[153] & b[11])^(a[152] & b[12])^(a[151] & b[13])^(a[150] & b[14])^(a[149] & b[15])^(a[148] & b[16])^(a[147] & b[17])^(a[146] & b[18])^(a[145] & b[19])^(a[144] & b[20])^(a[143] & b[21])^(a[142] & b[22])^(a[141] & b[23])^(a[140] & b[24])^(a[139] & b[25])^(a[138] & b[26])^(a[137] & b[27])^(a[136] & b[28])^(a[135] & b[29])^(a[134] & b[30])^(a[133] & b[31])^(a[132] & b[32])^(a[131] & b[33])^(a[130] & b[34])^(a[129] & b[35])^(a[128] & b[36])^(a[127] & b[37])^(a[126] & b[38])^(a[125] & b[39])^(a[124] & b[40])^(a[123] & b[41])^(a[122] & b[42])^(a[121] & b[43])^(a[120] & b[44])^(a[119] & b[45])^(a[118] & b[46])^(a[117] & b[47])^(a[116] & b[48])^(a[115] & b[49])^(a[114] & b[50])^(a[113] & b[51])^(a[112] & b[52])^(a[111] & b[53])^(a[110] & b[54])^(a[109] & b[55])^(a[108] & b[56])^(a[107] & b[57])^(a[106] & b[58])^(a[105] & b[59])^(a[104] & b[60])^(a[103] & b[61])^(a[102] & b[62])^(a[101] & b[63])^(a[100] & b[64])^(a[99] & b[65])^(a[98] & b[66])^(a[97] & b[67])^(a[96] & b[68])^(a[95] & b[69])^(a[94] & b[70])^(a[93] & b[71])^(a[92] & b[72])^(a[91] & b[73])^(a[90] & b[74])^(a[89] & b[75])^(a[88] & b[76])^(a[87] & b[77])^(a[86] & b[78])^(a[85] & b[79])^(a[84] & b[80])^(a[83] & b[81])^(a[82] & b[82])^(a[81] & b[83])^(a[80] & b[84])^(a[79] & b[85])^(a[78] & b[86])^(a[77] & b[87])^(a[76] & b[88])^(a[75] & b[89])^(a[74] & b[90])^(a[73] & b[91])^(a[72] & b[92])^(a[71] & b[93])^(a[70] & b[94])^(a[69] & b[95])^(a[68] & b[96])^(a[67] & b[97])^(a[66] & b[98])^(a[65] & b[99])^(a[64] & b[100])^(a[63] & b[101])^(a[62] & b[102])^(a[61] & b[103])^(a[60] & b[104])^(a[59] & b[105])^(a[58] & b[106])^(a[57] & b[107])^(a[56] & b[108])^(a[55] & b[109])^(a[54] & b[110])^(a[53] & b[111])^(a[52] & b[112])^(a[51] & b[113])^(a[50] & b[114])^(a[49] & b[115])^(a[48] & b[116])^(a[47] & b[117])^(a[46] & b[118])^(a[45] & b[119])^(a[44] & b[120])^(a[43] & b[121])^(a[42] & b[122])^(a[41] & b[123])^(a[40] & b[124])^(a[39] & b[125])^(a[38] & b[126])^(a[37] & b[127])^(a[36] & b[128])^(a[35] & b[129])^(a[34] & b[130])^(a[33] & b[131])^(a[32] & b[132])^(a[31] & b[133])^(a[30] & b[134])^(a[29] & b[135])^(a[28] & b[136])^(a[27] & b[137])^(a[26] & b[138])^(a[25] & b[139])^(a[24] & b[140])^(a[23] & b[141])^(a[22] & b[142])^(a[21] & b[143])^(a[20] & b[144])^(a[19] & b[145])^(a[18] & b[146])^(a[17] & b[147])^(a[16] & b[148])^(a[15] & b[149])^(a[14] & b[150])^(a[13] & b[151])^(a[12] & b[152])^(a[11] & b[153])^(a[10] & b[154])^(a[9] & b[155])^(a[8] & b[156])^(a[7] & b[157])^(a[6] & b[158])^(a[5] & b[159])^(a[4] & b[160])^(a[3] & b[161])^(a[2] & b[162]);
assign y[165] = (a[162] & b[3])^(a[161] & b[4])^(a[160] & b[5])^(a[159] & b[6])^(a[158] & b[7])^(a[157] & b[8])^(a[156] & b[9])^(a[155] & b[10])^(a[154] & b[11])^(a[153] & b[12])^(a[152] & b[13])^(a[151] & b[14])^(a[150] & b[15])^(a[149] & b[16])^(a[148] & b[17])^(a[147] & b[18])^(a[146] & b[19])^(a[145] & b[20])^(a[144] & b[21])^(a[143] & b[22])^(a[142] & b[23])^(a[141] & b[24])^(a[140] & b[25])^(a[139] & b[26])^(a[138] & b[27])^(a[137] & b[28])^(a[136] & b[29])^(a[135] & b[30])^(a[134] & b[31])^(a[133] & b[32])^(a[132] & b[33])^(a[131] & b[34])^(a[130] & b[35])^(a[129] & b[36])^(a[128] & b[37])^(a[127] & b[38])^(a[126] & b[39])^(a[125] & b[40])^(a[124] & b[41])^(a[123] & b[42])^(a[122] & b[43])^(a[121] & b[44])^(a[120] & b[45])^(a[119] & b[46])^(a[118] & b[47])^(a[117] & b[48])^(a[116] & b[49])^(a[115] & b[50])^(a[114] & b[51])^(a[113] & b[52])^(a[112] & b[53])^(a[111] & b[54])^(a[110] & b[55])^(a[109] & b[56])^(a[108] & b[57])^(a[107] & b[58])^(a[106] & b[59])^(a[105] & b[60])^(a[104] & b[61])^(a[103] & b[62])^(a[102] & b[63])^(a[101] & b[64])^(a[100] & b[65])^(a[99] & b[66])^(a[98] & b[67])^(a[97] & b[68])^(a[96] & b[69])^(a[95] & b[70])^(a[94] & b[71])^(a[93] & b[72])^(a[92] & b[73])^(a[91] & b[74])^(a[90] & b[75])^(a[89] & b[76])^(a[88] & b[77])^(a[87] & b[78])^(a[86] & b[79])^(a[85] & b[80])^(a[84] & b[81])^(a[83] & b[82])^(a[82] & b[83])^(a[81] & b[84])^(a[80] & b[85])^(a[79] & b[86])^(a[78] & b[87])^(a[77] & b[88])^(a[76] & b[89])^(a[75] & b[90])^(a[74] & b[91])^(a[73] & b[92])^(a[72] & b[93])^(a[71] & b[94])^(a[70] & b[95])^(a[69] & b[96])^(a[68] & b[97])^(a[67] & b[98])^(a[66] & b[99])^(a[65] & b[100])^(a[64] & b[101])^(a[63] & b[102])^(a[62] & b[103])^(a[61] & b[104])^(a[60] & b[105])^(a[59] & b[106])^(a[58] & b[107])^(a[57] & b[108])^(a[56] & b[109])^(a[55] & b[110])^(a[54] & b[111])^(a[53] & b[112])^(a[52] & b[113])^(a[51] & b[114])^(a[50] & b[115])^(a[49] & b[116])^(a[48] & b[117])^(a[47] & b[118])^(a[46] & b[119])^(a[45] & b[120])^(a[44] & b[121])^(a[43] & b[122])^(a[42] & b[123])^(a[41] & b[124])^(a[40] & b[125])^(a[39] & b[126])^(a[38] & b[127])^(a[37] & b[128])^(a[36] & b[129])^(a[35] & b[130])^(a[34] & b[131])^(a[33] & b[132])^(a[32] & b[133])^(a[31] & b[134])^(a[30] & b[135])^(a[29] & b[136])^(a[28] & b[137])^(a[27] & b[138])^(a[26] & b[139])^(a[25] & b[140])^(a[24] & b[141])^(a[23] & b[142])^(a[22] & b[143])^(a[21] & b[144])^(a[20] & b[145])^(a[19] & b[146])^(a[18] & b[147])^(a[17] & b[148])^(a[16] & b[149])^(a[15] & b[150])^(a[14] & b[151])^(a[13] & b[152])^(a[12] & b[153])^(a[11] & b[154])^(a[10] & b[155])^(a[9] & b[156])^(a[8] & b[157])^(a[7] & b[158])^(a[6] & b[159])^(a[5] & b[160])^(a[4] & b[161])^(a[3] & b[162]);
assign y[166] = (a[162] & b[4])^(a[161] & b[5])^(a[160] & b[6])^(a[159] & b[7])^(a[158] & b[8])^(a[157] & b[9])^(a[156] & b[10])^(a[155] & b[11])^(a[154] & b[12])^(a[153] & b[13])^(a[152] & b[14])^(a[151] & b[15])^(a[150] & b[16])^(a[149] & b[17])^(a[148] & b[18])^(a[147] & b[19])^(a[146] & b[20])^(a[145] & b[21])^(a[144] & b[22])^(a[143] & b[23])^(a[142] & b[24])^(a[141] & b[25])^(a[140] & b[26])^(a[139] & b[27])^(a[138] & b[28])^(a[137] & b[29])^(a[136] & b[30])^(a[135] & b[31])^(a[134] & b[32])^(a[133] & b[33])^(a[132] & b[34])^(a[131] & b[35])^(a[130] & b[36])^(a[129] & b[37])^(a[128] & b[38])^(a[127] & b[39])^(a[126] & b[40])^(a[125] & b[41])^(a[124] & b[42])^(a[123] & b[43])^(a[122] & b[44])^(a[121] & b[45])^(a[120] & b[46])^(a[119] & b[47])^(a[118] & b[48])^(a[117] & b[49])^(a[116] & b[50])^(a[115] & b[51])^(a[114] & b[52])^(a[113] & b[53])^(a[112] & b[54])^(a[111] & b[55])^(a[110] & b[56])^(a[109] & b[57])^(a[108] & b[58])^(a[107] & b[59])^(a[106] & b[60])^(a[105] & b[61])^(a[104] & b[62])^(a[103] & b[63])^(a[102] & b[64])^(a[101] & b[65])^(a[100] & b[66])^(a[99] & b[67])^(a[98] & b[68])^(a[97] & b[69])^(a[96] & b[70])^(a[95] & b[71])^(a[94] & b[72])^(a[93] & b[73])^(a[92] & b[74])^(a[91] & b[75])^(a[90] & b[76])^(a[89] & b[77])^(a[88] & b[78])^(a[87] & b[79])^(a[86] & b[80])^(a[85] & b[81])^(a[84] & b[82])^(a[83] & b[83])^(a[82] & b[84])^(a[81] & b[85])^(a[80] & b[86])^(a[79] & b[87])^(a[78] & b[88])^(a[77] & b[89])^(a[76] & b[90])^(a[75] & b[91])^(a[74] & b[92])^(a[73] & b[93])^(a[72] & b[94])^(a[71] & b[95])^(a[70] & b[96])^(a[69] & b[97])^(a[68] & b[98])^(a[67] & b[99])^(a[66] & b[100])^(a[65] & b[101])^(a[64] & b[102])^(a[63] & b[103])^(a[62] & b[104])^(a[61] & b[105])^(a[60] & b[106])^(a[59] & b[107])^(a[58] & b[108])^(a[57] & b[109])^(a[56] & b[110])^(a[55] & b[111])^(a[54] & b[112])^(a[53] & b[113])^(a[52] & b[114])^(a[51] & b[115])^(a[50] & b[116])^(a[49] & b[117])^(a[48] & b[118])^(a[47] & b[119])^(a[46] & b[120])^(a[45] & b[121])^(a[44] & b[122])^(a[43] & b[123])^(a[42] & b[124])^(a[41] & b[125])^(a[40] & b[126])^(a[39] & b[127])^(a[38] & b[128])^(a[37] & b[129])^(a[36] & b[130])^(a[35] & b[131])^(a[34] & b[132])^(a[33] & b[133])^(a[32] & b[134])^(a[31] & b[135])^(a[30] & b[136])^(a[29] & b[137])^(a[28] & b[138])^(a[27] & b[139])^(a[26] & b[140])^(a[25] & b[141])^(a[24] & b[142])^(a[23] & b[143])^(a[22] & b[144])^(a[21] & b[145])^(a[20] & b[146])^(a[19] & b[147])^(a[18] & b[148])^(a[17] & b[149])^(a[16] & b[150])^(a[15] & b[151])^(a[14] & b[152])^(a[13] & b[153])^(a[12] & b[154])^(a[11] & b[155])^(a[10] & b[156])^(a[9] & b[157])^(a[8] & b[158])^(a[7] & b[159])^(a[6] & b[160])^(a[5] & b[161])^(a[4] & b[162]);
assign y[167] = (a[162] & b[5])^(a[161] & b[6])^(a[160] & b[7])^(a[159] & b[8])^(a[158] & b[9])^(a[157] & b[10])^(a[156] & b[11])^(a[155] & b[12])^(a[154] & b[13])^(a[153] & b[14])^(a[152] & b[15])^(a[151] & b[16])^(a[150] & b[17])^(a[149] & b[18])^(a[148] & b[19])^(a[147] & b[20])^(a[146] & b[21])^(a[145] & b[22])^(a[144] & b[23])^(a[143] & b[24])^(a[142] & b[25])^(a[141] & b[26])^(a[140] & b[27])^(a[139] & b[28])^(a[138] & b[29])^(a[137] & b[30])^(a[136] & b[31])^(a[135] & b[32])^(a[134] & b[33])^(a[133] & b[34])^(a[132] & b[35])^(a[131] & b[36])^(a[130] & b[37])^(a[129] & b[38])^(a[128] & b[39])^(a[127] & b[40])^(a[126] & b[41])^(a[125] & b[42])^(a[124] & b[43])^(a[123] & b[44])^(a[122] & b[45])^(a[121] & b[46])^(a[120] & b[47])^(a[119] & b[48])^(a[118] & b[49])^(a[117] & b[50])^(a[116] & b[51])^(a[115] & b[52])^(a[114] & b[53])^(a[113] & b[54])^(a[112] & b[55])^(a[111] & b[56])^(a[110] & b[57])^(a[109] & b[58])^(a[108] & b[59])^(a[107] & b[60])^(a[106] & b[61])^(a[105] & b[62])^(a[104] & b[63])^(a[103] & b[64])^(a[102] & b[65])^(a[101] & b[66])^(a[100] & b[67])^(a[99] & b[68])^(a[98] & b[69])^(a[97] & b[70])^(a[96] & b[71])^(a[95] & b[72])^(a[94] & b[73])^(a[93] & b[74])^(a[92] & b[75])^(a[91] & b[76])^(a[90] & b[77])^(a[89] & b[78])^(a[88] & b[79])^(a[87] & b[80])^(a[86] & b[81])^(a[85] & b[82])^(a[84] & b[83])^(a[83] & b[84])^(a[82] & b[85])^(a[81] & b[86])^(a[80] & b[87])^(a[79] & b[88])^(a[78] & b[89])^(a[77] & b[90])^(a[76] & b[91])^(a[75] & b[92])^(a[74] & b[93])^(a[73] & b[94])^(a[72] & b[95])^(a[71] & b[96])^(a[70] & b[97])^(a[69] & b[98])^(a[68] & b[99])^(a[67] & b[100])^(a[66] & b[101])^(a[65] & b[102])^(a[64] & b[103])^(a[63] & b[104])^(a[62] & b[105])^(a[61] & b[106])^(a[60] & b[107])^(a[59] & b[108])^(a[58] & b[109])^(a[57] & b[110])^(a[56] & b[111])^(a[55] & b[112])^(a[54] & b[113])^(a[53] & b[114])^(a[52] & b[115])^(a[51] & b[116])^(a[50] & b[117])^(a[49] & b[118])^(a[48] & b[119])^(a[47] & b[120])^(a[46] & b[121])^(a[45] & b[122])^(a[44] & b[123])^(a[43] & b[124])^(a[42] & b[125])^(a[41] & b[126])^(a[40] & b[127])^(a[39] & b[128])^(a[38] & b[129])^(a[37] & b[130])^(a[36] & b[131])^(a[35] & b[132])^(a[34] & b[133])^(a[33] & b[134])^(a[32] & b[135])^(a[31] & b[136])^(a[30] & b[137])^(a[29] & b[138])^(a[28] & b[139])^(a[27] & b[140])^(a[26] & b[141])^(a[25] & b[142])^(a[24] & b[143])^(a[23] & b[144])^(a[22] & b[145])^(a[21] & b[146])^(a[20] & b[147])^(a[19] & b[148])^(a[18] & b[149])^(a[17] & b[150])^(a[16] & b[151])^(a[15] & b[152])^(a[14] & b[153])^(a[13] & b[154])^(a[12] & b[155])^(a[11] & b[156])^(a[10] & b[157])^(a[9] & b[158])^(a[8] & b[159])^(a[7] & b[160])^(a[6] & b[161])^(a[5] & b[162]);
assign y[168] = (a[162] & b[6])^(a[161] & b[7])^(a[160] & b[8])^(a[159] & b[9])^(a[158] & b[10])^(a[157] & b[11])^(a[156] & b[12])^(a[155] & b[13])^(a[154] & b[14])^(a[153] & b[15])^(a[152] & b[16])^(a[151] & b[17])^(a[150] & b[18])^(a[149] & b[19])^(a[148] & b[20])^(a[147] & b[21])^(a[146] & b[22])^(a[145] & b[23])^(a[144] & b[24])^(a[143] & b[25])^(a[142] & b[26])^(a[141] & b[27])^(a[140] & b[28])^(a[139] & b[29])^(a[138] & b[30])^(a[137] & b[31])^(a[136] & b[32])^(a[135] & b[33])^(a[134] & b[34])^(a[133] & b[35])^(a[132] & b[36])^(a[131] & b[37])^(a[130] & b[38])^(a[129] & b[39])^(a[128] & b[40])^(a[127] & b[41])^(a[126] & b[42])^(a[125] & b[43])^(a[124] & b[44])^(a[123] & b[45])^(a[122] & b[46])^(a[121] & b[47])^(a[120] & b[48])^(a[119] & b[49])^(a[118] & b[50])^(a[117] & b[51])^(a[116] & b[52])^(a[115] & b[53])^(a[114] & b[54])^(a[113] & b[55])^(a[112] & b[56])^(a[111] & b[57])^(a[110] & b[58])^(a[109] & b[59])^(a[108] & b[60])^(a[107] & b[61])^(a[106] & b[62])^(a[105] & b[63])^(a[104] & b[64])^(a[103] & b[65])^(a[102] & b[66])^(a[101] & b[67])^(a[100] & b[68])^(a[99] & b[69])^(a[98] & b[70])^(a[97] & b[71])^(a[96] & b[72])^(a[95] & b[73])^(a[94] & b[74])^(a[93] & b[75])^(a[92] & b[76])^(a[91] & b[77])^(a[90] & b[78])^(a[89] & b[79])^(a[88] & b[80])^(a[87] & b[81])^(a[86] & b[82])^(a[85] & b[83])^(a[84] & b[84])^(a[83] & b[85])^(a[82] & b[86])^(a[81] & b[87])^(a[80] & b[88])^(a[79] & b[89])^(a[78] & b[90])^(a[77] & b[91])^(a[76] & b[92])^(a[75] & b[93])^(a[74] & b[94])^(a[73] & b[95])^(a[72] & b[96])^(a[71] & b[97])^(a[70] & b[98])^(a[69] & b[99])^(a[68] & b[100])^(a[67] & b[101])^(a[66] & b[102])^(a[65] & b[103])^(a[64] & b[104])^(a[63] & b[105])^(a[62] & b[106])^(a[61] & b[107])^(a[60] & b[108])^(a[59] & b[109])^(a[58] & b[110])^(a[57] & b[111])^(a[56] & b[112])^(a[55] & b[113])^(a[54] & b[114])^(a[53] & b[115])^(a[52] & b[116])^(a[51] & b[117])^(a[50] & b[118])^(a[49] & b[119])^(a[48] & b[120])^(a[47] & b[121])^(a[46] & b[122])^(a[45] & b[123])^(a[44] & b[124])^(a[43] & b[125])^(a[42] & b[126])^(a[41] & b[127])^(a[40] & b[128])^(a[39] & b[129])^(a[38] & b[130])^(a[37] & b[131])^(a[36] & b[132])^(a[35] & b[133])^(a[34] & b[134])^(a[33] & b[135])^(a[32] & b[136])^(a[31] & b[137])^(a[30] & b[138])^(a[29] & b[139])^(a[28] & b[140])^(a[27] & b[141])^(a[26] & b[142])^(a[25] & b[143])^(a[24] & b[144])^(a[23] & b[145])^(a[22] & b[146])^(a[21] & b[147])^(a[20] & b[148])^(a[19] & b[149])^(a[18] & b[150])^(a[17] & b[151])^(a[16] & b[152])^(a[15] & b[153])^(a[14] & b[154])^(a[13] & b[155])^(a[12] & b[156])^(a[11] & b[157])^(a[10] & b[158])^(a[9] & b[159])^(a[8] & b[160])^(a[7] & b[161])^(a[6] & b[162]);
assign y[169] = (a[162] & b[7])^(a[161] & b[8])^(a[160] & b[9])^(a[159] & b[10])^(a[158] & b[11])^(a[157] & b[12])^(a[156] & b[13])^(a[155] & b[14])^(a[154] & b[15])^(a[153] & b[16])^(a[152] & b[17])^(a[151] & b[18])^(a[150] & b[19])^(a[149] & b[20])^(a[148] & b[21])^(a[147] & b[22])^(a[146] & b[23])^(a[145] & b[24])^(a[144] & b[25])^(a[143] & b[26])^(a[142] & b[27])^(a[141] & b[28])^(a[140] & b[29])^(a[139] & b[30])^(a[138] & b[31])^(a[137] & b[32])^(a[136] & b[33])^(a[135] & b[34])^(a[134] & b[35])^(a[133] & b[36])^(a[132] & b[37])^(a[131] & b[38])^(a[130] & b[39])^(a[129] & b[40])^(a[128] & b[41])^(a[127] & b[42])^(a[126] & b[43])^(a[125] & b[44])^(a[124] & b[45])^(a[123] & b[46])^(a[122] & b[47])^(a[121] & b[48])^(a[120] & b[49])^(a[119] & b[50])^(a[118] & b[51])^(a[117] & b[52])^(a[116] & b[53])^(a[115] & b[54])^(a[114] & b[55])^(a[113] & b[56])^(a[112] & b[57])^(a[111] & b[58])^(a[110] & b[59])^(a[109] & b[60])^(a[108] & b[61])^(a[107] & b[62])^(a[106] & b[63])^(a[105] & b[64])^(a[104] & b[65])^(a[103] & b[66])^(a[102] & b[67])^(a[101] & b[68])^(a[100] & b[69])^(a[99] & b[70])^(a[98] & b[71])^(a[97] & b[72])^(a[96] & b[73])^(a[95] & b[74])^(a[94] & b[75])^(a[93] & b[76])^(a[92] & b[77])^(a[91] & b[78])^(a[90] & b[79])^(a[89] & b[80])^(a[88] & b[81])^(a[87] & b[82])^(a[86] & b[83])^(a[85] & b[84])^(a[84] & b[85])^(a[83] & b[86])^(a[82] & b[87])^(a[81] & b[88])^(a[80] & b[89])^(a[79] & b[90])^(a[78] & b[91])^(a[77] & b[92])^(a[76] & b[93])^(a[75] & b[94])^(a[74] & b[95])^(a[73] & b[96])^(a[72] & b[97])^(a[71] & b[98])^(a[70] & b[99])^(a[69] & b[100])^(a[68] & b[101])^(a[67] & b[102])^(a[66] & b[103])^(a[65] & b[104])^(a[64] & b[105])^(a[63] & b[106])^(a[62] & b[107])^(a[61] & b[108])^(a[60] & b[109])^(a[59] & b[110])^(a[58] & b[111])^(a[57] & b[112])^(a[56] & b[113])^(a[55] & b[114])^(a[54] & b[115])^(a[53] & b[116])^(a[52] & b[117])^(a[51] & b[118])^(a[50] & b[119])^(a[49] & b[120])^(a[48] & b[121])^(a[47] & b[122])^(a[46] & b[123])^(a[45] & b[124])^(a[44] & b[125])^(a[43] & b[126])^(a[42] & b[127])^(a[41] & b[128])^(a[40] & b[129])^(a[39] & b[130])^(a[38] & b[131])^(a[37] & b[132])^(a[36] & b[133])^(a[35] & b[134])^(a[34] & b[135])^(a[33] & b[136])^(a[32] & b[137])^(a[31] & b[138])^(a[30] & b[139])^(a[29] & b[140])^(a[28] & b[141])^(a[27] & b[142])^(a[26] & b[143])^(a[25] & b[144])^(a[24] & b[145])^(a[23] & b[146])^(a[22] & b[147])^(a[21] & b[148])^(a[20] & b[149])^(a[19] & b[150])^(a[18] & b[151])^(a[17] & b[152])^(a[16] & b[153])^(a[15] & b[154])^(a[14] & b[155])^(a[13] & b[156])^(a[12] & b[157])^(a[11] & b[158])^(a[10] & b[159])^(a[9] & b[160])^(a[8] & b[161])^(a[7] & b[162]);
assign y[170] = (a[162] & b[8])^(a[161] & b[9])^(a[160] & b[10])^(a[159] & b[11])^(a[158] & b[12])^(a[157] & b[13])^(a[156] & b[14])^(a[155] & b[15])^(a[154] & b[16])^(a[153] & b[17])^(a[152] & b[18])^(a[151] & b[19])^(a[150] & b[20])^(a[149] & b[21])^(a[148] & b[22])^(a[147] & b[23])^(a[146] & b[24])^(a[145] & b[25])^(a[144] & b[26])^(a[143] & b[27])^(a[142] & b[28])^(a[141] & b[29])^(a[140] & b[30])^(a[139] & b[31])^(a[138] & b[32])^(a[137] & b[33])^(a[136] & b[34])^(a[135] & b[35])^(a[134] & b[36])^(a[133] & b[37])^(a[132] & b[38])^(a[131] & b[39])^(a[130] & b[40])^(a[129] & b[41])^(a[128] & b[42])^(a[127] & b[43])^(a[126] & b[44])^(a[125] & b[45])^(a[124] & b[46])^(a[123] & b[47])^(a[122] & b[48])^(a[121] & b[49])^(a[120] & b[50])^(a[119] & b[51])^(a[118] & b[52])^(a[117] & b[53])^(a[116] & b[54])^(a[115] & b[55])^(a[114] & b[56])^(a[113] & b[57])^(a[112] & b[58])^(a[111] & b[59])^(a[110] & b[60])^(a[109] & b[61])^(a[108] & b[62])^(a[107] & b[63])^(a[106] & b[64])^(a[105] & b[65])^(a[104] & b[66])^(a[103] & b[67])^(a[102] & b[68])^(a[101] & b[69])^(a[100] & b[70])^(a[99] & b[71])^(a[98] & b[72])^(a[97] & b[73])^(a[96] & b[74])^(a[95] & b[75])^(a[94] & b[76])^(a[93] & b[77])^(a[92] & b[78])^(a[91] & b[79])^(a[90] & b[80])^(a[89] & b[81])^(a[88] & b[82])^(a[87] & b[83])^(a[86] & b[84])^(a[85] & b[85])^(a[84] & b[86])^(a[83] & b[87])^(a[82] & b[88])^(a[81] & b[89])^(a[80] & b[90])^(a[79] & b[91])^(a[78] & b[92])^(a[77] & b[93])^(a[76] & b[94])^(a[75] & b[95])^(a[74] & b[96])^(a[73] & b[97])^(a[72] & b[98])^(a[71] & b[99])^(a[70] & b[100])^(a[69] & b[101])^(a[68] & b[102])^(a[67] & b[103])^(a[66] & b[104])^(a[65] & b[105])^(a[64] & b[106])^(a[63] & b[107])^(a[62] & b[108])^(a[61] & b[109])^(a[60] & b[110])^(a[59] & b[111])^(a[58] & b[112])^(a[57] & b[113])^(a[56] & b[114])^(a[55] & b[115])^(a[54] & b[116])^(a[53] & b[117])^(a[52] & b[118])^(a[51] & b[119])^(a[50] & b[120])^(a[49] & b[121])^(a[48] & b[122])^(a[47] & b[123])^(a[46] & b[124])^(a[45] & b[125])^(a[44] & b[126])^(a[43] & b[127])^(a[42] & b[128])^(a[41] & b[129])^(a[40] & b[130])^(a[39] & b[131])^(a[38] & b[132])^(a[37] & b[133])^(a[36] & b[134])^(a[35] & b[135])^(a[34] & b[136])^(a[33] & b[137])^(a[32] & b[138])^(a[31] & b[139])^(a[30] & b[140])^(a[29] & b[141])^(a[28] & b[142])^(a[27] & b[143])^(a[26] & b[144])^(a[25] & b[145])^(a[24] & b[146])^(a[23] & b[147])^(a[22] & b[148])^(a[21] & b[149])^(a[20] & b[150])^(a[19] & b[151])^(a[18] & b[152])^(a[17] & b[153])^(a[16] & b[154])^(a[15] & b[155])^(a[14] & b[156])^(a[13] & b[157])^(a[12] & b[158])^(a[11] & b[159])^(a[10] & b[160])^(a[9] & b[161])^(a[8] & b[162]);
assign y[171] = (a[162] & b[9])^(a[161] & b[10])^(a[160] & b[11])^(a[159] & b[12])^(a[158] & b[13])^(a[157] & b[14])^(a[156] & b[15])^(a[155] & b[16])^(a[154] & b[17])^(a[153] & b[18])^(a[152] & b[19])^(a[151] & b[20])^(a[150] & b[21])^(a[149] & b[22])^(a[148] & b[23])^(a[147] & b[24])^(a[146] & b[25])^(a[145] & b[26])^(a[144] & b[27])^(a[143] & b[28])^(a[142] & b[29])^(a[141] & b[30])^(a[140] & b[31])^(a[139] & b[32])^(a[138] & b[33])^(a[137] & b[34])^(a[136] & b[35])^(a[135] & b[36])^(a[134] & b[37])^(a[133] & b[38])^(a[132] & b[39])^(a[131] & b[40])^(a[130] & b[41])^(a[129] & b[42])^(a[128] & b[43])^(a[127] & b[44])^(a[126] & b[45])^(a[125] & b[46])^(a[124] & b[47])^(a[123] & b[48])^(a[122] & b[49])^(a[121] & b[50])^(a[120] & b[51])^(a[119] & b[52])^(a[118] & b[53])^(a[117] & b[54])^(a[116] & b[55])^(a[115] & b[56])^(a[114] & b[57])^(a[113] & b[58])^(a[112] & b[59])^(a[111] & b[60])^(a[110] & b[61])^(a[109] & b[62])^(a[108] & b[63])^(a[107] & b[64])^(a[106] & b[65])^(a[105] & b[66])^(a[104] & b[67])^(a[103] & b[68])^(a[102] & b[69])^(a[101] & b[70])^(a[100] & b[71])^(a[99] & b[72])^(a[98] & b[73])^(a[97] & b[74])^(a[96] & b[75])^(a[95] & b[76])^(a[94] & b[77])^(a[93] & b[78])^(a[92] & b[79])^(a[91] & b[80])^(a[90] & b[81])^(a[89] & b[82])^(a[88] & b[83])^(a[87] & b[84])^(a[86] & b[85])^(a[85] & b[86])^(a[84] & b[87])^(a[83] & b[88])^(a[82] & b[89])^(a[81] & b[90])^(a[80] & b[91])^(a[79] & b[92])^(a[78] & b[93])^(a[77] & b[94])^(a[76] & b[95])^(a[75] & b[96])^(a[74] & b[97])^(a[73] & b[98])^(a[72] & b[99])^(a[71] & b[100])^(a[70] & b[101])^(a[69] & b[102])^(a[68] & b[103])^(a[67] & b[104])^(a[66] & b[105])^(a[65] & b[106])^(a[64] & b[107])^(a[63] & b[108])^(a[62] & b[109])^(a[61] & b[110])^(a[60] & b[111])^(a[59] & b[112])^(a[58] & b[113])^(a[57] & b[114])^(a[56] & b[115])^(a[55] & b[116])^(a[54] & b[117])^(a[53] & b[118])^(a[52] & b[119])^(a[51] & b[120])^(a[50] & b[121])^(a[49] & b[122])^(a[48] & b[123])^(a[47] & b[124])^(a[46] & b[125])^(a[45] & b[126])^(a[44] & b[127])^(a[43] & b[128])^(a[42] & b[129])^(a[41] & b[130])^(a[40] & b[131])^(a[39] & b[132])^(a[38] & b[133])^(a[37] & b[134])^(a[36] & b[135])^(a[35] & b[136])^(a[34] & b[137])^(a[33] & b[138])^(a[32] & b[139])^(a[31] & b[140])^(a[30] & b[141])^(a[29] & b[142])^(a[28] & b[143])^(a[27] & b[144])^(a[26] & b[145])^(a[25] & b[146])^(a[24] & b[147])^(a[23] & b[148])^(a[22] & b[149])^(a[21] & b[150])^(a[20] & b[151])^(a[19] & b[152])^(a[18] & b[153])^(a[17] & b[154])^(a[16] & b[155])^(a[15] & b[156])^(a[14] & b[157])^(a[13] & b[158])^(a[12] & b[159])^(a[11] & b[160])^(a[10] & b[161])^(a[9] & b[162]);
assign y[172] = (a[162] & b[10])^(a[161] & b[11])^(a[160] & b[12])^(a[159] & b[13])^(a[158] & b[14])^(a[157] & b[15])^(a[156] & b[16])^(a[155] & b[17])^(a[154] & b[18])^(a[153] & b[19])^(a[152] & b[20])^(a[151] & b[21])^(a[150] & b[22])^(a[149] & b[23])^(a[148] & b[24])^(a[147] & b[25])^(a[146] & b[26])^(a[145] & b[27])^(a[144] & b[28])^(a[143] & b[29])^(a[142] & b[30])^(a[141] & b[31])^(a[140] & b[32])^(a[139] & b[33])^(a[138] & b[34])^(a[137] & b[35])^(a[136] & b[36])^(a[135] & b[37])^(a[134] & b[38])^(a[133] & b[39])^(a[132] & b[40])^(a[131] & b[41])^(a[130] & b[42])^(a[129] & b[43])^(a[128] & b[44])^(a[127] & b[45])^(a[126] & b[46])^(a[125] & b[47])^(a[124] & b[48])^(a[123] & b[49])^(a[122] & b[50])^(a[121] & b[51])^(a[120] & b[52])^(a[119] & b[53])^(a[118] & b[54])^(a[117] & b[55])^(a[116] & b[56])^(a[115] & b[57])^(a[114] & b[58])^(a[113] & b[59])^(a[112] & b[60])^(a[111] & b[61])^(a[110] & b[62])^(a[109] & b[63])^(a[108] & b[64])^(a[107] & b[65])^(a[106] & b[66])^(a[105] & b[67])^(a[104] & b[68])^(a[103] & b[69])^(a[102] & b[70])^(a[101] & b[71])^(a[100] & b[72])^(a[99] & b[73])^(a[98] & b[74])^(a[97] & b[75])^(a[96] & b[76])^(a[95] & b[77])^(a[94] & b[78])^(a[93] & b[79])^(a[92] & b[80])^(a[91] & b[81])^(a[90] & b[82])^(a[89] & b[83])^(a[88] & b[84])^(a[87] & b[85])^(a[86] & b[86])^(a[85] & b[87])^(a[84] & b[88])^(a[83] & b[89])^(a[82] & b[90])^(a[81] & b[91])^(a[80] & b[92])^(a[79] & b[93])^(a[78] & b[94])^(a[77] & b[95])^(a[76] & b[96])^(a[75] & b[97])^(a[74] & b[98])^(a[73] & b[99])^(a[72] & b[100])^(a[71] & b[101])^(a[70] & b[102])^(a[69] & b[103])^(a[68] & b[104])^(a[67] & b[105])^(a[66] & b[106])^(a[65] & b[107])^(a[64] & b[108])^(a[63] & b[109])^(a[62] & b[110])^(a[61] & b[111])^(a[60] & b[112])^(a[59] & b[113])^(a[58] & b[114])^(a[57] & b[115])^(a[56] & b[116])^(a[55] & b[117])^(a[54] & b[118])^(a[53] & b[119])^(a[52] & b[120])^(a[51] & b[121])^(a[50] & b[122])^(a[49] & b[123])^(a[48] & b[124])^(a[47] & b[125])^(a[46] & b[126])^(a[45] & b[127])^(a[44] & b[128])^(a[43] & b[129])^(a[42] & b[130])^(a[41] & b[131])^(a[40] & b[132])^(a[39] & b[133])^(a[38] & b[134])^(a[37] & b[135])^(a[36] & b[136])^(a[35] & b[137])^(a[34] & b[138])^(a[33] & b[139])^(a[32] & b[140])^(a[31] & b[141])^(a[30] & b[142])^(a[29] & b[143])^(a[28] & b[144])^(a[27] & b[145])^(a[26] & b[146])^(a[25] & b[147])^(a[24] & b[148])^(a[23] & b[149])^(a[22] & b[150])^(a[21] & b[151])^(a[20] & b[152])^(a[19] & b[153])^(a[18] & b[154])^(a[17] & b[155])^(a[16] & b[156])^(a[15] & b[157])^(a[14] & b[158])^(a[13] & b[159])^(a[12] & b[160])^(a[11] & b[161])^(a[10] & b[162]);
assign y[173] = (a[162] & b[11])^(a[161] & b[12])^(a[160] & b[13])^(a[159] & b[14])^(a[158] & b[15])^(a[157] & b[16])^(a[156] & b[17])^(a[155] & b[18])^(a[154] & b[19])^(a[153] & b[20])^(a[152] & b[21])^(a[151] & b[22])^(a[150] & b[23])^(a[149] & b[24])^(a[148] & b[25])^(a[147] & b[26])^(a[146] & b[27])^(a[145] & b[28])^(a[144] & b[29])^(a[143] & b[30])^(a[142] & b[31])^(a[141] & b[32])^(a[140] & b[33])^(a[139] & b[34])^(a[138] & b[35])^(a[137] & b[36])^(a[136] & b[37])^(a[135] & b[38])^(a[134] & b[39])^(a[133] & b[40])^(a[132] & b[41])^(a[131] & b[42])^(a[130] & b[43])^(a[129] & b[44])^(a[128] & b[45])^(a[127] & b[46])^(a[126] & b[47])^(a[125] & b[48])^(a[124] & b[49])^(a[123] & b[50])^(a[122] & b[51])^(a[121] & b[52])^(a[120] & b[53])^(a[119] & b[54])^(a[118] & b[55])^(a[117] & b[56])^(a[116] & b[57])^(a[115] & b[58])^(a[114] & b[59])^(a[113] & b[60])^(a[112] & b[61])^(a[111] & b[62])^(a[110] & b[63])^(a[109] & b[64])^(a[108] & b[65])^(a[107] & b[66])^(a[106] & b[67])^(a[105] & b[68])^(a[104] & b[69])^(a[103] & b[70])^(a[102] & b[71])^(a[101] & b[72])^(a[100] & b[73])^(a[99] & b[74])^(a[98] & b[75])^(a[97] & b[76])^(a[96] & b[77])^(a[95] & b[78])^(a[94] & b[79])^(a[93] & b[80])^(a[92] & b[81])^(a[91] & b[82])^(a[90] & b[83])^(a[89] & b[84])^(a[88] & b[85])^(a[87] & b[86])^(a[86] & b[87])^(a[85] & b[88])^(a[84] & b[89])^(a[83] & b[90])^(a[82] & b[91])^(a[81] & b[92])^(a[80] & b[93])^(a[79] & b[94])^(a[78] & b[95])^(a[77] & b[96])^(a[76] & b[97])^(a[75] & b[98])^(a[74] & b[99])^(a[73] & b[100])^(a[72] & b[101])^(a[71] & b[102])^(a[70] & b[103])^(a[69] & b[104])^(a[68] & b[105])^(a[67] & b[106])^(a[66] & b[107])^(a[65] & b[108])^(a[64] & b[109])^(a[63] & b[110])^(a[62] & b[111])^(a[61] & b[112])^(a[60] & b[113])^(a[59] & b[114])^(a[58] & b[115])^(a[57] & b[116])^(a[56] & b[117])^(a[55] & b[118])^(a[54] & b[119])^(a[53] & b[120])^(a[52] & b[121])^(a[51] & b[122])^(a[50] & b[123])^(a[49] & b[124])^(a[48] & b[125])^(a[47] & b[126])^(a[46] & b[127])^(a[45] & b[128])^(a[44] & b[129])^(a[43] & b[130])^(a[42] & b[131])^(a[41] & b[132])^(a[40] & b[133])^(a[39] & b[134])^(a[38] & b[135])^(a[37] & b[136])^(a[36] & b[137])^(a[35] & b[138])^(a[34] & b[139])^(a[33] & b[140])^(a[32] & b[141])^(a[31] & b[142])^(a[30] & b[143])^(a[29] & b[144])^(a[28] & b[145])^(a[27] & b[146])^(a[26] & b[147])^(a[25] & b[148])^(a[24] & b[149])^(a[23] & b[150])^(a[22] & b[151])^(a[21] & b[152])^(a[20] & b[153])^(a[19] & b[154])^(a[18] & b[155])^(a[17] & b[156])^(a[16] & b[157])^(a[15] & b[158])^(a[14] & b[159])^(a[13] & b[160])^(a[12] & b[161])^(a[11] & b[162]);
assign y[174] = (a[162] & b[12])^(a[161] & b[13])^(a[160] & b[14])^(a[159] & b[15])^(a[158] & b[16])^(a[157] & b[17])^(a[156] & b[18])^(a[155] & b[19])^(a[154] & b[20])^(a[153] & b[21])^(a[152] & b[22])^(a[151] & b[23])^(a[150] & b[24])^(a[149] & b[25])^(a[148] & b[26])^(a[147] & b[27])^(a[146] & b[28])^(a[145] & b[29])^(a[144] & b[30])^(a[143] & b[31])^(a[142] & b[32])^(a[141] & b[33])^(a[140] & b[34])^(a[139] & b[35])^(a[138] & b[36])^(a[137] & b[37])^(a[136] & b[38])^(a[135] & b[39])^(a[134] & b[40])^(a[133] & b[41])^(a[132] & b[42])^(a[131] & b[43])^(a[130] & b[44])^(a[129] & b[45])^(a[128] & b[46])^(a[127] & b[47])^(a[126] & b[48])^(a[125] & b[49])^(a[124] & b[50])^(a[123] & b[51])^(a[122] & b[52])^(a[121] & b[53])^(a[120] & b[54])^(a[119] & b[55])^(a[118] & b[56])^(a[117] & b[57])^(a[116] & b[58])^(a[115] & b[59])^(a[114] & b[60])^(a[113] & b[61])^(a[112] & b[62])^(a[111] & b[63])^(a[110] & b[64])^(a[109] & b[65])^(a[108] & b[66])^(a[107] & b[67])^(a[106] & b[68])^(a[105] & b[69])^(a[104] & b[70])^(a[103] & b[71])^(a[102] & b[72])^(a[101] & b[73])^(a[100] & b[74])^(a[99] & b[75])^(a[98] & b[76])^(a[97] & b[77])^(a[96] & b[78])^(a[95] & b[79])^(a[94] & b[80])^(a[93] & b[81])^(a[92] & b[82])^(a[91] & b[83])^(a[90] & b[84])^(a[89] & b[85])^(a[88] & b[86])^(a[87] & b[87])^(a[86] & b[88])^(a[85] & b[89])^(a[84] & b[90])^(a[83] & b[91])^(a[82] & b[92])^(a[81] & b[93])^(a[80] & b[94])^(a[79] & b[95])^(a[78] & b[96])^(a[77] & b[97])^(a[76] & b[98])^(a[75] & b[99])^(a[74] & b[100])^(a[73] & b[101])^(a[72] & b[102])^(a[71] & b[103])^(a[70] & b[104])^(a[69] & b[105])^(a[68] & b[106])^(a[67] & b[107])^(a[66] & b[108])^(a[65] & b[109])^(a[64] & b[110])^(a[63] & b[111])^(a[62] & b[112])^(a[61] & b[113])^(a[60] & b[114])^(a[59] & b[115])^(a[58] & b[116])^(a[57] & b[117])^(a[56] & b[118])^(a[55] & b[119])^(a[54] & b[120])^(a[53] & b[121])^(a[52] & b[122])^(a[51] & b[123])^(a[50] & b[124])^(a[49] & b[125])^(a[48] & b[126])^(a[47] & b[127])^(a[46] & b[128])^(a[45] & b[129])^(a[44] & b[130])^(a[43] & b[131])^(a[42] & b[132])^(a[41] & b[133])^(a[40] & b[134])^(a[39] & b[135])^(a[38] & b[136])^(a[37] & b[137])^(a[36] & b[138])^(a[35] & b[139])^(a[34] & b[140])^(a[33] & b[141])^(a[32] & b[142])^(a[31] & b[143])^(a[30] & b[144])^(a[29] & b[145])^(a[28] & b[146])^(a[27] & b[147])^(a[26] & b[148])^(a[25] & b[149])^(a[24] & b[150])^(a[23] & b[151])^(a[22] & b[152])^(a[21] & b[153])^(a[20] & b[154])^(a[19] & b[155])^(a[18] & b[156])^(a[17] & b[157])^(a[16] & b[158])^(a[15] & b[159])^(a[14] & b[160])^(a[13] & b[161])^(a[12] & b[162]);
assign y[175] = (a[162] & b[13])^(a[161] & b[14])^(a[160] & b[15])^(a[159] & b[16])^(a[158] & b[17])^(a[157] & b[18])^(a[156] & b[19])^(a[155] & b[20])^(a[154] & b[21])^(a[153] & b[22])^(a[152] & b[23])^(a[151] & b[24])^(a[150] & b[25])^(a[149] & b[26])^(a[148] & b[27])^(a[147] & b[28])^(a[146] & b[29])^(a[145] & b[30])^(a[144] & b[31])^(a[143] & b[32])^(a[142] & b[33])^(a[141] & b[34])^(a[140] & b[35])^(a[139] & b[36])^(a[138] & b[37])^(a[137] & b[38])^(a[136] & b[39])^(a[135] & b[40])^(a[134] & b[41])^(a[133] & b[42])^(a[132] & b[43])^(a[131] & b[44])^(a[130] & b[45])^(a[129] & b[46])^(a[128] & b[47])^(a[127] & b[48])^(a[126] & b[49])^(a[125] & b[50])^(a[124] & b[51])^(a[123] & b[52])^(a[122] & b[53])^(a[121] & b[54])^(a[120] & b[55])^(a[119] & b[56])^(a[118] & b[57])^(a[117] & b[58])^(a[116] & b[59])^(a[115] & b[60])^(a[114] & b[61])^(a[113] & b[62])^(a[112] & b[63])^(a[111] & b[64])^(a[110] & b[65])^(a[109] & b[66])^(a[108] & b[67])^(a[107] & b[68])^(a[106] & b[69])^(a[105] & b[70])^(a[104] & b[71])^(a[103] & b[72])^(a[102] & b[73])^(a[101] & b[74])^(a[100] & b[75])^(a[99] & b[76])^(a[98] & b[77])^(a[97] & b[78])^(a[96] & b[79])^(a[95] & b[80])^(a[94] & b[81])^(a[93] & b[82])^(a[92] & b[83])^(a[91] & b[84])^(a[90] & b[85])^(a[89] & b[86])^(a[88] & b[87])^(a[87] & b[88])^(a[86] & b[89])^(a[85] & b[90])^(a[84] & b[91])^(a[83] & b[92])^(a[82] & b[93])^(a[81] & b[94])^(a[80] & b[95])^(a[79] & b[96])^(a[78] & b[97])^(a[77] & b[98])^(a[76] & b[99])^(a[75] & b[100])^(a[74] & b[101])^(a[73] & b[102])^(a[72] & b[103])^(a[71] & b[104])^(a[70] & b[105])^(a[69] & b[106])^(a[68] & b[107])^(a[67] & b[108])^(a[66] & b[109])^(a[65] & b[110])^(a[64] & b[111])^(a[63] & b[112])^(a[62] & b[113])^(a[61] & b[114])^(a[60] & b[115])^(a[59] & b[116])^(a[58] & b[117])^(a[57] & b[118])^(a[56] & b[119])^(a[55] & b[120])^(a[54] & b[121])^(a[53] & b[122])^(a[52] & b[123])^(a[51] & b[124])^(a[50] & b[125])^(a[49] & b[126])^(a[48] & b[127])^(a[47] & b[128])^(a[46] & b[129])^(a[45] & b[130])^(a[44] & b[131])^(a[43] & b[132])^(a[42] & b[133])^(a[41] & b[134])^(a[40] & b[135])^(a[39] & b[136])^(a[38] & b[137])^(a[37] & b[138])^(a[36] & b[139])^(a[35] & b[140])^(a[34] & b[141])^(a[33] & b[142])^(a[32] & b[143])^(a[31] & b[144])^(a[30] & b[145])^(a[29] & b[146])^(a[28] & b[147])^(a[27] & b[148])^(a[26] & b[149])^(a[25] & b[150])^(a[24] & b[151])^(a[23] & b[152])^(a[22] & b[153])^(a[21] & b[154])^(a[20] & b[155])^(a[19] & b[156])^(a[18] & b[157])^(a[17] & b[158])^(a[16] & b[159])^(a[15] & b[160])^(a[14] & b[161])^(a[13] & b[162]);
assign y[176] = (a[162] & b[14])^(a[161] & b[15])^(a[160] & b[16])^(a[159] & b[17])^(a[158] & b[18])^(a[157] & b[19])^(a[156] & b[20])^(a[155] & b[21])^(a[154] & b[22])^(a[153] & b[23])^(a[152] & b[24])^(a[151] & b[25])^(a[150] & b[26])^(a[149] & b[27])^(a[148] & b[28])^(a[147] & b[29])^(a[146] & b[30])^(a[145] & b[31])^(a[144] & b[32])^(a[143] & b[33])^(a[142] & b[34])^(a[141] & b[35])^(a[140] & b[36])^(a[139] & b[37])^(a[138] & b[38])^(a[137] & b[39])^(a[136] & b[40])^(a[135] & b[41])^(a[134] & b[42])^(a[133] & b[43])^(a[132] & b[44])^(a[131] & b[45])^(a[130] & b[46])^(a[129] & b[47])^(a[128] & b[48])^(a[127] & b[49])^(a[126] & b[50])^(a[125] & b[51])^(a[124] & b[52])^(a[123] & b[53])^(a[122] & b[54])^(a[121] & b[55])^(a[120] & b[56])^(a[119] & b[57])^(a[118] & b[58])^(a[117] & b[59])^(a[116] & b[60])^(a[115] & b[61])^(a[114] & b[62])^(a[113] & b[63])^(a[112] & b[64])^(a[111] & b[65])^(a[110] & b[66])^(a[109] & b[67])^(a[108] & b[68])^(a[107] & b[69])^(a[106] & b[70])^(a[105] & b[71])^(a[104] & b[72])^(a[103] & b[73])^(a[102] & b[74])^(a[101] & b[75])^(a[100] & b[76])^(a[99] & b[77])^(a[98] & b[78])^(a[97] & b[79])^(a[96] & b[80])^(a[95] & b[81])^(a[94] & b[82])^(a[93] & b[83])^(a[92] & b[84])^(a[91] & b[85])^(a[90] & b[86])^(a[89] & b[87])^(a[88] & b[88])^(a[87] & b[89])^(a[86] & b[90])^(a[85] & b[91])^(a[84] & b[92])^(a[83] & b[93])^(a[82] & b[94])^(a[81] & b[95])^(a[80] & b[96])^(a[79] & b[97])^(a[78] & b[98])^(a[77] & b[99])^(a[76] & b[100])^(a[75] & b[101])^(a[74] & b[102])^(a[73] & b[103])^(a[72] & b[104])^(a[71] & b[105])^(a[70] & b[106])^(a[69] & b[107])^(a[68] & b[108])^(a[67] & b[109])^(a[66] & b[110])^(a[65] & b[111])^(a[64] & b[112])^(a[63] & b[113])^(a[62] & b[114])^(a[61] & b[115])^(a[60] & b[116])^(a[59] & b[117])^(a[58] & b[118])^(a[57] & b[119])^(a[56] & b[120])^(a[55] & b[121])^(a[54] & b[122])^(a[53] & b[123])^(a[52] & b[124])^(a[51] & b[125])^(a[50] & b[126])^(a[49] & b[127])^(a[48] & b[128])^(a[47] & b[129])^(a[46] & b[130])^(a[45] & b[131])^(a[44] & b[132])^(a[43] & b[133])^(a[42] & b[134])^(a[41] & b[135])^(a[40] & b[136])^(a[39] & b[137])^(a[38] & b[138])^(a[37] & b[139])^(a[36] & b[140])^(a[35] & b[141])^(a[34] & b[142])^(a[33] & b[143])^(a[32] & b[144])^(a[31] & b[145])^(a[30] & b[146])^(a[29] & b[147])^(a[28] & b[148])^(a[27] & b[149])^(a[26] & b[150])^(a[25] & b[151])^(a[24] & b[152])^(a[23] & b[153])^(a[22] & b[154])^(a[21] & b[155])^(a[20] & b[156])^(a[19] & b[157])^(a[18] & b[158])^(a[17] & b[159])^(a[16] & b[160])^(a[15] & b[161])^(a[14] & b[162]);
assign y[177] = (a[162] & b[15])^(a[161] & b[16])^(a[160] & b[17])^(a[159] & b[18])^(a[158] & b[19])^(a[157] & b[20])^(a[156] & b[21])^(a[155] & b[22])^(a[154] & b[23])^(a[153] & b[24])^(a[152] & b[25])^(a[151] & b[26])^(a[150] & b[27])^(a[149] & b[28])^(a[148] & b[29])^(a[147] & b[30])^(a[146] & b[31])^(a[145] & b[32])^(a[144] & b[33])^(a[143] & b[34])^(a[142] & b[35])^(a[141] & b[36])^(a[140] & b[37])^(a[139] & b[38])^(a[138] & b[39])^(a[137] & b[40])^(a[136] & b[41])^(a[135] & b[42])^(a[134] & b[43])^(a[133] & b[44])^(a[132] & b[45])^(a[131] & b[46])^(a[130] & b[47])^(a[129] & b[48])^(a[128] & b[49])^(a[127] & b[50])^(a[126] & b[51])^(a[125] & b[52])^(a[124] & b[53])^(a[123] & b[54])^(a[122] & b[55])^(a[121] & b[56])^(a[120] & b[57])^(a[119] & b[58])^(a[118] & b[59])^(a[117] & b[60])^(a[116] & b[61])^(a[115] & b[62])^(a[114] & b[63])^(a[113] & b[64])^(a[112] & b[65])^(a[111] & b[66])^(a[110] & b[67])^(a[109] & b[68])^(a[108] & b[69])^(a[107] & b[70])^(a[106] & b[71])^(a[105] & b[72])^(a[104] & b[73])^(a[103] & b[74])^(a[102] & b[75])^(a[101] & b[76])^(a[100] & b[77])^(a[99] & b[78])^(a[98] & b[79])^(a[97] & b[80])^(a[96] & b[81])^(a[95] & b[82])^(a[94] & b[83])^(a[93] & b[84])^(a[92] & b[85])^(a[91] & b[86])^(a[90] & b[87])^(a[89] & b[88])^(a[88] & b[89])^(a[87] & b[90])^(a[86] & b[91])^(a[85] & b[92])^(a[84] & b[93])^(a[83] & b[94])^(a[82] & b[95])^(a[81] & b[96])^(a[80] & b[97])^(a[79] & b[98])^(a[78] & b[99])^(a[77] & b[100])^(a[76] & b[101])^(a[75] & b[102])^(a[74] & b[103])^(a[73] & b[104])^(a[72] & b[105])^(a[71] & b[106])^(a[70] & b[107])^(a[69] & b[108])^(a[68] & b[109])^(a[67] & b[110])^(a[66] & b[111])^(a[65] & b[112])^(a[64] & b[113])^(a[63] & b[114])^(a[62] & b[115])^(a[61] & b[116])^(a[60] & b[117])^(a[59] & b[118])^(a[58] & b[119])^(a[57] & b[120])^(a[56] & b[121])^(a[55] & b[122])^(a[54] & b[123])^(a[53] & b[124])^(a[52] & b[125])^(a[51] & b[126])^(a[50] & b[127])^(a[49] & b[128])^(a[48] & b[129])^(a[47] & b[130])^(a[46] & b[131])^(a[45] & b[132])^(a[44] & b[133])^(a[43] & b[134])^(a[42] & b[135])^(a[41] & b[136])^(a[40] & b[137])^(a[39] & b[138])^(a[38] & b[139])^(a[37] & b[140])^(a[36] & b[141])^(a[35] & b[142])^(a[34] & b[143])^(a[33] & b[144])^(a[32] & b[145])^(a[31] & b[146])^(a[30] & b[147])^(a[29] & b[148])^(a[28] & b[149])^(a[27] & b[150])^(a[26] & b[151])^(a[25] & b[152])^(a[24] & b[153])^(a[23] & b[154])^(a[22] & b[155])^(a[21] & b[156])^(a[20] & b[157])^(a[19] & b[158])^(a[18] & b[159])^(a[17] & b[160])^(a[16] & b[161])^(a[15] & b[162]);
assign y[178] = (a[162] & b[16])^(a[161] & b[17])^(a[160] & b[18])^(a[159] & b[19])^(a[158] & b[20])^(a[157] & b[21])^(a[156] & b[22])^(a[155] & b[23])^(a[154] & b[24])^(a[153] & b[25])^(a[152] & b[26])^(a[151] & b[27])^(a[150] & b[28])^(a[149] & b[29])^(a[148] & b[30])^(a[147] & b[31])^(a[146] & b[32])^(a[145] & b[33])^(a[144] & b[34])^(a[143] & b[35])^(a[142] & b[36])^(a[141] & b[37])^(a[140] & b[38])^(a[139] & b[39])^(a[138] & b[40])^(a[137] & b[41])^(a[136] & b[42])^(a[135] & b[43])^(a[134] & b[44])^(a[133] & b[45])^(a[132] & b[46])^(a[131] & b[47])^(a[130] & b[48])^(a[129] & b[49])^(a[128] & b[50])^(a[127] & b[51])^(a[126] & b[52])^(a[125] & b[53])^(a[124] & b[54])^(a[123] & b[55])^(a[122] & b[56])^(a[121] & b[57])^(a[120] & b[58])^(a[119] & b[59])^(a[118] & b[60])^(a[117] & b[61])^(a[116] & b[62])^(a[115] & b[63])^(a[114] & b[64])^(a[113] & b[65])^(a[112] & b[66])^(a[111] & b[67])^(a[110] & b[68])^(a[109] & b[69])^(a[108] & b[70])^(a[107] & b[71])^(a[106] & b[72])^(a[105] & b[73])^(a[104] & b[74])^(a[103] & b[75])^(a[102] & b[76])^(a[101] & b[77])^(a[100] & b[78])^(a[99] & b[79])^(a[98] & b[80])^(a[97] & b[81])^(a[96] & b[82])^(a[95] & b[83])^(a[94] & b[84])^(a[93] & b[85])^(a[92] & b[86])^(a[91] & b[87])^(a[90] & b[88])^(a[89] & b[89])^(a[88] & b[90])^(a[87] & b[91])^(a[86] & b[92])^(a[85] & b[93])^(a[84] & b[94])^(a[83] & b[95])^(a[82] & b[96])^(a[81] & b[97])^(a[80] & b[98])^(a[79] & b[99])^(a[78] & b[100])^(a[77] & b[101])^(a[76] & b[102])^(a[75] & b[103])^(a[74] & b[104])^(a[73] & b[105])^(a[72] & b[106])^(a[71] & b[107])^(a[70] & b[108])^(a[69] & b[109])^(a[68] & b[110])^(a[67] & b[111])^(a[66] & b[112])^(a[65] & b[113])^(a[64] & b[114])^(a[63] & b[115])^(a[62] & b[116])^(a[61] & b[117])^(a[60] & b[118])^(a[59] & b[119])^(a[58] & b[120])^(a[57] & b[121])^(a[56] & b[122])^(a[55] & b[123])^(a[54] & b[124])^(a[53] & b[125])^(a[52] & b[126])^(a[51] & b[127])^(a[50] & b[128])^(a[49] & b[129])^(a[48] & b[130])^(a[47] & b[131])^(a[46] & b[132])^(a[45] & b[133])^(a[44] & b[134])^(a[43] & b[135])^(a[42] & b[136])^(a[41] & b[137])^(a[40] & b[138])^(a[39] & b[139])^(a[38] & b[140])^(a[37] & b[141])^(a[36] & b[142])^(a[35] & b[143])^(a[34] & b[144])^(a[33] & b[145])^(a[32] & b[146])^(a[31] & b[147])^(a[30] & b[148])^(a[29] & b[149])^(a[28] & b[150])^(a[27] & b[151])^(a[26] & b[152])^(a[25] & b[153])^(a[24] & b[154])^(a[23] & b[155])^(a[22] & b[156])^(a[21] & b[157])^(a[20] & b[158])^(a[19] & b[159])^(a[18] & b[160])^(a[17] & b[161])^(a[16] & b[162]);
assign y[179] = (a[162] & b[17])^(a[161] & b[18])^(a[160] & b[19])^(a[159] & b[20])^(a[158] & b[21])^(a[157] & b[22])^(a[156] & b[23])^(a[155] & b[24])^(a[154] & b[25])^(a[153] & b[26])^(a[152] & b[27])^(a[151] & b[28])^(a[150] & b[29])^(a[149] & b[30])^(a[148] & b[31])^(a[147] & b[32])^(a[146] & b[33])^(a[145] & b[34])^(a[144] & b[35])^(a[143] & b[36])^(a[142] & b[37])^(a[141] & b[38])^(a[140] & b[39])^(a[139] & b[40])^(a[138] & b[41])^(a[137] & b[42])^(a[136] & b[43])^(a[135] & b[44])^(a[134] & b[45])^(a[133] & b[46])^(a[132] & b[47])^(a[131] & b[48])^(a[130] & b[49])^(a[129] & b[50])^(a[128] & b[51])^(a[127] & b[52])^(a[126] & b[53])^(a[125] & b[54])^(a[124] & b[55])^(a[123] & b[56])^(a[122] & b[57])^(a[121] & b[58])^(a[120] & b[59])^(a[119] & b[60])^(a[118] & b[61])^(a[117] & b[62])^(a[116] & b[63])^(a[115] & b[64])^(a[114] & b[65])^(a[113] & b[66])^(a[112] & b[67])^(a[111] & b[68])^(a[110] & b[69])^(a[109] & b[70])^(a[108] & b[71])^(a[107] & b[72])^(a[106] & b[73])^(a[105] & b[74])^(a[104] & b[75])^(a[103] & b[76])^(a[102] & b[77])^(a[101] & b[78])^(a[100] & b[79])^(a[99] & b[80])^(a[98] & b[81])^(a[97] & b[82])^(a[96] & b[83])^(a[95] & b[84])^(a[94] & b[85])^(a[93] & b[86])^(a[92] & b[87])^(a[91] & b[88])^(a[90] & b[89])^(a[89] & b[90])^(a[88] & b[91])^(a[87] & b[92])^(a[86] & b[93])^(a[85] & b[94])^(a[84] & b[95])^(a[83] & b[96])^(a[82] & b[97])^(a[81] & b[98])^(a[80] & b[99])^(a[79] & b[100])^(a[78] & b[101])^(a[77] & b[102])^(a[76] & b[103])^(a[75] & b[104])^(a[74] & b[105])^(a[73] & b[106])^(a[72] & b[107])^(a[71] & b[108])^(a[70] & b[109])^(a[69] & b[110])^(a[68] & b[111])^(a[67] & b[112])^(a[66] & b[113])^(a[65] & b[114])^(a[64] & b[115])^(a[63] & b[116])^(a[62] & b[117])^(a[61] & b[118])^(a[60] & b[119])^(a[59] & b[120])^(a[58] & b[121])^(a[57] & b[122])^(a[56] & b[123])^(a[55] & b[124])^(a[54] & b[125])^(a[53] & b[126])^(a[52] & b[127])^(a[51] & b[128])^(a[50] & b[129])^(a[49] & b[130])^(a[48] & b[131])^(a[47] & b[132])^(a[46] & b[133])^(a[45] & b[134])^(a[44] & b[135])^(a[43] & b[136])^(a[42] & b[137])^(a[41] & b[138])^(a[40] & b[139])^(a[39] & b[140])^(a[38] & b[141])^(a[37] & b[142])^(a[36] & b[143])^(a[35] & b[144])^(a[34] & b[145])^(a[33] & b[146])^(a[32] & b[147])^(a[31] & b[148])^(a[30] & b[149])^(a[29] & b[150])^(a[28] & b[151])^(a[27] & b[152])^(a[26] & b[153])^(a[25] & b[154])^(a[24] & b[155])^(a[23] & b[156])^(a[22] & b[157])^(a[21] & b[158])^(a[20] & b[159])^(a[19] & b[160])^(a[18] & b[161])^(a[17] & b[162]);
assign y[180] = (a[162] & b[18])^(a[161] & b[19])^(a[160] & b[20])^(a[159] & b[21])^(a[158] & b[22])^(a[157] & b[23])^(a[156] & b[24])^(a[155] & b[25])^(a[154] & b[26])^(a[153] & b[27])^(a[152] & b[28])^(a[151] & b[29])^(a[150] & b[30])^(a[149] & b[31])^(a[148] & b[32])^(a[147] & b[33])^(a[146] & b[34])^(a[145] & b[35])^(a[144] & b[36])^(a[143] & b[37])^(a[142] & b[38])^(a[141] & b[39])^(a[140] & b[40])^(a[139] & b[41])^(a[138] & b[42])^(a[137] & b[43])^(a[136] & b[44])^(a[135] & b[45])^(a[134] & b[46])^(a[133] & b[47])^(a[132] & b[48])^(a[131] & b[49])^(a[130] & b[50])^(a[129] & b[51])^(a[128] & b[52])^(a[127] & b[53])^(a[126] & b[54])^(a[125] & b[55])^(a[124] & b[56])^(a[123] & b[57])^(a[122] & b[58])^(a[121] & b[59])^(a[120] & b[60])^(a[119] & b[61])^(a[118] & b[62])^(a[117] & b[63])^(a[116] & b[64])^(a[115] & b[65])^(a[114] & b[66])^(a[113] & b[67])^(a[112] & b[68])^(a[111] & b[69])^(a[110] & b[70])^(a[109] & b[71])^(a[108] & b[72])^(a[107] & b[73])^(a[106] & b[74])^(a[105] & b[75])^(a[104] & b[76])^(a[103] & b[77])^(a[102] & b[78])^(a[101] & b[79])^(a[100] & b[80])^(a[99] & b[81])^(a[98] & b[82])^(a[97] & b[83])^(a[96] & b[84])^(a[95] & b[85])^(a[94] & b[86])^(a[93] & b[87])^(a[92] & b[88])^(a[91] & b[89])^(a[90] & b[90])^(a[89] & b[91])^(a[88] & b[92])^(a[87] & b[93])^(a[86] & b[94])^(a[85] & b[95])^(a[84] & b[96])^(a[83] & b[97])^(a[82] & b[98])^(a[81] & b[99])^(a[80] & b[100])^(a[79] & b[101])^(a[78] & b[102])^(a[77] & b[103])^(a[76] & b[104])^(a[75] & b[105])^(a[74] & b[106])^(a[73] & b[107])^(a[72] & b[108])^(a[71] & b[109])^(a[70] & b[110])^(a[69] & b[111])^(a[68] & b[112])^(a[67] & b[113])^(a[66] & b[114])^(a[65] & b[115])^(a[64] & b[116])^(a[63] & b[117])^(a[62] & b[118])^(a[61] & b[119])^(a[60] & b[120])^(a[59] & b[121])^(a[58] & b[122])^(a[57] & b[123])^(a[56] & b[124])^(a[55] & b[125])^(a[54] & b[126])^(a[53] & b[127])^(a[52] & b[128])^(a[51] & b[129])^(a[50] & b[130])^(a[49] & b[131])^(a[48] & b[132])^(a[47] & b[133])^(a[46] & b[134])^(a[45] & b[135])^(a[44] & b[136])^(a[43] & b[137])^(a[42] & b[138])^(a[41] & b[139])^(a[40] & b[140])^(a[39] & b[141])^(a[38] & b[142])^(a[37] & b[143])^(a[36] & b[144])^(a[35] & b[145])^(a[34] & b[146])^(a[33] & b[147])^(a[32] & b[148])^(a[31] & b[149])^(a[30] & b[150])^(a[29] & b[151])^(a[28] & b[152])^(a[27] & b[153])^(a[26] & b[154])^(a[25] & b[155])^(a[24] & b[156])^(a[23] & b[157])^(a[22] & b[158])^(a[21] & b[159])^(a[20] & b[160])^(a[19] & b[161])^(a[18] & b[162]);
assign y[181] = (a[162] & b[19])^(a[161] & b[20])^(a[160] & b[21])^(a[159] & b[22])^(a[158] & b[23])^(a[157] & b[24])^(a[156] & b[25])^(a[155] & b[26])^(a[154] & b[27])^(a[153] & b[28])^(a[152] & b[29])^(a[151] & b[30])^(a[150] & b[31])^(a[149] & b[32])^(a[148] & b[33])^(a[147] & b[34])^(a[146] & b[35])^(a[145] & b[36])^(a[144] & b[37])^(a[143] & b[38])^(a[142] & b[39])^(a[141] & b[40])^(a[140] & b[41])^(a[139] & b[42])^(a[138] & b[43])^(a[137] & b[44])^(a[136] & b[45])^(a[135] & b[46])^(a[134] & b[47])^(a[133] & b[48])^(a[132] & b[49])^(a[131] & b[50])^(a[130] & b[51])^(a[129] & b[52])^(a[128] & b[53])^(a[127] & b[54])^(a[126] & b[55])^(a[125] & b[56])^(a[124] & b[57])^(a[123] & b[58])^(a[122] & b[59])^(a[121] & b[60])^(a[120] & b[61])^(a[119] & b[62])^(a[118] & b[63])^(a[117] & b[64])^(a[116] & b[65])^(a[115] & b[66])^(a[114] & b[67])^(a[113] & b[68])^(a[112] & b[69])^(a[111] & b[70])^(a[110] & b[71])^(a[109] & b[72])^(a[108] & b[73])^(a[107] & b[74])^(a[106] & b[75])^(a[105] & b[76])^(a[104] & b[77])^(a[103] & b[78])^(a[102] & b[79])^(a[101] & b[80])^(a[100] & b[81])^(a[99] & b[82])^(a[98] & b[83])^(a[97] & b[84])^(a[96] & b[85])^(a[95] & b[86])^(a[94] & b[87])^(a[93] & b[88])^(a[92] & b[89])^(a[91] & b[90])^(a[90] & b[91])^(a[89] & b[92])^(a[88] & b[93])^(a[87] & b[94])^(a[86] & b[95])^(a[85] & b[96])^(a[84] & b[97])^(a[83] & b[98])^(a[82] & b[99])^(a[81] & b[100])^(a[80] & b[101])^(a[79] & b[102])^(a[78] & b[103])^(a[77] & b[104])^(a[76] & b[105])^(a[75] & b[106])^(a[74] & b[107])^(a[73] & b[108])^(a[72] & b[109])^(a[71] & b[110])^(a[70] & b[111])^(a[69] & b[112])^(a[68] & b[113])^(a[67] & b[114])^(a[66] & b[115])^(a[65] & b[116])^(a[64] & b[117])^(a[63] & b[118])^(a[62] & b[119])^(a[61] & b[120])^(a[60] & b[121])^(a[59] & b[122])^(a[58] & b[123])^(a[57] & b[124])^(a[56] & b[125])^(a[55] & b[126])^(a[54] & b[127])^(a[53] & b[128])^(a[52] & b[129])^(a[51] & b[130])^(a[50] & b[131])^(a[49] & b[132])^(a[48] & b[133])^(a[47] & b[134])^(a[46] & b[135])^(a[45] & b[136])^(a[44] & b[137])^(a[43] & b[138])^(a[42] & b[139])^(a[41] & b[140])^(a[40] & b[141])^(a[39] & b[142])^(a[38] & b[143])^(a[37] & b[144])^(a[36] & b[145])^(a[35] & b[146])^(a[34] & b[147])^(a[33] & b[148])^(a[32] & b[149])^(a[31] & b[150])^(a[30] & b[151])^(a[29] & b[152])^(a[28] & b[153])^(a[27] & b[154])^(a[26] & b[155])^(a[25] & b[156])^(a[24] & b[157])^(a[23] & b[158])^(a[22] & b[159])^(a[21] & b[160])^(a[20] & b[161])^(a[19] & b[162]);
assign y[182] = (a[162] & b[20])^(a[161] & b[21])^(a[160] & b[22])^(a[159] & b[23])^(a[158] & b[24])^(a[157] & b[25])^(a[156] & b[26])^(a[155] & b[27])^(a[154] & b[28])^(a[153] & b[29])^(a[152] & b[30])^(a[151] & b[31])^(a[150] & b[32])^(a[149] & b[33])^(a[148] & b[34])^(a[147] & b[35])^(a[146] & b[36])^(a[145] & b[37])^(a[144] & b[38])^(a[143] & b[39])^(a[142] & b[40])^(a[141] & b[41])^(a[140] & b[42])^(a[139] & b[43])^(a[138] & b[44])^(a[137] & b[45])^(a[136] & b[46])^(a[135] & b[47])^(a[134] & b[48])^(a[133] & b[49])^(a[132] & b[50])^(a[131] & b[51])^(a[130] & b[52])^(a[129] & b[53])^(a[128] & b[54])^(a[127] & b[55])^(a[126] & b[56])^(a[125] & b[57])^(a[124] & b[58])^(a[123] & b[59])^(a[122] & b[60])^(a[121] & b[61])^(a[120] & b[62])^(a[119] & b[63])^(a[118] & b[64])^(a[117] & b[65])^(a[116] & b[66])^(a[115] & b[67])^(a[114] & b[68])^(a[113] & b[69])^(a[112] & b[70])^(a[111] & b[71])^(a[110] & b[72])^(a[109] & b[73])^(a[108] & b[74])^(a[107] & b[75])^(a[106] & b[76])^(a[105] & b[77])^(a[104] & b[78])^(a[103] & b[79])^(a[102] & b[80])^(a[101] & b[81])^(a[100] & b[82])^(a[99] & b[83])^(a[98] & b[84])^(a[97] & b[85])^(a[96] & b[86])^(a[95] & b[87])^(a[94] & b[88])^(a[93] & b[89])^(a[92] & b[90])^(a[91] & b[91])^(a[90] & b[92])^(a[89] & b[93])^(a[88] & b[94])^(a[87] & b[95])^(a[86] & b[96])^(a[85] & b[97])^(a[84] & b[98])^(a[83] & b[99])^(a[82] & b[100])^(a[81] & b[101])^(a[80] & b[102])^(a[79] & b[103])^(a[78] & b[104])^(a[77] & b[105])^(a[76] & b[106])^(a[75] & b[107])^(a[74] & b[108])^(a[73] & b[109])^(a[72] & b[110])^(a[71] & b[111])^(a[70] & b[112])^(a[69] & b[113])^(a[68] & b[114])^(a[67] & b[115])^(a[66] & b[116])^(a[65] & b[117])^(a[64] & b[118])^(a[63] & b[119])^(a[62] & b[120])^(a[61] & b[121])^(a[60] & b[122])^(a[59] & b[123])^(a[58] & b[124])^(a[57] & b[125])^(a[56] & b[126])^(a[55] & b[127])^(a[54] & b[128])^(a[53] & b[129])^(a[52] & b[130])^(a[51] & b[131])^(a[50] & b[132])^(a[49] & b[133])^(a[48] & b[134])^(a[47] & b[135])^(a[46] & b[136])^(a[45] & b[137])^(a[44] & b[138])^(a[43] & b[139])^(a[42] & b[140])^(a[41] & b[141])^(a[40] & b[142])^(a[39] & b[143])^(a[38] & b[144])^(a[37] & b[145])^(a[36] & b[146])^(a[35] & b[147])^(a[34] & b[148])^(a[33] & b[149])^(a[32] & b[150])^(a[31] & b[151])^(a[30] & b[152])^(a[29] & b[153])^(a[28] & b[154])^(a[27] & b[155])^(a[26] & b[156])^(a[25] & b[157])^(a[24] & b[158])^(a[23] & b[159])^(a[22] & b[160])^(a[21] & b[161])^(a[20] & b[162]);
assign y[183] = (a[162] & b[21])^(a[161] & b[22])^(a[160] & b[23])^(a[159] & b[24])^(a[158] & b[25])^(a[157] & b[26])^(a[156] & b[27])^(a[155] & b[28])^(a[154] & b[29])^(a[153] & b[30])^(a[152] & b[31])^(a[151] & b[32])^(a[150] & b[33])^(a[149] & b[34])^(a[148] & b[35])^(a[147] & b[36])^(a[146] & b[37])^(a[145] & b[38])^(a[144] & b[39])^(a[143] & b[40])^(a[142] & b[41])^(a[141] & b[42])^(a[140] & b[43])^(a[139] & b[44])^(a[138] & b[45])^(a[137] & b[46])^(a[136] & b[47])^(a[135] & b[48])^(a[134] & b[49])^(a[133] & b[50])^(a[132] & b[51])^(a[131] & b[52])^(a[130] & b[53])^(a[129] & b[54])^(a[128] & b[55])^(a[127] & b[56])^(a[126] & b[57])^(a[125] & b[58])^(a[124] & b[59])^(a[123] & b[60])^(a[122] & b[61])^(a[121] & b[62])^(a[120] & b[63])^(a[119] & b[64])^(a[118] & b[65])^(a[117] & b[66])^(a[116] & b[67])^(a[115] & b[68])^(a[114] & b[69])^(a[113] & b[70])^(a[112] & b[71])^(a[111] & b[72])^(a[110] & b[73])^(a[109] & b[74])^(a[108] & b[75])^(a[107] & b[76])^(a[106] & b[77])^(a[105] & b[78])^(a[104] & b[79])^(a[103] & b[80])^(a[102] & b[81])^(a[101] & b[82])^(a[100] & b[83])^(a[99] & b[84])^(a[98] & b[85])^(a[97] & b[86])^(a[96] & b[87])^(a[95] & b[88])^(a[94] & b[89])^(a[93] & b[90])^(a[92] & b[91])^(a[91] & b[92])^(a[90] & b[93])^(a[89] & b[94])^(a[88] & b[95])^(a[87] & b[96])^(a[86] & b[97])^(a[85] & b[98])^(a[84] & b[99])^(a[83] & b[100])^(a[82] & b[101])^(a[81] & b[102])^(a[80] & b[103])^(a[79] & b[104])^(a[78] & b[105])^(a[77] & b[106])^(a[76] & b[107])^(a[75] & b[108])^(a[74] & b[109])^(a[73] & b[110])^(a[72] & b[111])^(a[71] & b[112])^(a[70] & b[113])^(a[69] & b[114])^(a[68] & b[115])^(a[67] & b[116])^(a[66] & b[117])^(a[65] & b[118])^(a[64] & b[119])^(a[63] & b[120])^(a[62] & b[121])^(a[61] & b[122])^(a[60] & b[123])^(a[59] & b[124])^(a[58] & b[125])^(a[57] & b[126])^(a[56] & b[127])^(a[55] & b[128])^(a[54] & b[129])^(a[53] & b[130])^(a[52] & b[131])^(a[51] & b[132])^(a[50] & b[133])^(a[49] & b[134])^(a[48] & b[135])^(a[47] & b[136])^(a[46] & b[137])^(a[45] & b[138])^(a[44] & b[139])^(a[43] & b[140])^(a[42] & b[141])^(a[41] & b[142])^(a[40] & b[143])^(a[39] & b[144])^(a[38] & b[145])^(a[37] & b[146])^(a[36] & b[147])^(a[35] & b[148])^(a[34] & b[149])^(a[33] & b[150])^(a[32] & b[151])^(a[31] & b[152])^(a[30] & b[153])^(a[29] & b[154])^(a[28] & b[155])^(a[27] & b[156])^(a[26] & b[157])^(a[25] & b[158])^(a[24] & b[159])^(a[23] & b[160])^(a[22] & b[161])^(a[21] & b[162]);
assign y[184] = (a[162] & b[22])^(a[161] & b[23])^(a[160] & b[24])^(a[159] & b[25])^(a[158] & b[26])^(a[157] & b[27])^(a[156] & b[28])^(a[155] & b[29])^(a[154] & b[30])^(a[153] & b[31])^(a[152] & b[32])^(a[151] & b[33])^(a[150] & b[34])^(a[149] & b[35])^(a[148] & b[36])^(a[147] & b[37])^(a[146] & b[38])^(a[145] & b[39])^(a[144] & b[40])^(a[143] & b[41])^(a[142] & b[42])^(a[141] & b[43])^(a[140] & b[44])^(a[139] & b[45])^(a[138] & b[46])^(a[137] & b[47])^(a[136] & b[48])^(a[135] & b[49])^(a[134] & b[50])^(a[133] & b[51])^(a[132] & b[52])^(a[131] & b[53])^(a[130] & b[54])^(a[129] & b[55])^(a[128] & b[56])^(a[127] & b[57])^(a[126] & b[58])^(a[125] & b[59])^(a[124] & b[60])^(a[123] & b[61])^(a[122] & b[62])^(a[121] & b[63])^(a[120] & b[64])^(a[119] & b[65])^(a[118] & b[66])^(a[117] & b[67])^(a[116] & b[68])^(a[115] & b[69])^(a[114] & b[70])^(a[113] & b[71])^(a[112] & b[72])^(a[111] & b[73])^(a[110] & b[74])^(a[109] & b[75])^(a[108] & b[76])^(a[107] & b[77])^(a[106] & b[78])^(a[105] & b[79])^(a[104] & b[80])^(a[103] & b[81])^(a[102] & b[82])^(a[101] & b[83])^(a[100] & b[84])^(a[99] & b[85])^(a[98] & b[86])^(a[97] & b[87])^(a[96] & b[88])^(a[95] & b[89])^(a[94] & b[90])^(a[93] & b[91])^(a[92] & b[92])^(a[91] & b[93])^(a[90] & b[94])^(a[89] & b[95])^(a[88] & b[96])^(a[87] & b[97])^(a[86] & b[98])^(a[85] & b[99])^(a[84] & b[100])^(a[83] & b[101])^(a[82] & b[102])^(a[81] & b[103])^(a[80] & b[104])^(a[79] & b[105])^(a[78] & b[106])^(a[77] & b[107])^(a[76] & b[108])^(a[75] & b[109])^(a[74] & b[110])^(a[73] & b[111])^(a[72] & b[112])^(a[71] & b[113])^(a[70] & b[114])^(a[69] & b[115])^(a[68] & b[116])^(a[67] & b[117])^(a[66] & b[118])^(a[65] & b[119])^(a[64] & b[120])^(a[63] & b[121])^(a[62] & b[122])^(a[61] & b[123])^(a[60] & b[124])^(a[59] & b[125])^(a[58] & b[126])^(a[57] & b[127])^(a[56] & b[128])^(a[55] & b[129])^(a[54] & b[130])^(a[53] & b[131])^(a[52] & b[132])^(a[51] & b[133])^(a[50] & b[134])^(a[49] & b[135])^(a[48] & b[136])^(a[47] & b[137])^(a[46] & b[138])^(a[45] & b[139])^(a[44] & b[140])^(a[43] & b[141])^(a[42] & b[142])^(a[41] & b[143])^(a[40] & b[144])^(a[39] & b[145])^(a[38] & b[146])^(a[37] & b[147])^(a[36] & b[148])^(a[35] & b[149])^(a[34] & b[150])^(a[33] & b[151])^(a[32] & b[152])^(a[31] & b[153])^(a[30] & b[154])^(a[29] & b[155])^(a[28] & b[156])^(a[27] & b[157])^(a[26] & b[158])^(a[25] & b[159])^(a[24] & b[160])^(a[23] & b[161])^(a[22] & b[162]);
assign y[185] = (a[162] & b[23])^(a[161] & b[24])^(a[160] & b[25])^(a[159] & b[26])^(a[158] & b[27])^(a[157] & b[28])^(a[156] & b[29])^(a[155] & b[30])^(a[154] & b[31])^(a[153] & b[32])^(a[152] & b[33])^(a[151] & b[34])^(a[150] & b[35])^(a[149] & b[36])^(a[148] & b[37])^(a[147] & b[38])^(a[146] & b[39])^(a[145] & b[40])^(a[144] & b[41])^(a[143] & b[42])^(a[142] & b[43])^(a[141] & b[44])^(a[140] & b[45])^(a[139] & b[46])^(a[138] & b[47])^(a[137] & b[48])^(a[136] & b[49])^(a[135] & b[50])^(a[134] & b[51])^(a[133] & b[52])^(a[132] & b[53])^(a[131] & b[54])^(a[130] & b[55])^(a[129] & b[56])^(a[128] & b[57])^(a[127] & b[58])^(a[126] & b[59])^(a[125] & b[60])^(a[124] & b[61])^(a[123] & b[62])^(a[122] & b[63])^(a[121] & b[64])^(a[120] & b[65])^(a[119] & b[66])^(a[118] & b[67])^(a[117] & b[68])^(a[116] & b[69])^(a[115] & b[70])^(a[114] & b[71])^(a[113] & b[72])^(a[112] & b[73])^(a[111] & b[74])^(a[110] & b[75])^(a[109] & b[76])^(a[108] & b[77])^(a[107] & b[78])^(a[106] & b[79])^(a[105] & b[80])^(a[104] & b[81])^(a[103] & b[82])^(a[102] & b[83])^(a[101] & b[84])^(a[100] & b[85])^(a[99] & b[86])^(a[98] & b[87])^(a[97] & b[88])^(a[96] & b[89])^(a[95] & b[90])^(a[94] & b[91])^(a[93] & b[92])^(a[92] & b[93])^(a[91] & b[94])^(a[90] & b[95])^(a[89] & b[96])^(a[88] & b[97])^(a[87] & b[98])^(a[86] & b[99])^(a[85] & b[100])^(a[84] & b[101])^(a[83] & b[102])^(a[82] & b[103])^(a[81] & b[104])^(a[80] & b[105])^(a[79] & b[106])^(a[78] & b[107])^(a[77] & b[108])^(a[76] & b[109])^(a[75] & b[110])^(a[74] & b[111])^(a[73] & b[112])^(a[72] & b[113])^(a[71] & b[114])^(a[70] & b[115])^(a[69] & b[116])^(a[68] & b[117])^(a[67] & b[118])^(a[66] & b[119])^(a[65] & b[120])^(a[64] & b[121])^(a[63] & b[122])^(a[62] & b[123])^(a[61] & b[124])^(a[60] & b[125])^(a[59] & b[126])^(a[58] & b[127])^(a[57] & b[128])^(a[56] & b[129])^(a[55] & b[130])^(a[54] & b[131])^(a[53] & b[132])^(a[52] & b[133])^(a[51] & b[134])^(a[50] & b[135])^(a[49] & b[136])^(a[48] & b[137])^(a[47] & b[138])^(a[46] & b[139])^(a[45] & b[140])^(a[44] & b[141])^(a[43] & b[142])^(a[42] & b[143])^(a[41] & b[144])^(a[40] & b[145])^(a[39] & b[146])^(a[38] & b[147])^(a[37] & b[148])^(a[36] & b[149])^(a[35] & b[150])^(a[34] & b[151])^(a[33] & b[152])^(a[32] & b[153])^(a[31] & b[154])^(a[30] & b[155])^(a[29] & b[156])^(a[28] & b[157])^(a[27] & b[158])^(a[26] & b[159])^(a[25] & b[160])^(a[24] & b[161])^(a[23] & b[162]);
assign y[186] = (a[162] & b[24])^(a[161] & b[25])^(a[160] & b[26])^(a[159] & b[27])^(a[158] & b[28])^(a[157] & b[29])^(a[156] & b[30])^(a[155] & b[31])^(a[154] & b[32])^(a[153] & b[33])^(a[152] & b[34])^(a[151] & b[35])^(a[150] & b[36])^(a[149] & b[37])^(a[148] & b[38])^(a[147] & b[39])^(a[146] & b[40])^(a[145] & b[41])^(a[144] & b[42])^(a[143] & b[43])^(a[142] & b[44])^(a[141] & b[45])^(a[140] & b[46])^(a[139] & b[47])^(a[138] & b[48])^(a[137] & b[49])^(a[136] & b[50])^(a[135] & b[51])^(a[134] & b[52])^(a[133] & b[53])^(a[132] & b[54])^(a[131] & b[55])^(a[130] & b[56])^(a[129] & b[57])^(a[128] & b[58])^(a[127] & b[59])^(a[126] & b[60])^(a[125] & b[61])^(a[124] & b[62])^(a[123] & b[63])^(a[122] & b[64])^(a[121] & b[65])^(a[120] & b[66])^(a[119] & b[67])^(a[118] & b[68])^(a[117] & b[69])^(a[116] & b[70])^(a[115] & b[71])^(a[114] & b[72])^(a[113] & b[73])^(a[112] & b[74])^(a[111] & b[75])^(a[110] & b[76])^(a[109] & b[77])^(a[108] & b[78])^(a[107] & b[79])^(a[106] & b[80])^(a[105] & b[81])^(a[104] & b[82])^(a[103] & b[83])^(a[102] & b[84])^(a[101] & b[85])^(a[100] & b[86])^(a[99] & b[87])^(a[98] & b[88])^(a[97] & b[89])^(a[96] & b[90])^(a[95] & b[91])^(a[94] & b[92])^(a[93] & b[93])^(a[92] & b[94])^(a[91] & b[95])^(a[90] & b[96])^(a[89] & b[97])^(a[88] & b[98])^(a[87] & b[99])^(a[86] & b[100])^(a[85] & b[101])^(a[84] & b[102])^(a[83] & b[103])^(a[82] & b[104])^(a[81] & b[105])^(a[80] & b[106])^(a[79] & b[107])^(a[78] & b[108])^(a[77] & b[109])^(a[76] & b[110])^(a[75] & b[111])^(a[74] & b[112])^(a[73] & b[113])^(a[72] & b[114])^(a[71] & b[115])^(a[70] & b[116])^(a[69] & b[117])^(a[68] & b[118])^(a[67] & b[119])^(a[66] & b[120])^(a[65] & b[121])^(a[64] & b[122])^(a[63] & b[123])^(a[62] & b[124])^(a[61] & b[125])^(a[60] & b[126])^(a[59] & b[127])^(a[58] & b[128])^(a[57] & b[129])^(a[56] & b[130])^(a[55] & b[131])^(a[54] & b[132])^(a[53] & b[133])^(a[52] & b[134])^(a[51] & b[135])^(a[50] & b[136])^(a[49] & b[137])^(a[48] & b[138])^(a[47] & b[139])^(a[46] & b[140])^(a[45] & b[141])^(a[44] & b[142])^(a[43] & b[143])^(a[42] & b[144])^(a[41] & b[145])^(a[40] & b[146])^(a[39] & b[147])^(a[38] & b[148])^(a[37] & b[149])^(a[36] & b[150])^(a[35] & b[151])^(a[34] & b[152])^(a[33] & b[153])^(a[32] & b[154])^(a[31] & b[155])^(a[30] & b[156])^(a[29] & b[157])^(a[28] & b[158])^(a[27] & b[159])^(a[26] & b[160])^(a[25] & b[161])^(a[24] & b[162]);
assign y[187] = (a[162] & b[25])^(a[161] & b[26])^(a[160] & b[27])^(a[159] & b[28])^(a[158] & b[29])^(a[157] & b[30])^(a[156] & b[31])^(a[155] & b[32])^(a[154] & b[33])^(a[153] & b[34])^(a[152] & b[35])^(a[151] & b[36])^(a[150] & b[37])^(a[149] & b[38])^(a[148] & b[39])^(a[147] & b[40])^(a[146] & b[41])^(a[145] & b[42])^(a[144] & b[43])^(a[143] & b[44])^(a[142] & b[45])^(a[141] & b[46])^(a[140] & b[47])^(a[139] & b[48])^(a[138] & b[49])^(a[137] & b[50])^(a[136] & b[51])^(a[135] & b[52])^(a[134] & b[53])^(a[133] & b[54])^(a[132] & b[55])^(a[131] & b[56])^(a[130] & b[57])^(a[129] & b[58])^(a[128] & b[59])^(a[127] & b[60])^(a[126] & b[61])^(a[125] & b[62])^(a[124] & b[63])^(a[123] & b[64])^(a[122] & b[65])^(a[121] & b[66])^(a[120] & b[67])^(a[119] & b[68])^(a[118] & b[69])^(a[117] & b[70])^(a[116] & b[71])^(a[115] & b[72])^(a[114] & b[73])^(a[113] & b[74])^(a[112] & b[75])^(a[111] & b[76])^(a[110] & b[77])^(a[109] & b[78])^(a[108] & b[79])^(a[107] & b[80])^(a[106] & b[81])^(a[105] & b[82])^(a[104] & b[83])^(a[103] & b[84])^(a[102] & b[85])^(a[101] & b[86])^(a[100] & b[87])^(a[99] & b[88])^(a[98] & b[89])^(a[97] & b[90])^(a[96] & b[91])^(a[95] & b[92])^(a[94] & b[93])^(a[93] & b[94])^(a[92] & b[95])^(a[91] & b[96])^(a[90] & b[97])^(a[89] & b[98])^(a[88] & b[99])^(a[87] & b[100])^(a[86] & b[101])^(a[85] & b[102])^(a[84] & b[103])^(a[83] & b[104])^(a[82] & b[105])^(a[81] & b[106])^(a[80] & b[107])^(a[79] & b[108])^(a[78] & b[109])^(a[77] & b[110])^(a[76] & b[111])^(a[75] & b[112])^(a[74] & b[113])^(a[73] & b[114])^(a[72] & b[115])^(a[71] & b[116])^(a[70] & b[117])^(a[69] & b[118])^(a[68] & b[119])^(a[67] & b[120])^(a[66] & b[121])^(a[65] & b[122])^(a[64] & b[123])^(a[63] & b[124])^(a[62] & b[125])^(a[61] & b[126])^(a[60] & b[127])^(a[59] & b[128])^(a[58] & b[129])^(a[57] & b[130])^(a[56] & b[131])^(a[55] & b[132])^(a[54] & b[133])^(a[53] & b[134])^(a[52] & b[135])^(a[51] & b[136])^(a[50] & b[137])^(a[49] & b[138])^(a[48] & b[139])^(a[47] & b[140])^(a[46] & b[141])^(a[45] & b[142])^(a[44] & b[143])^(a[43] & b[144])^(a[42] & b[145])^(a[41] & b[146])^(a[40] & b[147])^(a[39] & b[148])^(a[38] & b[149])^(a[37] & b[150])^(a[36] & b[151])^(a[35] & b[152])^(a[34] & b[153])^(a[33] & b[154])^(a[32] & b[155])^(a[31] & b[156])^(a[30] & b[157])^(a[29] & b[158])^(a[28] & b[159])^(a[27] & b[160])^(a[26] & b[161])^(a[25] & b[162]);
assign y[188] = (a[162] & b[26])^(a[161] & b[27])^(a[160] & b[28])^(a[159] & b[29])^(a[158] & b[30])^(a[157] & b[31])^(a[156] & b[32])^(a[155] & b[33])^(a[154] & b[34])^(a[153] & b[35])^(a[152] & b[36])^(a[151] & b[37])^(a[150] & b[38])^(a[149] & b[39])^(a[148] & b[40])^(a[147] & b[41])^(a[146] & b[42])^(a[145] & b[43])^(a[144] & b[44])^(a[143] & b[45])^(a[142] & b[46])^(a[141] & b[47])^(a[140] & b[48])^(a[139] & b[49])^(a[138] & b[50])^(a[137] & b[51])^(a[136] & b[52])^(a[135] & b[53])^(a[134] & b[54])^(a[133] & b[55])^(a[132] & b[56])^(a[131] & b[57])^(a[130] & b[58])^(a[129] & b[59])^(a[128] & b[60])^(a[127] & b[61])^(a[126] & b[62])^(a[125] & b[63])^(a[124] & b[64])^(a[123] & b[65])^(a[122] & b[66])^(a[121] & b[67])^(a[120] & b[68])^(a[119] & b[69])^(a[118] & b[70])^(a[117] & b[71])^(a[116] & b[72])^(a[115] & b[73])^(a[114] & b[74])^(a[113] & b[75])^(a[112] & b[76])^(a[111] & b[77])^(a[110] & b[78])^(a[109] & b[79])^(a[108] & b[80])^(a[107] & b[81])^(a[106] & b[82])^(a[105] & b[83])^(a[104] & b[84])^(a[103] & b[85])^(a[102] & b[86])^(a[101] & b[87])^(a[100] & b[88])^(a[99] & b[89])^(a[98] & b[90])^(a[97] & b[91])^(a[96] & b[92])^(a[95] & b[93])^(a[94] & b[94])^(a[93] & b[95])^(a[92] & b[96])^(a[91] & b[97])^(a[90] & b[98])^(a[89] & b[99])^(a[88] & b[100])^(a[87] & b[101])^(a[86] & b[102])^(a[85] & b[103])^(a[84] & b[104])^(a[83] & b[105])^(a[82] & b[106])^(a[81] & b[107])^(a[80] & b[108])^(a[79] & b[109])^(a[78] & b[110])^(a[77] & b[111])^(a[76] & b[112])^(a[75] & b[113])^(a[74] & b[114])^(a[73] & b[115])^(a[72] & b[116])^(a[71] & b[117])^(a[70] & b[118])^(a[69] & b[119])^(a[68] & b[120])^(a[67] & b[121])^(a[66] & b[122])^(a[65] & b[123])^(a[64] & b[124])^(a[63] & b[125])^(a[62] & b[126])^(a[61] & b[127])^(a[60] & b[128])^(a[59] & b[129])^(a[58] & b[130])^(a[57] & b[131])^(a[56] & b[132])^(a[55] & b[133])^(a[54] & b[134])^(a[53] & b[135])^(a[52] & b[136])^(a[51] & b[137])^(a[50] & b[138])^(a[49] & b[139])^(a[48] & b[140])^(a[47] & b[141])^(a[46] & b[142])^(a[45] & b[143])^(a[44] & b[144])^(a[43] & b[145])^(a[42] & b[146])^(a[41] & b[147])^(a[40] & b[148])^(a[39] & b[149])^(a[38] & b[150])^(a[37] & b[151])^(a[36] & b[152])^(a[35] & b[153])^(a[34] & b[154])^(a[33] & b[155])^(a[32] & b[156])^(a[31] & b[157])^(a[30] & b[158])^(a[29] & b[159])^(a[28] & b[160])^(a[27] & b[161])^(a[26] & b[162]);
assign y[189] = (a[162] & b[27])^(a[161] & b[28])^(a[160] & b[29])^(a[159] & b[30])^(a[158] & b[31])^(a[157] & b[32])^(a[156] & b[33])^(a[155] & b[34])^(a[154] & b[35])^(a[153] & b[36])^(a[152] & b[37])^(a[151] & b[38])^(a[150] & b[39])^(a[149] & b[40])^(a[148] & b[41])^(a[147] & b[42])^(a[146] & b[43])^(a[145] & b[44])^(a[144] & b[45])^(a[143] & b[46])^(a[142] & b[47])^(a[141] & b[48])^(a[140] & b[49])^(a[139] & b[50])^(a[138] & b[51])^(a[137] & b[52])^(a[136] & b[53])^(a[135] & b[54])^(a[134] & b[55])^(a[133] & b[56])^(a[132] & b[57])^(a[131] & b[58])^(a[130] & b[59])^(a[129] & b[60])^(a[128] & b[61])^(a[127] & b[62])^(a[126] & b[63])^(a[125] & b[64])^(a[124] & b[65])^(a[123] & b[66])^(a[122] & b[67])^(a[121] & b[68])^(a[120] & b[69])^(a[119] & b[70])^(a[118] & b[71])^(a[117] & b[72])^(a[116] & b[73])^(a[115] & b[74])^(a[114] & b[75])^(a[113] & b[76])^(a[112] & b[77])^(a[111] & b[78])^(a[110] & b[79])^(a[109] & b[80])^(a[108] & b[81])^(a[107] & b[82])^(a[106] & b[83])^(a[105] & b[84])^(a[104] & b[85])^(a[103] & b[86])^(a[102] & b[87])^(a[101] & b[88])^(a[100] & b[89])^(a[99] & b[90])^(a[98] & b[91])^(a[97] & b[92])^(a[96] & b[93])^(a[95] & b[94])^(a[94] & b[95])^(a[93] & b[96])^(a[92] & b[97])^(a[91] & b[98])^(a[90] & b[99])^(a[89] & b[100])^(a[88] & b[101])^(a[87] & b[102])^(a[86] & b[103])^(a[85] & b[104])^(a[84] & b[105])^(a[83] & b[106])^(a[82] & b[107])^(a[81] & b[108])^(a[80] & b[109])^(a[79] & b[110])^(a[78] & b[111])^(a[77] & b[112])^(a[76] & b[113])^(a[75] & b[114])^(a[74] & b[115])^(a[73] & b[116])^(a[72] & b[117])^(a[71] & b[118])^(a[70] & b[119])^(a[69] & b[120])^(a[68] & b[121])^(a[67] & b[122])^(a[66] & b[123])^(a[65] & b[124])^(a[64] & b[125])^(a[63] & b[126])^(a[62] & b[127])^(a[61] & b[128])^(a[60] & b[129])^(a[59] & b[130])^(a[58] & b[131])^(a[57] & b[132])^(a[56] & b[133])^(a[55] & b[134])^(a[54] & b[135])^(a[53] & b[136])^(a[52] & b[137])^(a[51] & b[138])^(a[50] & b[139])^(a[49] & b[140])^(a[48] & b[141])^(a[47] & b[142])^(a[46] & b[143])^(a[45] & b[144])^(a[44] & b[145])^(a[43] & b[146])^(a[42] & b[147])^(a[41] & b[148])^(a[40] & b[149])^(a[39] & b[150])^(a[38] & b[151])^(a[37] & b[152])^(a[36] & b[153])^(a[35] & b[154])^(a[34] & b[155])^(a[33] & b[156])^(a[32] & b[157])^(a[31] & b[158])^(a[30] & b[159])^(a[29] & b[160])^(a[28] & b[161])^(a[27] & b[162]);
assign y[190] = (a[162] & b[28])^(a[161] & b[29])^(a[160] & b[30])^(a[159] & b[31])^(a[158] & b[32])^(a[157] & b[33])^(a[156] & b[34])^(a[155] & b[35])^(a[154] & b[36])^(a[153] & b[37])^(a[152] & b[38])^(a[151] & b[39])^(a[150] & b[40])^(a[149] & b[41])^(a[148] & b[42])^(a[147] & b[43])^(a[146] & b[44])^(a[145] & b[45])^(a[144] & b[46])^(a[143] & b[47])^(a[142] & b[48])^(a[141] & b[49])^(a[140] & b[50])^(a[139] & b[51])^(a[138] & b[52])^(a[137] & b[53])^(a[136] & b[54])^(a[135] & b[55])^(a[134] & b[56])^(a[133] & b[57])^(a[132] & b[58])^(a[131] & b[59])^(a[130] & b[60])^(a[129] & b[61])^(a[128] & b[62])^(a[127] & b[63])^(a[126] & b[64])^(a[125] & b[65])^(a[124] & b[66])^(a[123] & b[67])^(a[122] & b[68])^(a[121] & b[69])^(a[120] & b[70])^(a[119] & b[71])^(a[118] & b[72])^(a[117] & b[73])^(a[116] & b[74])^(a[115] & b[75])^(a[114] & b[76])^(a[113] & b[77])^(a[112] & b[78])^(a[111] & b[79])^(a[110] & b[80])^(a[109] & b[81])^(a[108] & b[82])^(a[107] & b[83])^(a[106] & b[84])^(a[105] & b[85])^(a[104] & b[86])^(a[103] & b[87])^(a[102] & b[88])^(a[101] & b[89])^(a[100] & b[90])^(a[99] & b[91])^(a[98] & b[92])^(a[97] & b[93])^(a[96] & b[94])^(a[95] & b[95])^(a[94] & b[96])^(a[93] & b[97])^(a[92] & b[98])^(a[91] & b[99])^(a[90] & b[100])^(a[89] & b[101])^(a[88] & b[102])^(a[87] & b[103])^(a[86] & b[104])^(a[85] & b[105])^(a[84] & b[106])^(a[83] & b[107])^(a[82] & b[108])^(a[81] & b[109])^(a[80] & b[110])^(a[79] & b[111])^(a[78] & b[112])^(a[77] & b[113])^(a[76] & b[114])^(a[75] & b[115])^(a[74] & b[116])^(a[73] & b[117])^(a[72] & b[118])^(a[71] & b[119])^(a[70] & b[120])^(a[69] & b[121])^(a[68] & b[122])^(a[67] & b[123])^(a[66] & b[124])^(a[65] & b[125])^(a[64] & b[126])^(a[63] & b[127])^(a[62] & b[128])^(a[61] & b[129])^(a[60] & b[130])^(a[59] & b[131])^(a[58] & b[132])^(a[57] & b[133])^(a[56] & b[134])^(a[55] & b[135])^(a[54] & b[136])^(a[53] & b[137])^(a[52] & b[138])^(a[51] & b[139])^(a[50] & b[140])^(a[49] & b[141])^(a[48] & b[142])^(a[47] & b[143])^(a[46] & b[144])^(a[45] & b[145])^(a[44] & b[146])^(a[43] & b[147])^(a[42] & b[148])^(a[41] & b[149])^(a[40] & b[150])^(a[39] & b[151])^(a[38] & b[152])^(a[37] & b[153])^(a[36] & b[154])^(a[35] & b[155])^(a[34] & b[156])^(a[33] & b[157])^(a[32] & b[158])^(a[31] & b[159])^(a[30] & b[160])^(a[29] & b[161])^(a[28] & b[162]);
assign y[191] = (a[162] & b[29])^(a[161] & b[30])^(a[160] & b[31])^(a[159] & b[32])^(a[158] & b[33])^(a[157] & b[34])^(a[156] & b[35])^(a[155] & b[36])^(a[154] & b[37])^(a[153] & b[38])^(a[152] & b[39])^(a[151] & b[40])^(a[150] & b[41])^(a[149] & b[42])^(a[148] & b[43])^(a[147] & b[44])^(a[146] & b[45])^(a[145] & b[46])^(a[144] & b[47])^(a[143] & b[48])^(a[142] & b[49])^(a[141] & b[50])^(a[140] & b[51])^(a[139] & b[52])^(a[138] & b[53])^(a[137] & b[54])^(a[136] & b[55])^(a[135] & b[56])^(a[134] & b[57])^(a[133] & b[58])^(a[132] & b[59])^(a[131] & b[60])^(a[130] & b[61])^(a[129] & b[62])^(a[128] & b[63])^(a[127] & b[64])^(a[126] & b[65])^(a[125] & b[66])^(a[124] & b[67])^(a[123] & b[68])^(a[122] & b[69])^(a[121] & b[70])^(a[120] & b[71])^(a[119] & b[72])^(a[118] & b[73])^(a[117] & b[74])^(a[116] & b[75])^(a[115] & b[76])^(a[114] & b[77])^(a[113] & b[78])^(a[112] & b[79])^(a[111] & b[80])^(a[110] & b[81])^(a[109] & b[82])^(a[108] & b[83])^(a[107] & b[84])^(a[106] & b[85])^(a[105] & b[86])^(a[104] & b[87])^(a[103] & b[88])^(a[102] & b[89])^(a[101] & b[90])^(a[100] & b[91])^(a[99] & b[92])^(a[98] & b[93])^(a[97] & b[94])^(a[96] & b[95])^(a[95] & b[96])^(a[94] & b[97])^(a[93] & b[98])^(a[92] & b[99])^(a[91] & b[100])^(a[90] & b[101])^(a[89] & b[102])^(a[88] & b[103])^(a[87] & b[104])^(a[86] & b[105])^(a[85] & b[106])^(a[84] & b[107])^(a[83] & b[108])^(a[82] & b[109])^(a[81] & b[110])^(a[80] & b[111])^(a[79] & b[112])^(a[78] & b[113])^(a[77] & b[114])^(a[76] & b[115])^(a[75] & b[116])^(a[74] & b[117])^(a[73] & b[118])^(a[72] & b[119])^(a[71] & b[120])^(a[70] & b[121])^(a[69] & b[122])^(a[68] & b[123])^(a[67] & b[124])^(a[66] & b[125])^(a[65] & b[126])^(a[64] & b[127])^(a[63] & b[128])^(a[62] & b[129])^(a[61] & b[130])^(a[60] & b[131])^(a[59] & b[132])^(a[58] & b[133])^(a[57] & b[134])^(a[56] & b[135])^(a[55] & b[136])^(a[54] & b[137])^(a[53] & b[138])^(a[52] & b[139])^(a[51] & b[140])^(a[50] & b[141])^(a[49] & b[142])^(a[48] & b[143])^(a[47] & b[144])^(a[46] & b[145])^(a[45] & b[146])^(a[44] & b[147])^(a[43] & b[148])^(a[42] & b[149])^(a[41] & b[150])^(a[40] & b[151])^(a[39] & b[152])^(a[38] & b[153])^(a[37] & b[154])^(a[36] & b[155])^(a[35] & b[156])^(a[34] & b[157])^(a[33] & b[158])^(a[32] & b[159])^(a[31] & b[160])^(a[30] & b[161])^(a[29] & b[162]);
assign y[192] = (a[162] & b[30])^(a[161] & b[31])^(a[160] & b[32])^(a[159] & b[33])^(a[158] & b[34])^(a[157] & b[35])^(a[156] & b[36])^(a[155] & b[37])^(a[154] & b[38])^(a[153] & b[39])^(a[152] & b[40])^(a[151] & b[41])^(a[150] & b[42])^(a[149] & b[43])^(a[148] & b[44])^(a[147] & b[45])^(a[146] & b[46])^(a[145] & b[47])^(a[144] & b[48])^(a[143] & b[49])^(a[142] & b[50])^(a[141] & b[51])^(a[140] & b[52])^(a[139] & b[53])^(a[138] & b[54])^(a[137] & b[55])^(a[136] & b[56])^(a[135] & b[57])^(a[134] & b[58])^(a[133] & b[59])^(a[132] & b[60])^(a[131] & b[61])^(a[130] & b[62])^(a[129] & b[63])^(a[128] & b[64])^(a[127] & b[65])^(a[126] & b[66])^(a[125] & b[67])^(a[124] & b[68])^(a[123] & b[69])^(a[122] & b[70])^(a[121] & b[71])^(a[120] & b[72])^(a[119] & b[73])^(a[118] & b[74])^(a[117] & b[75])^(a[116] & b[76])^(a[115] & b[77])^(a[114] & b[78])^(a[113] & b[79])^(a[112] & b[80])^(a[111] & b[81])^(a[110] & b[82])^(a[109] & b[83])^(a[108] & b[84])^(a[107] & b[85])^(a[106] & b[86])^(a[105] & b[87])^(a[104] & b[88])^(a[103] & b[89])^(a[102] & b[90])^(a[101] & b[91])^(a[100] & b[92])^(a[99] & b[93])^(a[98] & b[94])^(a[97] & b[95])^(a[96] & b[96])^(a[95] & b[97])^(a[94] & b[98])^(a[93] & b[99])^(a[92] & b[100])^(a[91] & b[101])^(a[90] & b[102])^(a[89] & b[103])^(a[88] & b[104])^(a[87] & b[105])^(a[86] & b[106])^(a[85] & b[107])^(a[84] & b[108])^(a[83] & b[109])^(a[82] & b[110])^(a[81] & b[111])^(a[80] & b[112])^(a[79] & b[113])^(a[78] & b[114])^(a[77] & b[115])^(a[76] & b[116])^(a[75] & b[117])^(a[74] & b[118])^(a[73] & b[119])^(a[72] & b[120])^(a[71] & b[121])^(a[70] & b[122])^(a[69] & b[123])^(a[68] & b[124])^(a[67] & b[125])^(a[66] & b[126])^(a[65] & b[127])^(a[64] & b[128])^(a[63] & b[129])^(a[62] & b[130])^(a[61] & b[131])^(a[60] & b[132])^(a[59] & b[133])^(a[58] & b[134])^(a[57] & b[135])^(a[56] & b[136])^(a[55] & b[137])^(a[54] & b[138])^(a[53] & b[139])^(a[52] & b[140])^(a[51] & b[141])^(a[50] & b[142])^(a[49] & b[143])^(a[48] & b[144])^(a[47] & b[145])^(a[46] & b[146])^(a[45] & b[147])^(a[44] & b[148])^(a[43] & b[149])^(a[42] & b[150])^(a[41] & b[151])^(a[40] & b[152])^(a[39] & b[153])^(a[38] & b[154])^(a[37] & b[155])^(a[36] & b[156])^(a[35] & b[157])^(a[34] & b[158])^(a[33] & b[159])^(a[32] & b[160])^(a[31] & b[161])^(a[30] & b[162]);
assign y[193] = (a[162] & b[31])^(a[161] & b[32])^(a[160] & b[33])^(a[159] & b[34])^(a[158] & b[35])^(a[157] & b[36])^(a[156] & b[37])^(a[155] & b[38])^(a[154] & b[39])^(a[153] & b[40])^(a[152] & b[41])^(a[151] & b[42])^(a[150] & b[43])^(a[149] & b[44])^(a[148] & b[45])^(a[147] & b[46])^(a[146] & b[47])^(a[145] & b[48])^(a[144] & b[49])^(a[143] & b[50])^(a[142] & b[51])^(a[141] & b[52])^(a[140] & b[53])^(a[139] & b[54])^(a[138] & b[55])^(a[137] & b[56])^(a[136] & b[57])^(a[135] & b[58])^(a[134] & b[59])^(a[133] & b[60])^(a[132] & b[61])^(a[131] & b[62])^(a[130] & b[63])^(a[129] & b[64])^(a[128] & b[65])^(a[127] & b[66])^(a[126] & b[67])^(a[125] & b[68])^(a[124] & b[69])^(a[123] & b[70])^(a[122] & b[71])^(a[121] & b[72])^(a[120] & b[73])^(a[119] & b[74])^(a[118] & b[75])^(a[117] & b[76])^(a[116] & b[77])^(a[115] & b[78])^(a[114] & b[79])^(a[113] & b[80])^(a[112] & b[81])^(a[111] & b[82])^(a[110] & b[83])^(a[109] & b[84])^(a[108] & b[85])^(a[107] & b[86])^(a[106] & b[87])^(a[105] & b[88])^(a[104] & b[89])^(a[103] & b[90])^(a[102] & b[91])^(a[101] & b[92])^(a[100] & b[93])^(a[99] & b[94])^(a[98] & b[95])^(a[97] & b[96])^(a[96] & b[97])^(a[95] & b[98])^(a[94] & b[99])^(a[93] & b[100])^(a[92] & b[101])^(a[91] & b[102])^(a[90] & b[103])^(a[89] & b[104])^(a[88] & b[105])^(a[87] & b[106])^(a[86] & b[107])^(a[85] & b[108])^(a[84] & b[109])^(a[83] & b[110])^(a[82] & b[111])^(a[81] & b[112])^(a[80] & b[113])^(a[79] & b[114])^(a[78] & b[115])^(a[77] & b[116])^(a[76] & b[117])^(a[75] & b[118])^(a[74] & b[119])^(a[73] & b[120])^(a[72] & b[121])^(a[71] & b[122])^(a[70] & b[123])^(a[69] & b[124])^(a[68] & b[125])^(a[67] & b[126])^(a[66] & b[127])^(a[65] & b[128])^(a[64] & b[129])^(a[63] & b[130])^(a[62] & b[131])^(a[61] & b[132])^(a[60] & b[133])^(a[59] & b[134])^(a[58] & b[135])^(a[57] & b[136])^(a[56] & b[137])^(a[55] & b[138])^(a[54] & b[139])^(a[53] & b[140])^(a[52] & b[141])^(a[51] & b[142])^(a[50] & b[143])^(a[49] & b[144])^(a[48] & b[145])^(a[47] & b[146])^(a[46] & b[147])^(a[45] & b[148])^(a[44] & b[149])^(a[43] & b[150])^(a[42] & b[151])^(a[41] & b[152])^(a[40] & b[153])^(a[39] & b[154])^(a[38] & b[155])^(a[37] & b[156])^(a[36] & b[157])^(a[35] & b[158])^(a[34] & b[159])^(a[33] & b[160])^(a[32] & b[161])^(a[31] & b[162]);
assign y[194] = (a[162] & b[32])^(a[161] & b[33])^(a[160] & b[34])^(a[159] & b[35])^(a[158] & b[36])^(a[157] & b[37])^(a[156] & b[38])^(a[155] & b[39])^(a[154] & b[40])^(a[153] & b[41])^(a[152] & b[42])^(a[151] & b[43])^(a[150] & b[44])^(a[149] & b[45])^(a[148] & b[46])^(a[147] & b[47])^(a[146] & b[48])^(a[145] & b[49])^(a[144] & b[50])^(a[143] & b[51])^(a[142] & b[52])^(a[141] & b[53])^(a[140] & b[54])^(a[139] & b[55])^(a[138] & b[56])^(a[137] & b[57])^(a[136] & b[58])^(a[135] & b[59])^(a[134] & b[60])^(a[133] & b[61])^(a[132] & b[62])^(a[131] & b[63])^(a[130] & b[64])^(a[129] & b[65])^(a[128] & b[66])^(a[127] & b[67])^(a[126] & b[68])^(a[125] & b[69])^(a[124] & b[70])^(a[123] & b[71])^(a[122] & b[72])^(a[121] & b[73])^(a[120] & b[74])^(a[119] & b[75])^(a[118] & b[76])^(a[117] & b[77])^(a[116] & b[78])^(a[115] & b[79])^(a[114] & b[80])^(a[113] & b[81])^(a[112] & b[82])^(a[111] & b[83])^(a[110] & b[84])^(a[109] & b[85])^(a[108] & b[86])^(a[107] & b[87])^(a[106] & b[88])^(a[105] & b[89])^(a[104] & b[90])^(a[103] & b[91])^(a[102] & b[92])^(a[101] & b[93])^(a[100] & b[94])^(a[99] & b[95])^(a[98] & b[96])^(a[97] & b[97])^(a[96] & b[98])^(a[95] & b[99])^(a[94] & b[100])^(a[93] & b[101])^(a[92] & b[102])^(a[91] & b[103])^(a[90] & b[104])^(a[89] & b[105])^(a[88] & b[106])^(a[87] & b[107])^(a[86] & b[108])^(a[85] & b[109])^(a[84] & b[110])^(a[83] & b[111])^(a[82] & b[112])^(a[81] & b[113])^(a[80] & b[114])^(a[79] & b[115])^(a[78] & b[116])^(a[77] & b[117])^(a[76] & b[118])^(a[75] & b[119])^(a[74] & b[120])^(a[73] & b[121])^(a[72] & b[122])^(a[71] & b[123])^(a[70] & b[124])^(a[69] & b[125])^(a[68] & b[126])^(a[67] & b[127])^(a[66] & b[128])^(a[65] & b[129])^(a[64] & b[130])^(a[63] & b[131])^(a[62] & b[132])^(a[61] & b[133])^(a[60] & b[134])^(a[59] & b[135])^(a[58] & b[136])^(a[57] & b[137])^(a[56] & b[138])^(a[55] & b[139])^(a[54] & b[140])^(a[53] & b[141])^(a[52] & b[142])^(a[51] & b[143])^(a[50] & b[144])^(a[49] & b[145])^(a[48] & b[146])^(a[47] & b[147])^(a[46] & b[148])^(a[45] & b[149])^(a[44] & b[150])^(a[43] & b[151])^(a[42] & b[152])^(a[41] & b[153])^(a[40] & b[154])^(a[39] & b[155])^(a[38] & b[156])^(a[37] & b[157])^(a[36] & b[158])^(a[35] & b[159])^(a[34] & b[160])^(a[33] & b[161])^(a[32] & b[162]);
assign y[195] = (a[162] & b[33])^(a[161] & b[34])^(a[160] & b[35])^(a[159] & b[36])^(a[158] & b[37])^(a[157] & b[38])^(a[156] & b[39])^(a[155] & b[40])^(a[154] & b[41])^(a[153] & b[42])^(a[152] & b[43])^(a[151] & b[44])^(a[150] & b[45])^(a[149] & b[46])^(a[148] & b[47])^(a[147] & b[48])^(a[146] & b[49])^(a[145] & b[50])^(a[144] & b[51])^(a[143] & b[52])^(a[142] & b[53])^(a[141] & b[54])^(a[140] & b[55])^(a[139] & b[56])^(a[138] & b[57])^(a[137] & b[58])^(a[136] & b[59])^(a[135] & b[60])^(a[134] & b[61])^(a[133] & b[62])^(a[132] & b[63])^(a[131] & b[64])^(a[130] & b[65])^(a[129] & b[66])^(a[128] & b[67])^(a[127] & b[68])^(a[126] & b[69])^(a[125] & b[70])^(a[124] & b[71])^(a[123] & b[72])^(a[122] & b[73])^(a[121] & b[74])^(a[120] & b[75])^(a[119] & b[76])^(a[118] & b[77])^(a[117] & b[78])^(a[116] & b[79])^(a[115] & b[80])^(a[114] & b[81])^(a[113] & b[82])^(a[112] & b[83])^(a[111] & b[84])^(a[110] & b[85])^(a[109] & b[86])^(a[108] & b[87])^(a[107] & b[88])^(a[106] & b[89])^(a[105] & b[90])^(a[104] & b[91])^(a[103] & b[92])^(a[102] & b[93])^(a[101] & b[94])^(a[100] & b[95])^(a[99] & b[96])^(a[98] & b[97])^(a[97] & b[98])^(a[96] & b[99])^(a[95] & b[100])^(a[94] & b[101])^(a[93] & b[102])^(a[92] & b[103])^(a[91] & b[104])^(a[90] & b[105])^(a[89] & b[106])^(a[88] & b[107])^(a[87] & b[108])^(a[86] & b[109])^(a[85] & b[110])^(a[84] & b[111])^(a[83] & b[112])^(a[82] & b[113])^(a[81] & b[114])^(a[80] & b[115])^(a[79] & b[116])^(a[78] & b[117])^(a[77] & b[118])^(a[76] & b[119])^(a[75] & b[120])^(a[74] & b[121])^(a[73] & b[122])^(a[72] & b[123])^(a[71] & b[124])^(a[70] & b[125])^(a[69] & b[126])^(a[68] & b[127])^(a[67] & b[128])^(a[66] & b[129])^(a[65] & b[130])^(a[64] & b[131])^(a[63] & b[132])^(a[62] & b[133])^(a[61] & b[134])^(a[60] & b[135])^(a[59] & b[136])^(a[58] & b[137])^(a[57] & b[138])^(a[56] & b[139])^(a[55] & b[140])^(a[54] & b[141])^(a[53] & b[142])^(a[52] & b[143])^(a[51] & b[144])^(a[50] & b[145])^(a[49] & b[146])^(a[48] & b[147])^(a[47] & b[148])^(a[46] & b[149])^(a[45] & b[150])^(a[44] & b[151])^(a[43] & b[152])^(a[42] & b[153])^(a[41] & b[154])^(a[40] & b[155])^(a[39] & b[156])^(a[38] & b[157])^(a[37] & b[158])^(a[36] & b[159])^(a[35] & b[160])^(a[34] & b[161])^(a[33] & b[162]);
assign y[196] = (a[162] & b[34])^(a[161] & b[35])^(a[160] & b[36])^(a[159] & b[37])^(a[158] & b[38])^(a[157] & b[39])^(a[156] & b[40])^(a[155] & b[41])^(a[154] & b[42])^(a[153] & b[43])^(a[152] & b[44])^(a[151] & b[45])^(a[150] & b[46])^(a[149] & b[47])^(a[148] & b[48])^(a[147] & b[49])^(a[146] & b[50])^(a[145] & b[51])^(a[144] & b[52])^(a[143] & b[53])^(a[142] & b[54])^(a[141] & b[55])^(a[140] & b[56])^(a[139] & b[57])^(a[138] & b[58])^(a[137] & b[59])^(a[136] & b[60])^(a[135] & b[61])^(a[134] & b[62])^(a[133] & b[63])^(a[132] & b[64])^(a[131] & b[65])^(a[130] & b[66])^(a[129] & b[67])^(a[128] & b[68])^(a[127] & b[69])^(a[126] & b[70])^(a[125] & b[71])^(a[124] & b[72])^(a[123] & b[73])^(a[122] & b[74])^(a[121] & b[75])^(a[120] & b[76])^(a[119] & b[77])^(a[118] & b[78])^(a[117] & b[79])^(a[116] & b[80])^(a[115] & b[81])^(a[114] & b[82])^(a[113] & b[83])^(a[112] & b[84])^(a[111] & b[85])^(a[110] & b[86])^(a[109] & b[87])^(a[108] & b[88])^(a[107] & b[89])^(a[106] & b[90])^(a[105] & b[91])^(a[104] & b[92])^(a[103] & b[93])^(a[102] & b[94])^(a[101] & b[95])^(a[100] & b[96])^(a[99] & b[97])^(a[98] & b[98])^(a[97] & b[99])^(a[96] & b[100])^(a[95] & b[101])^(a[94] & b[102])^(a[93] & b[103])^(a[92] & b[104])^(a[91] & b[105])^(a[90] & b[106])^(a[89] & b[107])^(a[88] & b[108])^(a[87] & b[109])^(a[86] & b[110])^(a[85] & b[111])^(a[84] & b[112])^(a[83] & b[113])^(a[82] & b[114])^(a[81] & b[115])^(a[80] & b[116])^(a[79] & b[117])^(a[78] & b[118])^(a[77] & b[119])^(a[76] & b[120])^(a[75] & b[121])^(a[74] & b[122])^(a[73] & b[123])^(a[72] & b[124])^(a[71] & b[125])^(a[70] & b[126])^(a[69] & b[127])^(a[68] & b[128])^(a[67] & b[129])^(a[66] & b[130])^(a[65] & b[131])^(a[64] & b[132])^(a[63] & b[133])^(a[62] & b[134])^(a[61] & b[135])^(a[60] & b[136])^(a[59] & b[137])^(a[58] & b[138])^(a[57] & b[139])^(a[56] & b[140])^(a[55] & b[141])^(a[54] & b[142])^(a[53] & b[143])^(a[52] & b[144])^(a[51] & b[145])^(a[50] & b[146])^(a[49] & b[147])^(a[48] & b[148])^(a[47] & b[149])^(a[46] & b[150])^(a[45] & b[151])^(a[44] & b[152])^(a[43] & b[153])^(a[42] & b[154])^(a[41] & b[155])^(a[40] & b[156])^(a[39] & b[157])^(a[38] & b[158])^(a[37] & b[159])^(a[36] & b[160])^(a[35] & b[161])^(a[34] & b[162]);
assign y[197] = (a[162] & b[35])^(a[161] & b[36])^(a[160] & b[37])^(a[159] & b[38])^(a[158] & b[39])^(a[157] & b[40])^(a[156] & b[41])^(a[155] & b[42])^(a[154] & b[43])^(a[153] & b[44])^(a[152] & b[45])^(a[151] & b[46])^(a[150] & b[47])^(a[149] & b[48])^(a[148] & b[49])^(a[147] & b[50])^(a[146] & b[51])^(a[145] & b[52])^(a[144] & b[53])^(a[143] & b[54])^(a[142] & b[55])^(a[141] & b[56])^(a[140] & b[57])^(a[139] & b[58])^(a[138] & b[59])^(a[137] & b[60])^(a[136] & b[61])^(a[135] & b[62])^(a[134] & b[63])^(a[133] & b[64])^(a[132] & b[65])^(a[131] & b[66])^(a[130] & b[67])^(a[129] & b[68])^(a[128] & b[69])^(a[127] & b[70])^(a[126] & b[71])^(a[125] & b[72])^(a[124] & b[73])^(a[123] & b[74])^(a[122] & b[75])^(a[121] & b[76])^(a[120] & b[77])^(a[119] & b[78])^(a[118] & b[79])^(a[117] & b[80])^(a[116] & b[81])^(a[115] & b[82])^(a[114] & b[83])^(a[113] & b[84])^(a[112] & b[85])^(a[111] & b[86])^(a[110] & b[87])^(a[109] & b[88])^(a[108] & b[89])^(a[107] & b[90])^(a[106] & b[91])^(a[105] & b[92])^(a[104] & b[93])^(a[103] & b[94])^(a[102] & b[95])^(a[101] & b[96])^(a[100] & b[97])^(a[99] & b[98])^(a[98] & b[99])^(a[97] & b[100])^(a[96] & b[101])^(a[95] & b[102])^(a[94] & b[103])^(a[93] & b[104])^(a[92] & b[105])^(a[91] & b[106])^(a[90] & b[107])^(a[89] & b[108])^(a[88] & b[109])^(a[87] & b[110])^(a[86] & b[111])^(a[85] & b[112])^(a[84] & b[113])^(a[83] & b[114])^(a[82] & b[115])^(a[81] & b[116])^(a[80] & b[117])^(a[79] & b[118])^(a[78] & b[119])^(a[77] & b[120])^(a[76] & b[121])^(a[75] & b[122])^(a[74] & b[123])^(a[73] & b[124])^(a[72] & b[125])^(a[71] & b[126])^(a[70] & b[127])^(a[69] & b[128])^(a[68] & b[129])^(a[67] & b[130])^(a[66] & b[131])^(a[65] & b[132])^(a[64] & b[133])^(a[63] & b[134])^(a[62] & b[135])^(a[61] & b[136])^(a[60] & b[137])^(a[59] & b[138])^(a[58] & b[139])^(a[57] & b[140])^(a[56] & b[141])^(a[55] & b[142])^(a[54] & b[143])^(a[53] & b[144])^(a[52] & b[145])^(a[51] & b[146])^(a[50] & b[147])^(a[49] & b[148])^(a[48] & b[149])^(a[47] & b[150])^(a[46] & b[151])^(a[45] & b[152])^(a[44] & b[153])^(a[43] & b[154])^(a[42] & b[155])^(a[41] & b[156])^(a[40] & b[157])^(a[39] & b[158])^(a[38] & b[159])^(a[37] & b[160])^(a[36] & b[161])^(a[35] & b[162]);
assign y[198] = (a[162] & b[36])^(a[161] & b[37])^(a[160] & b[38])^(a[159] & b[39])^(a[158] & b[40])^(a[157] & b[41])^(a[156] & b[42])^(a[155] & b[43])^(a[154] & b[44])^(a[153] & b[45])^(a[152] & b[46])^(a[151] & b[47])^(a[150] & b[48])^(a[149] & b[49])^(a[148] & b[50])^(a[147] & b[51])^(a[146] & b[52])^(a[145] & b[53])^(a[144] & b[54])^(a[143] & b[55])^(a[142] & b[56])^(a[141] & b[57])^(a[140] & b[58])^(a[139] & b[59])^(a[138] & b[60])^(a[137] & b[61])^(a[136] & b[62])^(a[135] & b[63])^(a[134] & b[64])^(a[133] & b[65])^(a[132] & b[66])^(a[131] & b[67])^(a[130] & b[68])^(a[129] & b[69])^(a[128] & b[70])^(a[127] & b[71])^(a[126] & b[72])^(a[125] & b[73])^(a[124] & b[74])^(a[123] & b[75])^(a[122] & b[76])^(a[121] & b[77])^(a[120] & b[78])^(a[119] & b[79])^(a[118] & b[80])^(a[117] & b[81])^(a[116] & b[82])^(a[115] & b[83])^(a[114] & b[84])^(a[113] & b[85])^(a[112] & b[86])^(a[111] & b[87])^(a[110] & b[88])^(a[109] & b[89])^(a[108] & b[90])^(a[107] & b[91])^(a[106] & b[92])^(a[105] & b[93])^(a[104] & b[94])^(a[103] & b[95])^(a[102] & b[96])^(a[101] & b[97])^(a[100] & b[98])^(a[99] & b[99])^(a[98] & b[100])^(a[97] & b[101])^(a[96] & b[102])^(a[95] & b[103])^(a[94] & b[104])^(a[93] & b[105])^(a[92] & b[106])^(a[91] & b[107])^(a[90] & b[108])^(a[89] & b[109])^(a[88] & b[110])^(a[87] & b[111])^(a[86] & b[112])^(a[85] & b[113])^(a[84] & b[114])^(a[83] & b[115])^(a[82] & b[116])^(a[81] & b[117])^(a[80] & b[118])^(a[79] & b[119])^(a[78] & b[120])^(a[77] & b[121])^(a[76] & b[122])^(a[75] & b[123])^(a[74] & b[124])^(a[73] & b[125])^(a[72] & b[126])^(a[71] & b[127])^(a[70] & b[128])^(a[69] & b[129])^(a[68] & b[130])^(a[67] & b[131])^(a[66] & b[132])^(a[65] & b[133])^(a[64] & b[134])^(a[63] & b[135])^(a[62] & b[136])^(a[61] & b[137])^(a[60] & b[138])^(a[59] & b[139])^(a[58] & b[140])^(a[57] & b[141])^(a[56] & b[142])^(a[55] & b[143])^(a[54] & b[144])^(a[53] & b[145])^(a[52] & b[146])^(a[51] & b[147])^(a[50] & b[148])^(a[49] & b[149])^(a[48] & b[150])^(a[47] & b[151])^(a[46] & b[152])^(a[45] & b[153])^(a[44] & b[154])^(a[43] & b[155])^(a[42] & b[156])^(a[41] & b[157])^(a[40] & b[158])^(a[39] & b[159])^(a[38] & b[160])^(a[37] & b[161])^(a[36] & b[162]);
assign y[199] = (a[162] & b[37])^(a[161] & b[38])^(a[160] & b[39])^(a[159] & b[40])^(a[158] & b[41])^(a[157] & b[42])^(a[156] & b[43])^(a[155] & b[44])^(a[154] & b[45])^(a[153] & b[46])^(a[152] & b[47])^(a[151] & b[48])^(a[150] & b[49])^(a[149] & b[50])^(a[148] & b[51])^(a[147] & b[52])^(a[146] & b[53])^(a[145] & b[54])^(a[144] & b[55])^(a[143] & b[56])^(a[142] & b[57])^(a[141] & b[58])^(a[140] & b[59])^(a[139] & b[60])^(a[138] & b[61])^(a[137] & b[62])^(a[136] & b[63])^(a[135] & b[64])^(a[134] & b[65])^(a[133] & b[66])^(a[132] & b[67])^(a[131] & b[68])^(a[130] & b[69])^(a[129] & b[70])^(a[128] & b[71])^(a[127] & b[72])^(a[126] & b[73])^(a[125] & b[74])^(a[124] & b[75])^(a[123] & b[76])^(a[122] & b[77])^(a[121] & b[78])^(a[120] & b[79])^(a[119] & b[80])^(a[118] & b[81])^(a[117] & b[82])^(a[116] & b[83])^(a[115] & b[84])^(a[114] & b[85])^(a[113] & b[86])^(a[112] & b[87])^(a[111] & b[88])^(a[110] & b[89])^(a[109] & b[90])^(a[108] & b[91])^(a[107] & b[92])^(a[106] & b[93])^(a[105] & b[94])^(a[104] & b[95])^(a[103] & b[96])^(a[102] & b[97])^(a[101] & b[98])^(a[100] & b[99])^(a[99] & b[100])^(a[98] & b[101])^(a[97] & b[102])^(a[96] & b[103])^(a[95] & b[104])^(a[94] & b[105])^(a[93] & b[106])^(a[92] & b[107])^(a[91] & b[108])^(a[90] & b[109])^(a[89] & b[110])^(a[88] & b[111])^(a[87] & b[112])^(a[86] & b[113])^(a[85] & b[114])^(a[84] & b[115])^(a[83] & b[116])^(a[82] & b[117])^(a[81] & b[118])^(a[80] & b[119])^(a[79] & b[120])^(a[78] & b[121])^(a[77] & b[122])^(a[76] & b[123])^(a[75] & b[124])^(a[74] & b[125])^(a[73] & b[126])^(a[72] & b[127])^(a[71] & b[128])^(a[70] & b[129])^(a[69] & b[130])^(a[68] & b[131])^(a[67] & b[132])^(a[66] & b[133])^(a[65] & b[134])^(a[64] & b[135])^(a[63] & b[136])^(a[62] & b[137])^(a[61] & b[138])^(a[60] & b[139])^(a[59] & b[140])^(a[58] & b[141])^(a[57] & b[142])^(a[56] & b[143])^(a[55] & b[144])^(a[54] & b[145])^(a[53] & b[146])^(a[52] & b[147])^(a[51] & b[148])^(a[50] & b[149])^(a[49] & b[150])^(a[48] & b[151])^(a[47] & b[152])^(a[46] & b[153])^(a[45] & b[154])^(a[44] & b[155])^(a[43] & b[156])^(a[42] & b[157])^(a[41] & b[158])^(a[40] & b[159])^(a[39] & b[160])^(a[38] & b[161])^(a[37] & b[162]);
assign y[200] = (a[162] & b[38])^(a[161] & b[39])^(a[160] & b[40])^(a[159] & b[41])^(a[158] & b[42])^(a[157] & b[43])^(a[156] & b[44])^(a[155] & b[45])^(a[154] & b[46])^(a[153] & b[47])^(a[152] & b[48])^(a[151] & b[49])^(a[150] & b[50])^(a[149] & b[51])^(a[148] & b[52])^(a[147] & b[53])^(a[146] & b[54])^(a[145] & b[55])^(a[144] & b[56])^(a[143] & b[57])^(a[142] & b[58])^(a[141] & b[59])^(a[140] & b[60])^(a[139] & b[61])^(a[138] & b[62])^(a[137] & b[63])^(a[136] & b[64])^(a[135] & b[65])^(a[134] & b[66])^(a[133] & b[67])^(a[132] & b[68])^(a[131] & b[69])^(a[130] & b[70])^(a[129] & b[71])^(a[128] & b[72])^(a[127] & b[73])^(a[126] & b[74])^(a[125] & b[75])^(a[124] & b[76])^(a[123] & b[77])^(a[122] & b[78])^(a[121] & b[79])^(a[120] & b[80])^(a[119] & b[81])^(a[118] & b[82])^(a[117] & b[83])^(a[116] & b[84])^(a[115] & b[85])^(a[114] & b[86])^(a[113] & b[87])^(a[112] & b[88])^(a[111] & b[89])^(a[110] & b[90])^(a[109] & b[91])^(a[108] & b[92])^(a[107] & b[93])^(a[106] & b[94])^(a[105] & b[95])^(a[104] & b[96])^(a[103] & b[97])^(a[102] & b[98])^(a[101] & b[99])^(a[100] & b[100])^(a[99] & b[101])^(a[98] & b[102])^(a[97] & b[103])^(a[96] & b[104])^(a[95] & b[105])^(a[94] & b[106])^(a[93] & b[107])^(a[92] & b[108])^(a[91] & b[109])^(a[90] & b[110])^(a[89] & b[111])^(a[88] & b[112])^(a[87] & b[113])^(a[86] & b[114])^(a[85] & b[115])^(a[84] & b[116])^(a[83] & b[117])^(a[82] & b[118])^(a[81] & b[119])^(a[80] & b[120])^(a[79] & b[121])^(a[78] & b[122])^(a[77] & b[123])^(a[76] & b[124])^(a[75] & b[125])^(a[74] & b[126])^(a[73] & b[127])^(a[72] & b[128])^(a[71] & b[129])^(a[70] & b[130])^(a[69] & b[131])^(a[68] & b[132])^(a[67] & b[133])^(a[66] & b[134])^(a[65] & b[135])^(a[64] & b[136])^(a[63] & b[137])^(a[62] & b[138])^(a[61] & b[139])^(a[60] & b[140])^(a[59] & b[141])^(a[58] & b[142])^(a[57] & b[143])^(a[56] & b[144])^(a[55] & b[145])^(a[54] & b[146])^(a[53] & b[147])^(a[52] & b[148])^(a[51] & b[149])^(a[50] & b[150])^(a[49] & b[151])^(a[48] & b[152])^(a[47] & b[153])^(a[46] & b[154])^(a[45] & b[155])^(a[44] & b[156])^(a[43] & b[157])^(a[42] & b[158])^(a[41] & b[159])^(a[40] & b[160])^(a[39] & b[161])^(a[38] & b[162]);
assign y[201] = (a[162] & b[39])^(a[161] & b[40])^(a[160] & b[41])^(a[159] & b[42])^(a[158] & b[43])^(a[157] & b[44])^(a[156] & b[45])^(a[155] & b[46])^(a[154] & b[47])^(a[153] & b[48])^(a[152] & b[49])^(a[151] & b[50])^(a[150] & b[51])^(a[149] & b[52])^(a[148] & b[53])^(a[147] & b[54])^(a[146] & b[55])^(a[145] & b[56])^(a[144] & b[57])^(a[143] & b[58])^(a[142] & b[59])^(a[141] & b[60])^(a[140] & b[61])^(a[139] & b[62])^(a[138] & b[63])^(a[137] & b[64])^(a[136] & b[65])^(a[135] & b[66])^(a[134] & b[67])^(a[133] & b[68])^(a[132] & b[69])^(a[131] & b[70])^(a[130] & b[71])^(a[129] & b[72])^(a[128] & b[73])^(a[127] & b[74])^(a[126] & b[75])^(a[125] & b[76])^(a[124] & b[77])^(a[123] & b[78])^(a[122] & b[79])^(a[121] & b[80])^(a[120] & b[81])^(a[119] & b[82])^(a[118] & b[83])^(a[117] & b[84])^(a[116] & b[85])^(a[115] & b[86])^(a[114] & b[87])^(a[113] & b[88])^(a[112] & b[89])^(a[111] & b[90])^(a[110] & b[91])^(a[109] & b[92])^(a[108] & b[93])^(a[107] & b[94])^(a[106] & b[95])^(a[105] & b[96])^(a[104] & b[97])^(a[103] & b[98])^(a[102] & b[99])^(a[101] & b[100])^(a[100] & b[101])^(a[99] & b[102])^(a[98] & b[103])^(a[97] & b[104])^(a[96] & b[105])^(a[95] & b[106])^(a[94] & b[107])^(a[93] & b[108])^(a[92] & b[109])^(a[91] & b[110])^(a[90] & b[111])^(a[89] & b[112])^(a[88] & b[113])^(a[87] & b[114])^(a[86] & b[115])^(a[85] & b[116])^(a[84] & b[117])^(a[83] & b[118])^(a[82] & b[119])^(a[81] & b[120])^(a[80] & b[121])^(a[79] & b[122])^(a[78] & b[123])^(a[77] & b[124])^(a[76] & b[125])^(a[75] & b[126])^(a[74] & b[127])^(a[73] & b[128])^(a[72] & b[129])^(a[71] & b[130])^(a[70] & b[131])^(a[69] & b[132])^(a[68] & b[133])^(a[67] & b[134])^(a[66] & b[135])^(a[65] & b[136])^(a[64] & b[137])^(a[63] & b[138])^(a[62] & b[139])^(a[61] & b[140])^(a[60] & b[141])^(a[59] & b[142])^(a[58] & b[143])^(a[57] & b[144])^(a[56] & b[145])^(a[55] & b[146])^(a[54] & b[147])^(a[53] & b[148])^(a[52] & b[149])^(a[51] & b[150])^(a[50] & b[151])^(a[49] & b[152])^(a[48] & b[153])^(a[47] & b[154])^(a[46] & b[155])^(a[45] & b[156])^(a[44] & b[157])^(a[43] & b[158])^(a[42] & b[159])^(a[41] & b[160])^(a[40] & b[161])^(a[39] & b[162]);
assign y[202] = (a[162] & b[40])^(a[161] & b[41])^(a[160] & b[42])^(a[159] & b[43])^(a[158] & b[44])^(a[157] & b[45])^(a[156] & b[46])^(a[155] & b[47])^(a[154] & b[48])^(a[153] & b[49])^(a[152] & b[50])^(a[151] & b[51])^(a[150] & b[52])^(a[149] & b[53])^(a[148] & b[54])^(a[147] & b[55])^(a[146] & b[56])^(a[145] & b[57])^(a[144] & b[58])^(a[143] & b[59])^(a[142] & b[60])^(a[141] & b[61])^(a[140] & b[62])^(a[139] & b[63])^(a[138] & b[64])^(a[137] & b[65])^(a[136] & b[66])^(a[135] & b[67])^(a[134] & b[68])^(a[133] & b[69])^(a[132] & b[70])^(a[131] & b[71])^(a[130] & b[72])^(a[129] & b[73])^(a[128] & b[74])^(a[127] & b[75])^(a[126] & b[76])^(a[125] & b[77])^(a[124] & b[78])^(a[123] & b[79])^(a[122] & b[80])^(a[121] & b[81])^(a[120] & b[82])^(a[119] & b[83])^(a[118] & b[84])^(a[117] & b[85])^(a[116] & b[86])^(a[115] & b[87])^(a[114] & b[88])^(a[113] & b[89])^(a[112] & b[90])^(a[111] & b[91])^(a[110] & b[92])^(a[109] & b[93])^(a[108] & b[94])^(a[107] & b[95])^(a[106] & b[96])^(a[105] & b[97])^(a[104] & b[98])^(a[103] & b[99])^(a[102] & b[100])^(a[101] & b[101])^(a[100] & b[102])^(a[99] & b[103])^(a[98] & b[104])^(a[97] & b[105])^(a[96] & b[106])^(a[95] & b[107])^(a[94] & b[108])^(a[93] & b[109])^(a[92] & b[110])^(a[91] & b[111])^(a[90] & b[112])^(a[89] & b[113])^(a[88] & b[114])^(a[87] & b[115])^(a[86] & b[116])^(a[85] & b[117])^(a[84] & b[118])^(a[83] & b[119])^(a[82] & b[120])^(a[81] & b[121])^(a[80] & b[122])^(a[79] & b[123])^(a[78] & b[124])^(a[77] & b[125])^(a[76] & b[126])^(a[75] & b[127])^(a[74] & b[128])^(a[73] & b[129])^(a[72] & b[130])^(a[71] & b[131])^(a[70] & b[132])^(a[69] & b[133])^(a[68] & b[134])^(a[67] & b[135])^(a[66] & b[136])^(a[65] & b[137])^(a[64] & b[138])^(a[63] & b[139])^(a[62] & b[140])^(a[61] & b[141])^(a[60] & b[142])^(a[59] & b[143])^(a[58] & b[144])^(a[57] & b[145])^(a[56] & b[146])^(a[55] & b[147])^(a[54] & b[148])^(a[53] & b[149])^(a[52] & b[150])^(a[51] & b[151])^(a[50] & b[152])^(a[49] & b[153])^(a[48] & b[154])^(a[47] & b[155])^(a[46] & b[156])^(a[45] & b[157])^(a[44] & b[158])^(a[43] & b[159])^(a[42] & b[160])^(a[41] & b[161])^(a[40] & b[162]);
assign y[203] = (a[162] & b[41])^(a[161] & b[42])^(a[160] & b[43])^(a[159] & b[44])^(a[158] & b[45])^(a[157] & b[46])^(a[156] & b[47])^(a[155] & b[48])^(a[154] & b[49])^(a[153] & b[50])^(a[152] & b[51])^(a[151] & b[52])^(a[150] & b[53])^(a[149] & b[54])^(a[148] & b[55])^(a[147] & b[56])^(a[146] & b[57])^(a[145] & b[58])^(a[144] & b[59])^(a[143] & b[60])^(a[142] & b[61])^(a[141] & b[62])^(a[140] & b[63])^(a[139] & b[64])^(a[138] & b[65])^(a[137] & b[66])^(a[136] & b[67])^(a[135] & b[68])^(a[134] & b[69])^(a[133] & b[70])^(a[132] & b[71])^(a[131] & b[72])^(a[130] & b[73])^(a[129] & b[74])^(a[128] & b[75])^(a[127] & b[76])^(a[126] & b[77])^(a[125] & b[78])^(a[124] & b[79])^(a[123] & b[80])^(a[122] & b[81])^(a[121] & b[82])^(a[120] & b[83])^(a[119] & b[84])^(a[118] & b[85])^(a[117] & b[86])^(a[116] & b[87])^(a[115] & b[88])^(a[114] & b[89])^(a[113] & b[90])^(a[112] & b[91])^(a[111] & b[92])^(a[110] & b[93])^(a[109] & b[94])^(a[108] & b[95])^(a[107] & b[96])^(a[106] & b[97])^(a[105] & b[98])^(a[104] & b[99])^(a[103] & b[100])^(a[102] & b[101])^(a[101] & b[102])^(a[100] & b[103])^(a[99] & b[104])^(a[98] & b[105])^(a[97] & b[106])^(a[96] & b[107])^(a[95] & b[108])^(a[94] & b[109])^(a[93] & b[110])^(a[92] & b[111])^(a[91] & b[112])^(a[90] & b[113])^(a[89] & b[114])^(a[88] & b[115])^(a[87] & b[116])^(a[86] & b[117])^(a[85] & b[118])^(a[84] & b[119])^(a[83] & b[120])^(a[82] & b[121])^(a[81] & b[122])^(a[80] & b[123])^(a[79] & b[124])^(a[78] & b[125])^(a[77] & b[126])^(a[76] & b[127])^(a[75] & b[128])^(a[74] & b[129])^(a[73] & b[130])^(a[72] & b[131])^(a[71] & b[132])^(a[70] & b[133])^(a[69] & b[134])^(a[68] & b[135])^(a[67] & b[136])^(a[66] & b[137])^(a[65] & b[138])^(a[64] & b[139])^(a[63] & b[140])^(a[62] & b[141])^(a[61] & b[142])^(a[60] & b[143])^(a[59] & b[144])^(a[58] & b[145])^(a[57] & b[146])^(a[56] & b[147])^(a[55] & b[148])^(a[54] & b[149])^(a[53] & b[150])^(a[52] & b[151])^(a[51] & b[152])^(a[50] & b[153])^(a[49] & b[154])^(a[48] & b[155])^(a[47] & b[156])^(a[46] & b[157])^(a[45] & b[158])^(a[44] & b[159])^(a[43] & b[160])^(a[42] & b[161])^(a[41] & b[162]);
assign y[204] = (a[162] & b[42])^(a[161] & b[43])^(a[160] & b[44])^(a[159] & b[45])^(a[158] & b[46])^(a[157] & b[47])^(a[156] & b[48])^(a[155] & b[49])^(a[154] & b[50])^(a[153] & b[51])^(a[152] & b[52])^(a[151] & b[53])^(a[150] & b[54])^(a[149] & b[55])^(a[148] & b[56])^(a[147] & b[57])^(a[146] & b[58])^(a[145] & b[59])^(a[144] & b[60])^(a[143] & b[61])^(a[142] & b[62])^(a[141] & b[63])^(a[140] & b[64])^(a[139] & b[65])^(a[138] & b[66])^(a[137] & b[67])^(a[136] & b[68])^(a[135] & b[69])^(a[134] & b[70])^(a[133] & b[71])^(a[132] & b[72])^(a[131] & b[73])^(a[130] & b[74])^(a[129] & b[75])^(a[128] & b[76])^(a[127] & b[77])^(a[126] & b[78])^(a[125] & b[79])^(a[124] & b[80])^(a[123] & b[81])^(a[122] & b[82])^(a[121] & b[83])^(a[120] & b[84])^(a[119] & b[85])^(a[118] & b[86])^(a[117] & b[87])^(a[116] & b[88])^(a[115] & b[89])^(a[114] & b[90])^(a[113] & b[91])^(a[112] & b[92])^(a[111] & b[93])^(a[110] & b[94])^(a[109] & b[95])^(a[108] & b[96])^(a[107] & b[97])^(a[106] & b[98])^(a[105] & b[99])^(a[104] & b[100])^(a[103] & b[101])^(a[102] & b[102])^(a[101] & b[103])^(a[100] & b[104])^(a[99] & b[105])^(a[98] & b[106])^(a[97] & b[107])^(a[96] & b[108])^(a[95] & b[109])^(a[94] & b[110])^(a[93] & b[111])^(a[92] & b[112])^(a[91] & b[113])^(a[90] & b[114])^(a[89] & b[115])^(a[88] & b[116])^(a[87] & b[117])^(a[86] & b[118])^(a[85] & b[119])^(a[84] & b[120])^(a[83] & b[121])^(a[82] & b[122])^(a[81] & b[123])^(a[80] & b[124])^(a[79] & b[125])^(a[78] & b[126])^(a[77] & b[127])^(a[76] & b[128])^(a[75] & b[129])^(a[74] & b[130])^(a[73] & b[131])^(a[72] & b[132])^(a[71] & b[133])^(a[70] & b[134])^(a[69] & b[135])^(a[68] & b[136])^(a[67] & b[137])^(a[66] & b[138])^(a[65] & b[139])^(a[64] & b[140])^(a[63] & b[141])^(a[62] & b[142])^(a[61] & b[143])^(a[60] & b[144])^(a[59] & b[145])^(a[58] & b[146])^(a[57] & b[147])^(a[56] & b[148])^(a[55] & b[149])^(a[54] & b[150])^(a[53] & b[151])^(a[52] & b[152])^(a[51] & b[153])^(a[50] & b[154])^(a[49] & b[155])^(a[48] & b[156])^(a[47] & b[157])^(a[46] & b[158])^(a[45] & b[159])^(a[44] & b[160])^(a[43] & b[161])^(a[42] & b[162]);
assign y[205] = (a[162] & b[43])^(a[161] & b[44])^(a[160] & b[45])^(a[159] & b[46])^(a[158] & b[47])^(a[157] & b[48])^(a[156] & b[49])^(a[155] & b[50])^(a[154] & b[51])^(a[153] & b[52])^(a[152] & b[53])^(a[151] & b[54])^(a[150] & b[55])^(a[149] & b[56])^(a[148] & b[57])^(a[147] & b[58])^(a[146] & b[59])^(a[145] & b[60])^(a[144] & b[61])^(a[143] & b[62])^(a[142] & b[63])^(a[141] & b[64])^(a[140] & b[65])^(a[139] & b[66])^(a[138] & b[67])^(a[137] & b[68])^(a[136] & b[69])^(a[135] & b[70])^(a[134] & b[71])^(a[133] & b[72])^(a[132] & b[73])^(a[131] & b[74])^(a[130] & b[75])^(a[129] & b[76])^(a[128] & b[77])^(a[127] & b[78])^(a[126] & b[79])^(a[125] & b[80])^(a[124] & b[81])^(a[123] & b[82])^(a[122] & b[83])^(a[121] & b[84])^(a[120] & b[85])^(a[119] & b[86])^(a[118] & b[87])^(a[117] & b[88])^(a[116] & b[89])^(a[115] & b[90])^(a[114] & b[91])^(a[113] & b[92])^(a[112] & b[93])^(a[111] & b[94])^(a[110] & b[95])^(a[109] & b[96])^(a[108] & b[97])^(a[107] & b[98])^(a[106] & b[99])^(a[105] & b[100])^(a[104] & b[101])^(a[103] & b[102])^(a[102] & b[103])^(a[101] & b[104])^(a[100] & b[105])^(a[99] & b[106])^(a[98] & b[107])^(a[97] & b[108])^(a[96] & b[109])^(a[95] & b[110])^(a[94] & b[111])^(a[93] & b[112])^(a[92] & b[113])^(a[91] & b[114])^(a[90] & b[115])^(a[89] & b[116])^(a[88] & b[117])^(a[87] & b[118])^(a[86] & b[119])^(a[85] & b[120])^(a[84] & b[121])^(a[83] & b[122])^(a[82] & b[123])^(a[81] & b[124])^(a[80] & b[125])^(a[79] & b[126])^(a[78] & b[127])^(a[77] & b[128])^(a[76] & b[129])^(a[75] & b[130])^(a[74] & b[131])^(a[73] & b[132])^(a[72] & b[133])^(a[71] & b[134])^(a[70] & b[135])^(a[69] & b[136])^(a[68] & b[137])^(a[67] & b[138])^(a[66] & b[139])^(a[65] & b[140])^(a[64] & b[141])^(a[63] & b[142])^(a[62] & b[143])^(a[61] & b[144])^(a[60] & b[145])^(a[59] & b[146])^(a[58] & b[147])^(a[57] & b[148])^(a[56] & b[149])^(a[55] & b[150])^(a[54] & b[151])^(a[53] & b[152])^(a[52] & b[153])^(a[51] & b[154])^(a[50] & b[155])^(a[49] & b[156])^(a[48] & b[157])^(a[47] & b[158])^(a[46] & b[159])^(a[45] & b[160])^(a[44] & b[161])^(a[43] & b[162]);
assign y[206] = (a[162] & b[44])^(a[161] & b[45])^(a[160] & b[46])^(a[159] & b[47])^(a[158] & b[48])^(a[157] & b[49])^(a[156] & b[50])^(a[155] & b[51])^(a[154] & b[52])^(a[153] & b[53])^(a[152] & b[54])^(a[151] & b[55])^(a[150] & b[56])^(a[149] & b[57])^(a[148] & b[58])^(a[147] & b[59])^(a[146] & b[60])^(a[145] & b[61])^(a[144] & b[62])^(a[143] & b[63])^(a[142] & b[64])^(a[141] & b[65])^(a[140] & b[66])^(a[139] & b[67])^(a[138] & b[68])^(a[137] & b[69])^(a[136] & b[70])^(a[135] & b[71])^(a[134] & b[72])^(a[133] & b[73])^(a[132] & b[74])^(a[131] & b[75])^(a[130] & b[76])^(a[129] & b[77])^(a[128] & b[78])^(a[127] & b[79])^(a[126] & b[80])^(a[125] & b[81])^(a[124] & b[82])^(a[123] & b[83])^(a[122] & b[84])^(a[121] & b[85])^(a[120] & b[86])^(a[119] & b[87])^(a[118] & b[88])^(a[117] & b[89])^(a[116] & b[90])^(a[115] & b[91])^(a[114] & b[92])^(a[113] & b[93])^(a[112] & b[94])^(a[111] & b[95])^(a[110] & b[96])^(a[109] & b[97])^(a[108] & b[98])^(a[107] & b[99])^(a[106] & b[100])^(a[105] & b[101])^(a[104] & b[102])^(a[103] & b[103])^(a[102] & b[104])^(a[101] & b[105])^(a[100] & b[106])^(a[99] & b[107])^(a[98] & b[108])^(a[97] & b[109])^(a[96] & b[110])^(a[95] & b[111])^(a[94] & b[112])^(a[93] & b[113])^(a[92] & b[114])^(a[91] & b[115])^(a[90] & b[116])^(a[89] & b[117])^(a[88] & b[118])^(a[87] & b[119])^(a[86] & b[120])^(a[85] & b[121])^(a[84] & b[122])^(a[83] & b[123])^(a[82] & b[124])^(a[81] & b[125])^(a[80] & b[126])^(a[79] & b[127])^(a[78] & b[128])^(a[77] & b[129])^(a[76] & b[130])^(a[75] & b[131])^(a[74] & b[132])^(a[73] & b[133])^(a[72] & b[134])^(a[71] & b[135])^(a[70] & b[136])^(a[69] & b[137])^(a[68] & b[138])^(a[67] & b[139])^(a[66] & b[140])^(a[65] & b[141])^(a[64] & b[142])^(a[63] & b[143])^(a[62] & b[144])^(a[61] & b[145])^(a[60] & b[146])^(a[59] & b[147])^(a[58] & b[148])^(a[57] & b[149])^(a[56] & b[150])^(a[55] & b[151])^(a[54] & b[152])^(a[53] & b[153])^(a[52] & b[154])^(a[51] & b[155])^(a[50] & b[156])^(a[49] & b[157])^(a[48] & b[158])^(a[47] & b[159])^(a[46] & b[160])^(a[45] & b[161])^(a[44] & b[162]);
assign y[207] = (a[162] & b[45])^(a[161] & b[46])^(a[160] & b[47])^(a[159] & b[48])^(a[158] & b[49])^(a[157] & b[50])^(a[156] & b[51])^(a[155] & b[52])^(a[154] & b[53])^(a[153] & b[54])^(a[152] & b[55])^(a[151] & b[56])^(a[150] & b[57])^(a[149] & b[58])^(a[148] & b[59])^(a[147] & b[60])^(a[146] & b[61])^(a[145] & b[62])^(a[144] & b[63])^(a[143] & b[64])^(a[142] & b[65])^(a[141] & b[66])^(a[140] & b[67])^(a[139] & b[68])^(a[138] & b[69])^(a[137] & b[70])^(a[136] & b[71])^(a[135] & b[72])^(a[134] & b[73])^(a[133] & b[74])^(a[132] & b[75])^(a[131] & b[76])^(a[130] & b[77])^(a[129] & b[78])^(a[128] & b[79])^(a[127] & b[80])^(a[126] & b[81])^(a[125] & b[82])^(a[124] & b[83])^(a[123] & b[84])^(a[122] & b[85])^(a[121] & b[86])^(a[120] & b[87])^(a[119] & b[88])^(a[118] & b[89])^(a[117] & b[90])^(a[116] & b[91])^(a[115] & b[92])^(a[114] & b[93])^(a[113] & b[94])^(a[112] & b[95])^(a[111] & b[96])^(a[110] & b[97])^(a[109] & b[98])^(a[108] & b[99])^(a[107] & b[100])^(a[106] & b[101])^(a[105] & b[102])^(a[104] & b[103])^(a[103] & b[104])^(a[102] & b[105])^(a[101] & b[106])^(a[100] & b[107])^(a[99] & b[108])^(a[98] & b[109])^(a[97] & b[110])^(a[96] & b[111])^(a[95] & b[112])^(a[94] & b[113])^(a[93] & b[114])^(a[92] & b[115])^(a[91] & b[116])^(a[90] & b[117])^(a[89] & b[118])^(a[88] & b[119])^(a[87] & b[120])^(a[86] & b[121])^(a[85] & b[122])^(a[84] & b[123])^(a[83] & b[124])^(a[82] & b[125])^(a[81] & b[126])^(a[80] & b[127])^(a[79] & b[128])^(a[78] & b[129])^(a[77] & b[130])^(a[76] & b[131])^(a[75] & b[132])^(a[74] & b[133])^(a[73] & b[134])^(a[72] & b[135])^(a[71] & b[136])^(a[70] & b[137])^(a[69] & b[138])^(a[68] & b[139])^(a[67] & b[140])^(a[66] & b[141])^(a[65] & b[142])^(a[64] & b[143])^(a[63] & b[144])^(a[62] & b[145])^(a[61] & b[146])^(a[60] & b[147])^(a[59] & b[148])^(a[58] & b[149])^(a[57] & b[150])^(a[56] & b[151])^(a[55] & b[152])^(a[54] & b[153])^(a[53] & b[154])^(a[52] & b[155])^(a[51] & b[156])^(a[50] & b[157])^(a[49] & b[158])^(a[48] & b[159])^(a[47] & b[160])^(a[46] & b[161])^(a[45] & b[162]);
assign y[208] = (a[162] & b[46])^(a[161] & b[47])^(a[160] & b[48])^(a[159] & b[49])^(a[158] & b[50])^(a[157] & b[51])^(a[156] & b[52])^(a[155] & b[53])^(a[154] & b[54])^(a[153] & b[55])^(a[152] & b[56])^(a[151] & b[57])^(a[150] & b[58])^(a[149] & b[59])^(a[148] & b[60])^(a[147] & b[61])^(a[146] & b[62])^(a[145] & b[63])^(a[144] & b[64])^(a[143] & b[65])^(a[142] & b[66])^(a[141] & b[67])^(a[140] & b[68])^(a[139] & b[69])^(a[138] & b[70])^(a[137] & b[71])^(a[136] & b[72])^(a[135] & b[73])^(a[134] & b[74])^(a[133] & b[75])^(a[132] & b[76])^(a[131] & b[77])^(a[130] & b[78])^(a[129] & b[79])^(a[128] & b[80])^(a[127] & b[81])^(a[126] & b[82])^(a[125] & b[83])^(a[124] & b[84])^(a[123] & b[85])^(a[122] & b[86])^(a[121] & b[87])^(a[120] & b[88])^(a[119] & b[89])^(a[118] & b[90])^(a[117] & b[91])^(a[116] & b[92])^(a[115] & b[93])^(a[114] & b[94])^(a[113] & b[95])^(a[112] & b[96])^(a[111] & b[97])^(a[110] & b[98])^(a[109] & b[99])^(a[108] & b[100])^(a[107] & b[101])^(a[106] & b[102])^(a[105] & b[103])^(a[104] & b[104])^(a[103] & b[105])^(a[102] & b[106])^(a[101] & b[107])^(a[100] & b[108])^(a[99] & b[109])^(a[98] & b[110])^(a[97] & b[111])^(a[96] & b[112])^(a[95] & b[113])^(a[94] & b[114])^(a[93] & b[115])^(a[92] & b[116])^(a[91] & b[117])^(a[90] & b[118])^(a[89] & b[119])^(a[88] & b[120])^(a[87] & b[121])^(a[86] & b[122])^(a[85] & b[123])^(a[84] & b[124])^(a[83] & b[125])^(a[82] & b[126])^(a[81] & b[127])^(a[80] & b[128])^(a[79] & b[129])^(a[78] & b[130])^(a[77] & b[131])^(a[76] & b[132])^(a[75] & b[133])^(a[74] & b[134])^(a[73] & b[135])^(a[72] & b[136])^(a[71] & b[137])^(a[70] & b[138])^(a[69] & b[139])^(a[68] & b[140])^(a[67] & b[141])^(a[66] & b[142])^(a[65] & b[143])^(a[64] & b[144])^(a[63] & b[145])^(a[62] & b[146])^(a[61] & b[147])^(a[60] & b[148])^(a[59] & b[149])^(a[58] & b[150])^(a[57] & b[151])^(a[56] & b[152])^(a[55] & b[153])^(a[54] & b[154])^(a[53] & b[155])^(a[52] & b[156])^(a[51] & b[157])^(a[50] & b[158])^(a[49] & b[159])^(a[48] & b[160])^(a[47] & b[161])^(a[46] & b[162]);
assign y[209] = (a[162] & b[47])^(a[161] & b[48])^(a[160] & b[49])^(a[159] & b[50])^(a[158] & b[51])^(a[157] & b[52])^(a[156] & b[53])^(a[155] & b[54])^(a[154] & b[55])^(a[153] & b[56])^(a[152] & b[57])^(a[151] & b[58])^(a[150] & b[59])^(a[149] & b[60])^(a[148] & b[61])^(a[147] & b[62])^(a[146] & b[63])^(a[145] & b[64])^(a[144] & b[65])^(a[143] & b[66])^(a[142] & b[67])^(a[141] & b[68])^(a[140] & b[69])^(a[139] & b[70])^(a[138] & b[71])^(a[137] & b[72])^(a[136] & b[73])^(a[135] & b[74])^(a[134] & b[75])^(a[133] & b[76])^(a[132] & b[77])^(a[131] & b[78])^(a[130] & b[79])^(a[129] & b[80])^(a[128] & b[81])^(a[127] & b[82])^(a[126] & b[83])^(a[125] & b[84])^(a[124] & b[85])^(a[123] & b[86])^(a[122] & b[87])^(a[121] & b[88])^(a[120] & b[89])^(a[119] & b[90])^(a[118] & b[91])^(a[117] & b[92])^(a[116] & b[93])^(a[115] & b[94])^(a[114] & b[95])^(a[113] & b[96])^(a[112] & b[97])^(a[111] & b[98])^(a[110] & b[99])^(a[109] & b[100])^(a[108] & b[101])^(a[107] & b[102])^(a[106] & b[103])^(a[105] & b[104])^(a[104] & b[105])^(a[103] & b[106])^(a[102] & b[107])^(a[101] & b[108])^(a[100] & b[109])^(a[99] & b[110])^(a[98] & b[111])^(a[97] & b[112])^(a[96] & b[113])^(a[95] & b[114])^(a[94] & b[115])^(a[93] & b[116])^(a[92] & b[117])^(a[91] & b[118])^(a[90] & b[119])^(a[89] & b[120])^(a[88] & b[121])^(a[87] & b[122])^(a[86] & b[123])^(a[85] & b[124])^(a[84] & b[125])^(a[83] & b[126])^(a[82] & b[127])^(a[81] & b[128])^(a[80] & b[129])^(a[79] & b[130])^(a[78] & b[131])^(a[77] & b[132])^(a[76] & b[133])^(a[75] & b[134])^(a[74] & b[135])^(a[73] & b[136])^(a[72] & b[137])^(a[71] & b[138])^(a[70] & b[139])^(a[69] & b[140])^(a[68] & b[141])^(a[67] & b[142])^(a[66] & b[143])^(a[65] & b[144])^(a[64] & b[145])^(a[63] & b[146])^(a[62] & b[147])^(a[61] & b[148])^(a[60] & b[149])^(a[59] & b[150])^(a[58] & b[151])^(a[57] & b[152])^(a[56] & b[153])^(a[55] & b[154])^(a[54] & b[155])^(a[53] & b[156])^(a[52] & b[157])^(a[51] & b[158])^(a[50] & b[159])^(a[49] & b[160])^(a[48] & b[161])^(a[47] & b[162]);
assign y[210] = (a[162] & b[48])^(a[161] & b[49])^(a[160] & b[50])^(a[159] & b[51])^(a[158] & b[52])^(a[157] & b[53])^(a[156] & b[54])^(a[155] & b[55])^(a[154] & b[56])^(a[153] & b[57])^(a[152] & b[58])^(a[151] & b[59])^(a[150] & b[60])^(a[149] & b[61])^(a[148] & b[62])^(a[147] & b[63])^(a[146] & b[64])^(a[145] & b[65])^(a[144] & b[66])^(a[143] & b[67])^(a[142] & b[68])^(a[141] & b[69])^(a[140] & b[70])^(a[139] & b[71])^(a[138] & b[72])^(a[137] & b[73])^(a[136] & b[74])^(a[135] & b[75])^(a[134] & b[76])^(a[133] & b[77])^(a[132] & b[78])^(a[131] & b[79])^(a[130] & b[80])^(a[129] & b[81])^(a[128] & b[82])^(a[127] & b[83])^(a[126] & b[84])^(a[125] & b[85])^(a[124] & b[86])^(a[123] & b[87])^(a[122] & b[88])^(a[121] & b[89])^(a[120] & b[90])^(a[119] & b[91])^(a[118] & b[92])^(a[117] & b[93])^(a[116] & b[94])^(a[115] & b[95])^(a[114] & b[96])^(a[113] & b[97])^(a[112] & b[98])^(a[111] & b[99])^(a[110] & b[100])^(a[109] & b[101])^(a[108] & b[102])^(a[107] & b[103])^(a[106] & b[104])^(a[105] & b[105])^(a[104] & b[106])^(a[103] & b[107])^(a[102] & b[108])^(a[101] & b[109])^(a[100] & b[110])^(a[99] & b[111])^(a[98] & b[112])^(a[97] & b[113])^(a[96] & b[114])^(a[95] & b[115])^(a[94] & b[116])^(a[93] & b[117])^(a[92] & b[118])^(a[91] & b[119])^(a[90] & b[120])^(a[89] & b[121])^(a[88] & b[122])^(a[87] & b[123])^(a[86] & b[124])^(a[85] & b[125])^(a[84] & b[126])^(a[83] & b[127])^(a[82] & b[128])^(a[81] & b[129])^(a[80] & b[130])^(a[79] & b[131])^(a[78] & b[132])^(a[77] & b[133])^(a[76] & b[134])^(a[75] & b[135])^(a[74] & b[136])^(a[73] & b[137])^(a[72] & b[138])^(a[71] & b[139])^(a[70] & b[140])^(a[69] & b[141])^(a[68] & b[142])^(a[67] & b[143])^(a[66] & b[144])^(a[65] & b[145])^(a[64] & b[146])^(a[63] & b[147])^(a[62] & b[148])^(a[61] & b[149])^(a[60] & b[150])^(a[59] & b[151])^(a[58] & b[152])^(a[57] & b[153])^(a[56] & b[154])^(a[55] & b[155])^(a[54] & b[156])^(a[53] & b[157])^(a[52] & b[158])^(a[51] & b[159])^(a[50] & b[160])^(a[49] & b[161])^(a[48] & b[162]);
assign y[211] = (a[162] & b[49])^(a[161] & b[50])^(a[160] & b[51])^(a[159] & b[52])^(a[158] & b[53])^(a[157] & b[54])^(a[156] & b[55])^(a[155] & b[56])^(a[154] & b[57])^(a[153] & b[58])^(a[152] & b[59])^(a[151] & b[60])^(a[150] & b[61])^(a[149] & b[62])^(a[148] & b[63])^(a[147] & b[64])^(a[146] & b[65])^(a[145] & b[66])^(a[144] & b[67])^(a[143] & b[68])^(a[142] & b[69])^(a[141] & b[70])^(a[140] & b[71])^(a[139] & b[72])^(a[138] & b[73])^(a[137] & b[74])^(a[136] & b[75])^(a[135] & b[76])^(a[134] & b[77])^(a[133] & b[78])^(a[132] & b[79])^(a[131] & b[80])^(a[130] & b[81])^(a[129] & b[82])^(a[128] & b[83])^(a[127] & b[84])^(a[126] & b[85])^(a[125] & b[86])^(a[124] & b[87])^(a[123] & b[88])^(a[122] & b[89])^(a[121] & b[90])^(a[120] & b[91])^(a[119] & b[92])^(a[118] & b[93])^(a[117] & b[94])^(a[116] & b[95])^(a[115] & b[96])^(a[114] & b[97])^(a[113] & b[98])^(a[112] & b[99])^(a[111] & b[100])^(a[110] & b[101])^(a[109] & b[102])^(a[108] & b[103])^(a[107] & b[104])^(a[106] & b[105])^(a[105] & b[106])^(a[104] & b[107])^(a[103] & b[108])^(a[102] & b[109])^(a[101] & b[110])^(a[100] & b[111])^(a[99] & b[112])^(a[98] & b[113])^(a[97] & b[114])^(a[96] & b[115])^(a[95] & b[116])^(a[94] & b[117])^(a[93] & b[118])^(a[92] & b[119])^(a[91] & b[120])^(a[90] & b[121])^(a[89] & b[122])^(a[88] & b[123])^(a[87] & b[124])^(a[86] & b[125])^(a[85] & b[126])^(a[84] & b[127])^(a[83] & b[128])^(a[82] & b[129])^(a[81] & b[130])^(a[80] & b[131])^(a[79] & b[132])^(a[78] & b[133])^(a[77] & b[134])^(a[76] & b[135])^(a[75] & b[136])^(a[74] & b[137])^(a[73] & b[138])^(a[72] & b[139])^(a[71] & b[140])^(a[70] & b[141])^(a[69] & b[142])^(a[68] & b[143])^(a[67] & b[144])^(a[66] & b[145])^(a[65] & b[146])^(a[64] & b[147])^(a[63] & b[148])^(a[62] & b[149])^(a[61] & b[150])^(a[60] & b[151])^(a[59] & b[152])^(a[58] & b[153])^(a[57] & b[154])^(a[56] & b[155])^(a[55] & b[156])^(a[54] & b[157])^(a[53] & b[158])^(a[52] & b[159])^(a[51] & b[160])^(a[50] & b[161])^(a[49] & b[162]);
assign y[212] = (a[162] & b[50])^(a[161] & b[51])^(a[160] & b[52])^(a[159] & b[53])^(a[158] & b[54])^(a[157] & b[55])^(a[156] & b[56])^(a[155] & b[57])^(a[154] & b[58])^(a[153] & b[59])^(a[152] & b[60])^(a[151] & b[61])^(a[150] & b[62])^(a[149] & b[63])^(a[148] & b[64])^(a[147] & b[65])^(a[146] & b[66])^(a[145] & b[67])^(a[144] & b[68])^(a[143] & b[69])^(a[142] & b[70])^(a[141] & b[71])^(a[140] & b[72])^(a[139] & b[73])^(a[138] & b[74])^(a[137] & b[75])^(a[136] & b[76])^(a[135] & b[77])^(a[134] & b[78])^(a[133] & b[79])^(a[132] & b[80])^(a[131] & b[81])^(a[130] & b[82])^(a[129] & b[83])^(a[128] & b[84])^(a[127] & b[85])^(a[126] & b[86])^(a[125] & b[87])^(a[124] & b[88])^(a[123] & b[89])^(a[122] & b[90])^(a[121] & b[91])^(a[120] & b[92])^(a[119] & b[93])^(a[118] & b[94])^(a[117] & b[95])^(a[116] & b[96])^(a[115] & b[97])^(a[114] & b[98])^(a[113] & b[99])^(a[112] & b[100])^(a[111] & b[101])^(a[110] & b[102])^(a[109] & b[103])^(a[108] & b[104])^(a[107] & b[105])^(a[106] & b[106])^(a[105] & b[107])^(a[104] & b[108])^(a[103] & b[109])^(a[102] & b[110])^(a[101] & b[111])^(a[100] & b[112])^(a[99] & b[113])^(a[98] & b[114])^(a[97] & b[115])^(a[96] & b[116])^(a[95] & b[117])^(a[94] & b[118])^(a[93] & b[119])^(a[92] & b[120])^(a[91] & b[121])^(a[90] & b[122])^(a[89] & b[123])^(a[88] & b[124])^(a[87] & b[125])^(a[86] & b[126])^(a[85] & b[127])^(a[84] & b[128])^(a[83] & b[129])^(a[82] & b[130])^(a[81] & b[131])^(a[80] & b[132])^(a[79] & b[133])^(a[78] & b[134])^(a[77] & b[135])^(a[76] & b[136])^(a[75] & b[137])^(a[74] & b[138])^(a[73] & b[139])^(a[72] & b[140])^(a[71] & b[141])^(a[70] & b[142])^(a[69] & b[143])^(a[68] & b[144])^(a[67] & b[145])^(a[66] & b[146])^(a[65] & b[147])^(a[64] & b[148])^(a[63] & b[149])^(a[62] & b[150])^(a[61] & b[151])^(a[60] & b[152])^(a[59] & b[153])^(a[58] & b[154])^(a[57] & b[155])^(a[56] & b[156])^(a[55] & b[157])^(a[54] & b[158])^(a[53] & b[159])^(a[52] & b[160])^(a[51] & b[161])^(a[50] & b[162]);
assign y[213] = (a[162] & b[51])^(a[161] & b[52])^(a[160] & b[53])^(a[159] & b[54])^(a[158] & b[55])^(a[157] & b[56])^(a[156] & b[57])^(a[155] & b[58])^(a[154] & b[59])^(a[153] & b[60])^(a[152] & b[61])^(a[151] & b[62])^(a[150] & b[63])^(a[149] & b[64])^(a[148] & b[65])^(a[147] & b[66])^(a[146] & b[67])^(a[145] & b[68])^(a[144] & b[69])^(a[143] & b[70])^(a[142] & b[71])^(a[141] & b[72])^(a[140] & b[73])^(a[139] & b[74])^(a[138] & b[75])^(a[137] & b[76])^(a[136] & b[77])^(a[135] & b[78])^(a[134] & b[79])^(a[133] & b[80])^(a[132] & b[81])^(a[131] & b[82])^(a[130] & b[83])^(a[129] & b[84])^(a[128] & b[85])^(a[127] & b[86])^(a[126] & b[87])^(a[125] & b[88])^(a[124] & b[89])^(a[123] & b[90])^(a[122] & b[91])^(a[121] & b[92])^(a[120] & b[93])^(a[119] & b[94])^(a[118] & b[95])^(a[117] & b[96])^(a[116] & b[97])^(a[115] & b[98])^(a[114] & b[99])^(a[113] & b[100])^(a[112] & b[101])^(a[111] & b[102])^(a[110] & b[103])^(a[109] & b[104])^(a[108] & b[105])^(a[107] & b[106])^(a[106] & b[107])^(a[105] & b[108])^(a[104] & b[109])^(a[103] & b[110])^(a[102] & b[111])^(a[101] & b[112])^(a[100] & b[113])^(a[99] & b[114])^(a[98] & b[115])^(a[97] & b[116])^(a[96] & b[117])^(a[95] & b[118])^(a[94] & b[119])^(a[93] & b[120])^(a[92] & b[121])^(a[91] & b[122])^(a[90] & b[123])^(a[89] & b[124])^(a[88] & b[125])^(a[87] & b[126])^(a[86] & b[127])^(a[85] & b[128])^(a[84] & b[129])^(a[83] & b[130])^(a[82] & b[131])^(a[81] & b[132])^(a[80] & b[133])^(a[79] & b[134])^(a[78] & b[135])^(a[77] & b[136])^(a[76] & b[137])^(a[75] & b[138])^(a[74] & b[139])^(a[73] & b[140])^(a[72] & b[141])^(a[71] & b[142])^(a[70] & b[143])^(a[69] & b[144])^(a[68] & b[145])^(a[67] & b[146])^(a[66] & b[147])^(a[65] & b[148])^(a[64] & b[149])^(a[63] & b[150])^(a[62] & b[151])^(a[61] & b[152])^(a[60] & b[153])^(a[59] & b[154])^(a[58] & b[155])^(a[57] & b[156])^(a[56] & b[157])^(a[55] & b[158])^(a[54] & b[159])^(a[53] & b[160])^(a[52] & b[161])^(a[51] & b[162]);
assign y[214] = (a[162] & b[52])^(a[161] & b[53])^(a[160] & b[54])^(a[159] & b[55])^(a[158] & b[56])^(a[157] & b[57])^(a[156] & b[58])^(a[155] & b[59])^(a[154] & b[60])^(a[153] & b[61])^(a[152] & b[62])^(a[151] & b[63])^(a[150] & b[64])^(a[149] & b[65])^(a[148] & b[66])^(a[147] & b[67])^(a[146] & b[68])^(a[145] & b[69])^(a[144] & b[70])^(a[143] & b[71])^(a[142] & b[72])^(a[141] & b[73])^(a[140] & b[74])^(a[139] & b[75])^(a[138] & b[76])^(a[137] & b[77])^(a[136] & b[78])^(a[135] & b[79])^(a[134] & b[80])^(a[133] & b[81])^(a[132] & b[82])^(a[131] & b[83])^(a[130] & b[84])^(a[129] & b[85])^(a[128] & b[86])^(a[127] & b[87])^(a[126] & b[88])^(a[125] & b[89])^(a[124] & b[90])^(a[123] & b[91])^(a[122] & b[92])^(a[121] & b[93])^(a[120] & b[94])^(a[119] & b[95])^(a[118] & b[96])^(a[117] & b[97])^(a[116] & b[98])^(a[115] & b[99])^(a[114] & b[100])^(a[113] & b[101])^(a[112] & b[102])^(a[111] & b[103])^(a[110] & b[104])^(a[109] & b[105])^(a[108] & b[106])^(a[107] & b[107])^(a[106] & b[108])^(a[105] & b[109])^(a[104] & b[110])^(a[103] & b[111])^(a[102] & b[112])^(a[101] & b[113])^(a[100] & b[114])^(a[99] & b[115])^(a[98] & b[116])^(a[97] & b[117])^(a[96] & b[118])^(a[95] & b[119])^(a[94] & b[120])^(a[93] & b[121])^(a[92] & b[122])^(a[91] & b[123])^(a[90] & b[124])^(a[89] & b[125])^(a[88] & b[126])^(a[87] & b[127])^(a[86] & b[128])^(a[85] & b[129])^(a[84] & b[130])^(a[83] & b[131])^(a[82] & b[132])^(a[81] & b[133])^(a[80] & b[134])^(a[79] & b[135])^(a[78] & b[136])^(a[77] & b[137])^(a[76] & b[138])^(a[75] & b[139])^(a[74] & b[140])^(a[73] & b[141])^(a[72] & b[142])^(a[71] & b[143])^(a[70] & b[144])^(a[69] & b[145])^(a[68] & b[146])^(a[67] & b[147])^(a[66] & b[148])^(a[65] & b[149])^(a[64] & b[150])^(a[63] & b[151])^(a[62] & b[152])^(a[61] & b[153])^(a[60] & b[154])^(a[59] & b[155])^(a[58] & b[156])^(a[57] & b[157])^(a[56] & b[158])^(a[55] & b[159])^(a[54] & b[160])^(a[53] & b[161])^(a[52] & b[162]);
assign y[215] = (a[162] & b[53])^(a[161] & b[54])^(a[160] & b[55])^(a[159] & b[56])^(a[158] & b[57])^(a[157] & b[58])^(a[156] & b[59])^(a[155] & b[60])^(a[154] & b[61])^(a[153] & b[62])^(a[152] & b[63])^(a[151] & b[64])^(a[150] & b[65])^(a[149] & b[66])^(a[148] & b[67])^(a[147] & b[68])^(a[146] & b[69])^(a[145] & b[70])^(a[144] & b[71])^(a[143] & b[72])^(a[142] & b[73])^(a[141] & b[74])^(a[140] & b[75])^(a[139] & b[76])^(a[138] & b[77])^(a[137] & b[78])^(a[136] & b[79])^(a[135] & b[80])^(a[134] & b[81])^(a[133] & b[82])^(a[132] & b[83])^(a[131] & b[84])^(a[130] & b[85])^(a[129] & b[86])^(a[128] & b[87])^(a[127] & b[88])^(a[126] & b[89])^(a[125] & b[90])^(a[124] & b[91])^(a[123] & b[92])^(a[122] & b[93])^(a[121] & b[94])^(a[120] & b[95])^(a[119] & b[96])^(a[118] & b[97])^(a[117] & b[98])^(a[116] & b[99])^(a[115] & b[100])^(a[114] & b[101])^(a[113] & b[102])^(a[112] & b[103])^(a[111] & b[104])^(a[110] & b[105])^(a[109] & b[106])^(a[108] & b[107])^(a[107] & b[108])^(a[106] & b[109])^(a[105] & b[110])^(a[104] & b[111])^(a[103] & b[112])^(a[102] & b[113])^(a[101] & b[114])^(a[100] & b[115])^(a[99] & b[116])^(a[98] & b[117])^(a[97] & b[118])^(a[96] & b[119])^(a[95] & b[120])^(a[94] & b[121])^(a[93] & b[122])^(a[92] & b[123])^(a[91] & b[124])^(a[90] & b[125])^(a[89] & b[126])^(a[88] & b[127])^(a[87] & b[128])^(a[86] & b[129])^(a[85] & b[130])^(a[84] & b[131])^(a[83] & b[132])^(a[82] & b[133])^(a[81] & b[134])^(a[80] & b[135])^(a[79] & b[136])^(a[78] & b[137])^(a[77] & b[138])^(a[76] & b[139])^(a[75] & b[140])^(a[74] & b[141])^(a[73] & b[142])^(a[72] & b[143])^(a[71] & b[144])^(a[70] & b[145])^(a[69] & b[146])^(a[68] & b[147])^(a[67] & b[148])^(a[66] & b[149])^(a[65] & b[150])^(a[64] & b[151])^(a[63] & b[152])^(a[62] & b[153])^(a[61] & b[154])^(a[60] & b[155])^(a[59] & b[156])^(a[58] & b[157])^(a[57] & b[158])^(a[56] & b[159])^(a[55] & b[160])^(a[54] & b[161])^(a[53] & b[162]);
assign y[216] = (a[162] & b[54])^(a[161] & b[55])^(a[160] & b[56])^(a[159] & b[57])^(a[158] & b[58])^(a[157] & b[59])^(a[156] & b[60])^(a[155] & b[61])^(a[154] & b[62])^(a[153] & b[63])^(a[152] & b[64])^(a[151] & b[65])^(a[150] & b[66])^(a[149] & b[67])^(a[148] & b[68])^(a[147] & b[69])^(a[146] & b[70])^(a[145] & b[71])^(a[144] & b[72])^(a[143] & b[73])^(a[142] & b[74])^(a[141] & b[75])^(a[140] & b[76])^(a[139] & b[77])^(a[138] & b[78])^(a[137] & b[79])^(a[136] & b[80])^(a[135] & b[81])^(a[134] & b[82])^(a[133] & b[83])^(a[132] & b[84])^(a[131] & b[85])^(a[130] & b[86])^(a[129] & b[87])^(a[128] & b[88])^(a[127] & b[89])^(a[126] & b[90])^(a[125] & b[91])^(a[124] & b[92])^(a[123] & b[93])^(a[122] & b[94])^(a[121] & b[95])^(a[120] & b[96])^(a[119] & b[97])^(a[118] & b[98])^(a[117] & b[99])^(a[116] & b[100])^(a[115] & b[101])^(a[114] & b[102])^(a[113] & b[103])^(a[112] & b[104])^(a[111] & b[105])^(a[110] & b[106])^(a[109] & b[107])^(a[108] & b[108])^(a[107] & b[109])^(a[106] & b[110])^(a[105] & b[111])^(a[104] & b[112])^(a[103] & b[113])^(a[102] & b[114])^(a[101] & b[115])^(a[100] & b[116])^(a[99] & b[117])^(a[98] & b[118])^(a[97] & b[119])^(a[96] & b[120])^(a[95] & b[121])^(a[94] & b[122])^(a[93] & b[123])^(a[92] & b[124])^(a[91] & b[125])^(a[90] & b[126])^(a[89] & b[127])^(a[88] & b[128])^(a[87] & b[129])^(a[86] & b[130])^(a[85] & b[131])^(a[84] & b[132])^(a[83] & b[133])^(a[82] & b[134])^(a[81] & b[135])^(a[80] & b[136])^(a[79] & b[137])^(a[78] & b[138])^(a[77] & b[139])^(a[76] & b[140])^(a[75] & b[141])^(a[74] & b[142])^(a[73] & b[143])^(a[72] & b[144])^(a[71] & b[145])^(a[70] & b[146])^(a[69] & b[147])^(a[68] & b[148])^(a[67] & b[149])^(a[66] & b[150])^(a[65] & b[151])^(a[64] & b[152])^(a[63] & b[153])^(a[62] & b[154])^(a[61] & b[155])^(a[60] & b[156])^(a[59] & b[157])^(a[58] & b[158])^(a[57] & b[159])^(a[56] & b[160])^(a[55] & b[161])^(a[54] & b[162]);
assign y[217] = (a[162] & b[55])^(a[161] & b[56])^(a[160] & b[57])^(a[159] & b[58])^(a[158] & b[59])^(a[157] & b[60])^(a[156] & b[61])^(a[155] & b[62])^(a[154] & b[63])^(a[153] & b[64])^(a[152] & b[65])^(a[151] & b[66])^(a[150] & b[67])^(a[149] & b[68])^(a[148] & b[69])^(a[147] & b[70])^(a[146] & b[71])^(a[145] & b[72])^(a[144] & b[73])^(a[143] & b[74])^(a[142] & b[75])^(a[141] & b[76])^(a[140] & b[77])^(a[139] & b[78])^(a[138] & b[79])^(a[137] & b[80])^(a[136] & b[81])^(a[135] & b[82])^(a[134] & b[83])^(a[133] & b[84])^(a[132] & b[85])^(a[131] & b[86])^(a[130] & b[87])^(a[129] & b[88])^(a[128] & b[89])^(a[127] & b[90])^(a[126] & b[91])^(a[125] & b[92])^(a[124] & b[93])^(a[123] & b[94])^(a[122] & b[95])^(a[121] & b[96])^(a[120] & b[97])^(a[119] & b[98])^(a[118] & b[99])^(a[117] & b[100])^(a[116] & b[101])^(a[115] & b[102])^(a[114] & b[103])^(a[113] & b[104])^(a[112] & b[105])^(a[111] & b[106])^(a[110] & b[107])^(a[109] & b[108])^(a[108] & b[109])^(a[107] & b[110])^(a[106] & b[111])^(a[105] & b[112])^(a[104] & b[113])^(a[103] & b[114])^(a[102] & b[115])^(a[101] & b[116])^(a[100] & b[117])^(a[99] & b[118])^(a[98] & b[119])^(a[97] & b[120])^(a[96] & b[121])^(a[95] & b[122])^(a[94] & b[123])^(a[93] & b[124])^(a[92] & b[125])^(a[91] & b[126])^(a[90] & b[127])^(a[89] & b[128])^(a[88] & b[129])^(a[87] & b[130])^(a[86] & b[131])^(a[85] & b[132])^(a[84] & b[133])^(a[83] & b[134])^(a[82] & b[135])^(a[81] & b[136])^(a[80] & b[137])^(a[79] & b[138])^(a[78] & b[139])^(a[77] & b[140])^(a[76] & b[141])^(a[75] & b[142])^(a[74] & b[143])^(a[73] & b[144])^(a[72] & b[145])^(a[71] & b[146])^(a[70] & b[147])^(a[69] & b[148])^(a[68] & b[149])^(a[67] & b[150])^(a[66] & b[151])^(a[65] & b[152])^(a[64] & b[153])^(a[63] & b[154])^(a[62] & b[155])^(a[61] & b[156])^(a[60] & b[157])^(a[59] & b[158])^(a[58] & b[159])^(a[57] & b[160])^(a[56] & b[161])^(a[55] & b[162]);
assign y[218] = (a[162] & b[56])^(a[161] & b[57])^(a[160] & b[58])^(a[159] & b[59])^(a[158] & b[60])^(a[157] & b[61])^(a[156] & b[62])^(a[155] & b[63])^(a[154] & b[64])^(a[153] & b[65])^(a[152] & b[66])^(a[151] & b[67])^(a[150] & b[68])^(a[149] & b[69])^(a[148] & b[70])^(a[147] & b[71])^(a[146] & b[72])^(a[145] & b[73])^(a[144] & b[74])^(a[143] & b[75])^(a[142] & b[76])^(a[141] & b[77])^(a[140] & b[78])^(a[139] & b[79])^(a[138] & b[80])^(a[137] & b[81])^(a[136] & b[82])^(a[135] & b[83])^(a[134] & b[84])^(a[133] & b[85])^(a[132] & b[86])^(a[131] & b[87])^(a[130] & b[88])^(a[129] & b[89])^(a[128] & b[90])^(a[127] & b[91])^(a[126] & b[92])^(a[125] & b[93])^(a[124] & b[94])^(a[123] & b[95])^(a[122] & b[96])^(a[121] & b[97])^(a[120] & b[98])^(a[119] & b[99])^(a[118] & b[100])^(a[117] & b[101])^(a[116] & b[102])^(a[115] & b[103])^(a[114] & b[104])^(a[113] & b[105])^(a[112] & b[106])^(a[111] & b[107])^(a[110] & b[108])^(a[109] & b[109])^(a[108] & b[110])^(a[107] & b[111])^(a[106] & b[112])^(a[105] & b[113])^(a[104] & b[114])^(a[103] & b[115])^(a[102] & b[116])^(a[101] & b[117])^(a[100] & b[118])^(a[99] & b[119])^(a[98] & b[120])^(a[97] & b[121])^(a[96] & b[122])^(a[95] & b[123])^(a[94] & b[124])^(a[93] & b[125])^(a[92] & b[126])^(a[91] & b[127])^(a[90] & b[128])^(a[89] & b[129])^(a[88] & b[130])^(a[87] & b[131])^(a[86] & b[132])^(a[85] & b[133])^(a[84] & b[134])^(a[83] & b[135])^(a[82] & b[136])^(a[81] & b[137])^(a[80] & b[138])^(a[79] & b[139])^(a[78] & b[140])^(a[77] & b[141])^(a[76] & b[142])^(a[75] & b[143])^(a[74] & b[144])^(a[73] & b[145])^(a[72] & b[146])^(a[71] & b[147])^(a[70] & b[148])^(a[69] & b[149])^(a[68] & b[150])^(a[67] & b[151])^(a[66] & b[152])^(a[65] & b[153])^(a[64] & b[154])^(a[63] & b[155])^(a[62] & b[156])^(a[61] & b[157])^(a[60] & b[158])^(a[59] & b[159])^(a[58] & b[160])^(a[57] & b[161])^(a[56] & b[162]);
assign y[219] = (a[162] & b[57])^(a[161] & b[58])^(a[160] & b[59])^(a[159] & b[60])^(a[158] & b[61])^(a[157] & b[62])^(a[156] & b[63])^(a[155] & b[64])^(a[154] & b[65])^(a[153] & b[66])^(a[152] & b[67])^(a[151] & b[68])^(a[150] & b[69])^(a[149] & b[70])^(a[148] & b[71])^(a[147] & b[72])^(a[146] & b[73])^(a[145] & b[74])^(a[144] & b[75])^(a[143] & b[76])^(a[142] & b[77])^(a[141] & b[78])^(a[140] & b[79])^(a[139] & b[80])^(a[138] & b[81])^(a[137] & b[82])^(a[136] & b[83])^(a[135] & b[84])^(a[134] & b[85])^(a[133] & b[86])^(a[132] & b[87])^(a[131] & b[88])^(a[130] & b[89])^(a[129] & b[90])^(a[128] & b[91])^(a[127] & b[92])^(a[126] & b[93])^(a[125] & b[94])^(a[124] & b[95])^(a[123] & b[96])^(a[122] & b[97])^(a[121] & b[98])^(a[120] & b[99])^(a[119] & b[100])^(a[118] & b[101])^(a[117] & b[102])^(a[116] & b[103])^(a[115] & b[104])^(a[114] & b[105])^(a[113] & b[106])^(a[112] & b[107])^(a[111] & b[108])^(a[110] & b[109])^(a[109] & b[110])^(a[108] & b[111])^(a[107] & b[112])^(a[106] & b[113])^(a[105] & b[114])^(a[104] & b[115])^(a[103] & b[116])^(a[102] & b[117])^(a[101] & b[118])^(a[100] & b[119])^(a[99] & b[120])^(a[98] & b[121])^(a[97] & b[122])^(a[96] & b[123])^(a[95] & b[124])^(a[94] & b[125])^(a[93] & b[126])^(a[92] & b[127])^(a[91] & b[128])^(a[90] & b[129])^(a[89] & b[130])^(a[88] & b[131])^(a[87] & b[132])^(a[86] & b[133])^(a[85] & b[134])^(a[84] & b[135])^(a[83] & b[136])^(a[82] & b[137])^(a[81] & b[138])^(a[80] & b[139])^(a[79] & b[140])^(a[78] & b[141])^(a[77] & b[142])^(a[76] & b[143])^(a[75] & b[144])^(a[74] & b[145])^(a[73] & b[146])^(a[72] & b[147])^(a[71] & b[148])^(a[70] & b[149])^(a[69] & b[150])^(a[68] & b[151])^(a[67] & b[152])^(a[66] & b[153])^(a[65] & b[154])^(a[64] & b[155])^(a[63] & b[156])^(a[62] & b[157])^(a[61] & b[158])^(a[60] & b[159])^(a[59] & b[160])^(a[58] & b[161])^(a[57] & b[162]);
assign y[220] = (a[162] & b[58])^(a[161] & b[59])^(a[160] & b[60])^(a[159] & b[61])^(a[158] & b[62])^(a[157] & b[63])^(a[156] & b[64])^(a[155] & b[65])^(a[154] & b[66])^(a[153] & b[67])^(a[152] & b[68])^(a[151] & b[69])^(a[150] & b[70])^(a[149] & b[71])^(a[148] & b[72])^(a[147] & b[73])^(a[146] & b[74])^(a[145] & b[75])^(a[144] & b[76])^(a[143] & b[77])^(a[142] & b[78])^(a[141] & b[79])^(a[140] & b[80])^(a[139] & b[81])^(a[138] & b[82])^(a[137] & b[83])^(a[136] & b[84])^(a[135] & b[85])^(a[134] & b[86])^(a[133] & b[87])^(a[132] & b[88])^(a[131] & b[89])^(a[130] & b[90])^(a[129] & b[91])^(a[128] & b[92])^(a[127] & b[93])^(a[126] & b[94])^(a[125] & b[95])^(a[124] & b[96])^(a[123] & b[97])^(a[122] & b[98])^(a[121] & b[99])^(a[120] & b[100])^(a[119] & b[101])^(a[118] & b[102])^(a[117] & b[103])^(a[116] & b[104])^(a[115] & b[105])^(a[114] & b[106])^(a[113] & b[107])^(a[112] & b[108])^(a[111] & b[109])^(a[110] & b[110])^(a[109] & b[111])^(a[108] & b[112])^(a[107] & b[113])^(a[106] & b[114])^(a[105] & b[115])^(a[104] & b[116])^(a[103] & b[117])^(a[102] & b[118])^(a[101] & b[119])^(a[100] & b[120])^(a[99] & b[121])^(a[98] & b[122])^(a[97] & b[123])^(a[96] & b[124])^(a[95] & b[125])^(a[94] & b[126])^(a[93] & b[127])^(a[92] & b[128])^(a[91] & b[129])^(a[90] & b[130])^(a[89] & b[131])^(a[88] & b[132])^(a[87] & b[133])^(a[86] & b[134])^(a[85] & b[135])^(a[84] & b[136])^(a[83] & b[137])^(a[82] & b[138])^(a[81] & b[139])^(a[80] & b[140])^(a[79] & b[141])^(a[78] & b[142])^(a[77] & b[143])^(a[76] & b[144])^(a[75] & b[145])^(a[74] & b[146])^(a[73] & b[147])^(a[72] & b[148])^(a[71] & b[149])^(a[70] & b[150])^(a[69] & b[151])^(a[68] & b[152])^(a[67] & b[153])^(a[66] & b[154])^(a[65] & b[155])^(a[64] & b[156])^(a[63] & b[157])^(a[62] & b[158])^(a[61] & b[159])^(a[60] & b[160])^(a[59] & b[161])^(a[58] & b[162]);
assign y[221] = (a[162] & b[59])^(a[161] & b[60])^(a[160] & b[61])^(a[159] & b[62])^(a[158] & b[63])^(a[157] & b[64])^(a[156] & b[65])^(a[155] & b[66])^(a[154] & b[67])^(a[153] & b[68])^(a[152] & b[69])^(a[151] & b[70])^(a[150] & b[71])^(a[149] & b[72])^(a[148] & b[73])^(a[147] & b[74])^(a[146] & b[75])^(a[145] & b[76])^(a[144] & b[77])^(a[143] & b[78])^(a[142] & b[79])^(a[141] & b[80])^(a[140] & b[81])^(a[139] & b[82])^(a[138] & b[83])^(a[137] & b[84])^(a[136] & b[85])^(a[135] & b[86])^(a[134] & b[87])^(a[133] & b[88])^(a[132] & b[89])^(a[131] & b[90])^(a[130] & b[91])^(a[129] & b[92])^(a[128] & b[93])^(a[127] & b[94])^(a[126] & b[95])^(a[125] & b[96])^(a[124] & b[97])^(a[123] & b[98])^(a[122] & b[99])^(a[121] & b[100])^(a[120] & b[101])^(a[119] & b[102])^(a[118] & b[103])^(a[117] & b[104])^(a[116] & b[105])^(a[115] & b[106])^(a[114] & b[107])^(a[113] & b[108])^(a[112] & b[109])^(a[111] & b[110])^(a[110] & b[111])^(a[109] & b[112])^(a[108] & b[113])^(a[107] & b[114])^(a[106] & b[115])^(a[105] & b[116])^(a[104] & b[117])^(a[103] & b[118])^(a[102] & b[119])^(a[101] & b[120])^(a[100] & b[121])^(a[99] & b[122])^(a[98] & b[123])^(a[97] & b[124])^(a[96] & b[125])^(a[95] & b[126])^(a[94] & b[127])^(a[93] & b[128])^(a[92] & b[129])^(a[91] & b[130])^(a[90] & b[131])^(a[89] & b[132])^(a[88] & b[133])^(a[87] & b[134])^(a[86] & b[135])^(a[85] & b[136])^(a[84] & b[137])^(a[83] & b[138])^(a[82] & b[139])^(a[81] & b[140])^(a[80] & b[141])^(a[79] & b[142])^(a[78] & b[143])^(a[77] & b[144])^(a[76] & b[145])^(a[75] & b[146])^(a[74] & b[147])^(a[73] & b[148])^(a[72] & b[149])^(a[71] & b[150])^(a[70] & b[151])^(a[69] & b[152])^(a[68] & b[153])^(a[67] & b[154])^(a[66] & b[155])^(a[65] & b[156])^(a[64] & b[157])^(a[63] & b[158])^(a[62] & b[159])^(a[61] & b[160])^(a[60] & b[161])^(a[59] & b[162]);
assign y[222] = (a[162] & b[60])^(a[161] & b[61])^(a[160] & b[62])^(a[159] & b[63])^(a[158] & b[64])^(a[157] & b[65])^(a[156] & b[66])^(a[155] & b[67])^(a[154] & b[68])^(a[153] & b[69])^(a[152] & b[70])^(a[151] & b[71])^(a[150] & b[72])^(a[149] & b[73])^(a[148] & b[74])^(a[147] & b[75])^(a[146] & b[76])^(a[145] & b[77])^(a[144] & b[78])^(a[143] & b[79])^(a[142] & b[80])^(a[141] & b[81])^(a[140] & b[82])^(a[139] & b[83])^(a[138] & b[84])^(a[137] & b[85])^(a[136] & b[86])^(a[135] & b[87])^(a[134] & b[88])^(a[133] & b[89])^(a[132] & b[90])^(a[131] & b[91])^(a[130] & b[92])^(a[129] & b[93])^(a[128] & b[94])^(a[127] & b[95])^(a[126] & b[96])^(a[125] & b[97])^(a[124] & b[98])^(a[123] & b[99])^(a[122] & b[100])^(a[121] & b[101])^(a[120] & b[102])^(a[119] & b[103])^(a[118] & b[104])^(a[117] & b[105])^(a[116] & b[106])^(a[115] & b[107])^(a[114] & b[108])^(a[113] & b[109])^(a[112] & b[110])^(a[111] & b[111])^(a[110] & b[112])^(a[109] & b[113])^(a[108] & b[114])^(a[107] & b[115])^(a[106] & b[116])^(a[105] & b[117])^(a[104] & b[118])^(a[103] & b[119])^(a[102] & b[120])^(a[101] & b[121])^(a[100] & b[122])^(a[99] & b[123])^(a[98] & b[124])^(a[97] & b[125])^(a[96] & b[126])^(a[95] & b[127])^(a[94] & b[128])^(a[93] & b[129])^(a[92] & b[130])^(a[91] & b[131])^(a[90] & b[132])^(a[89] & b[133])^(a[88] & b[134])^(a[87] & b[135])^(a[86] & b[136])^(a[85] & b[137])^(a[84] & b[138])^(a[83] & b[139])^(a[82] & b[140])^(a[81] & b[141])^(a[80] & b[142])^(a[79] & b[143])^(a[78] & b[144])^(a[77] & b[145])^(a[76] & b[146])^(a[75] & b[147])^(a[74] & b[148])^(a[73] & b[149])^(a[72] & b[150])^(a[71] & b[151])^(a[70] & b[152])^(a[69] & b[153])^(a[68] & b[154])^(a[67] & b[155])^(a[66] & b[156])^(a[65] & b[157])^(a[64] & b[158])^(a[63] & b[159])^(a[62] & b[160])^(a[61] & b[161])^(a[60] & b[162]);
assign y[223] = (a[162] & b[61])^(a[161] & b[62])^(a[160] & b[63])^(a[159] & b[64])^(a[158] & b[65])^(a[157] & b[66])^(a[156] & b[67])^(a[155] & b[68])^(a[154] & b[69])^(a[153] & b[70])^(a[152] & b[71])^(a[151] & b[72])^(a[150] & b[73])^(a[149] & b[74])^(a[148] & b[75])^(a[147] & b[76])^(a[146] & b[77])^(a[145] & b[78])^(a[144] & b[79])^(a[143] & b[80])^(a[142] & b[81])^(a[141] & b[82])^(a[140] & b[83])^(a[139] & b[84])^(a[138] & b[85])^(a[137] & b[86])^(a[136] & b[87])^(a[135] & b[88])^(a[134] & b[89])^(a[133] & b[90])^(a[132] & b[91])^(a[131] & b[92])^(a[130] & b[93])^(a[129] & b[94])^(a[128] & b[95])^(a[127] & b[96])^(a[126] & b[97])^(a[125] & b[98])^(a[124] & b[99])^(a[123] & b[100])^(a[122] & b[101])^(a[121] & b[102])^(a[120] & b[103])^(a[119] & b[104])^(a[118] & b[105])^(a[117] & b[106])^(a[116] & b[107])^(a[115] & b[108])^(a[114] & b[109])^(a[113] & b[110])^(a[112] & b[111])^(a[111] & b[112])^(a[110] & b[113])^(a[109] & b[114])^(a[108] & b[115])^(a[107] & b[116])^(a[106] & b[117])^(a[105] & b[118])^(a[104] & b[119])^(a[103] & b[120])^(a[102] & b[121])^(a[101] & b[122])^(a[100] & b[123])^(a[99] & b[124])^(a[98] & b[125])^(a[97] & b[126])^(a[96] & b[127])^(a[95] & b[128])^(a[94] & b[129])^(a[93] & b[130])^(a[92] & b[131])^(a[91] & b[132])^(a[90] & b[133])^(a[89] & b[134])^(a[88] & b[135])^(a[87] & b[136])^(a[86] & b[137])^(a[85] & b[138])^(a[84] & b[139])^(a[83] & b[140])^(a[82] & b[141])^(a[81] & b[142])^(a[80] & b[143])^(a[79] & b[144])^(a[78] & b[145])^(a[77] & b[146])^(a[76] & b[147])^(a[75] & b[148])^(a[74] & b[149])^(a[73] & b[150])^(a[72] & b[151])^(a[71] & b[152])^(a[70] & b[153])^(a[69] & b[154])^(a[68] & b[155])^(a[67] & b[156])^(a[66] & b[157])^(a[65] & b[158])^(a[64] & b[159])^(a[63] & b[160])^(a[62] & b[161])^(a[61] & b[162]);
assign y[224] = (a[162] & b[62])^(a[161] & b[63])^(a[160] & b[64])^(a[159] & b[65])^(a[158] & b[66])^(a[157] & b[67])^(a[156] & b[68])^(a[155] & b[69])^(a[154] & b[70])^(a[153] & b[71])^(a[152] & b[72])^(a[151] & b[73])^(a[150] & b[74])^(a[149] & b[75])^(a[148] & b[76])^(a[147] & b[77])^(a[146] & b[78])^(a[145] & b[79])^(a[144] & b[80])^(a[143] & b[81])^(a[142] & b[82])^(a[141] & b[83])^(a[140] & b[84])^(a[139] & b[85])^(a[138] & b[86])^(a[137] & b[87])^(a[136] & b[88])^(a[135] & b[89])^(a[134] & b[90])^(a[133] & b[91])^(a[132] & b[92])^(a[131] & b[93])^(a[130] & b[94])^(a[129] & b[95])^(a[128] & b[96])^(a[127] & b[97])^(a[126] & b[98])^(a[125] & b[99])^(a[124] & b[100])^(a[123] & b[101])^(a[122] & b[102])^(a[121] & b[103])^(a[120] & b[104])^(a[119] & b[105])^(a[118] & b[106])^(a[117] & b[107])^(a[116] & b[108])^(a[115] & b[109])^(a[114] & b[110])^(a[113] & b[111])^(a[112] & b[112])^(a[111] & b[113])^(a[110] & b[114])^(a[109] & b[115])^(a[108] & b[116])^(a[107] & b[117])^(a[106] & b[118])^(a[105] & b[119])^(a[104] & b[120])^(a[103] & b[121])^(a[102] & b[122])^(a[101] & b[123])^(a[100] & b[124])^(a[99] & b[125])^(a[98] & b[126])^(a[97] & b[127])^(a[96] & b[128])^(a[95] & b[129])^(a[94] & b[130])^(a[93] & b[131])^(a[92] & b[132])^(a[91] & b[133])^(a[90] & b[134])^(a[89] & b[135])^(a[88] & b[136])^(a[87] & b[137])^(a[86] & b[138])^(a[85] & b[139])^(a[84] & b[140])^(a[83] & b[141])^(a[82] & b[142])^(a[81] & b[143])^(a[80] & b[144])^(a[79] & b[145])^(a[78] & b[146])^(a[77] & b[147])^(a[76] & b[148])^(a[75] & b[149])^(a[74] & b[150])^(a[73] & b[151])^(a[72] & b[152])^(a[71] & b[153])^(a[70] & b[154])^(a[69] & b[155])^(a[68] & b[156])^(a[67] & b[157])^(a[66] & b[158])^(a[65] & b[159])^(a[64] & b[160])^(a[63] & b[161])^(a[62] & b[162]);
assign y[225] = (a[162] & b[63])^(a[161] & b[64])^(a[160] & b[65])^(a[159] & b[66])^(a[158] & b[67])^(a[157] & b[68])^(a[156] & b[69])^(a[155] & b[70])^(a[154] & b[71])^(a[153] & b[72])^(a[152] & b[73])^(a[151] & b[74])^(a[150] & b[75])^(a[149] & b[76])^(a[148] & b[77])^(a[147] & b[78])^(a[146] & b[79])^(a[145] & b[80])^(a[144] & b[81])^(a[143] & b[82])^(a[142] & b[83])^(a[141] & b[84])^(a[140] & b[85])^(a[139] & b[86])^(a[138] & b[87])^(a[137] & b[88])^(a[136] & b[89])^(a[135] & b[90])^(a[134] & b[91])^(a[133] & b[92])^(a[132] & b[93])^(a[131] & b[94])^(a[130] & b[95])^(a[129] & b[96])^(a[128] & b[97])^(a[127] & b[98])^(a[126] & b[99])^(a[125] & b[100])^(a[124] & b[101])^(a[123] & b[102])^(a[122] & b[103])^(a[121] & b[104])^(a[120] & b[105])^(a[119] & b[106])^(a[118] & b[107])^(a[117] & b[108])^(a[116] & b[109])^(a[115] & b[110])^(a[114] & b[111])^(a[113] & b[112])^(a[112] & b[113])^(a[111] & b[114])^(a[110] & b[115])^(a[109] & b[116])^(a[108] & b[117])^(a[107] & b[118])^(a[106] & b[119])^(a[105] & b[120])^(a[104] & b[121])^(a[103] & b[122])^(a[102] & b[123])^(a[101] & b[124])^(a[100] & b[125])^(a[99] & b[126])^(a[98] & b[127])^(a[97] & b[128])^(a[96] & b[129])^(a[95] & b[130])^(a[94] & b[131])^(a[93] & b[132])^(a[92] & b[133])^(a[91] & b[134])^(a[90] & b[135])^(a[89] & b[136])^(a[88] & b[137])^(a[87] & b[138])^(a[86] & b[139])^(a[85] & b[140])^(a[84] & b[141])^(a[83] & b[142])^(a[82] & b[143])^(a[81] & b[144])^(a[80] & b[145])^(a[79] & b[146])^(a[78] & b[147])^(a[77] & b[148])^(a[76] & b[149])^(a[75] & b[150])^(a[74] & b[151])^(a[73] & b[152])^(a[72] & b[153])^(a[71] & b[154])^(a[70] & b[155])^(a[69] & b[156])^(a[68] & b[157])^(a[67] & b[158])^(a[66] & b[159])^(a[65] & b[160])^(a[64] & b[161])^(a[63] & b[162]);
assign y[226] = (a[162] & b[64])^(a[161] & b[65])^(a[160] & b[66])^(a[159] & b[67])^(a[158] & b[68])^(a[157] & b[69])^(a[156] & b[70])^(a[155] & b[71])^(a[154] & b[72])^(a[153] & b[73])^(a[152] & b[74])^(a[151] & b[75])^(a[150] & b[76])^(a[149] & b[77])^(a[148] & b[78])^(a[147] & b[79])^(a[146] & b[80])^(a[145] & b[81])^(a[144] & b[82])^(a[143] & b[83])^(a[142] & b[84])^(a[141] & b[85])^(a[140] & b[86])^(a[139] & b[87])^(a[138] & b[88])^(a[137] & b[89])^(a[136] & b[90])^(a[135] & b[91])^(a[134] & b[92])^(a[133] & b[93])^(a[132] & b[94])^(a[131] & b[95])^(a[130] & b[96])^(a[129] & b[97])^(a[128] & b[98])^(a[127] & b[99])^(a[126] & b[100])^(a[125] & b[101])^(a[124] & b[102])^(a[123] & b[103])^(a[122] & b[104])^(a[121] & b[105])^(a[120] & b[106])^(a[119] & b[107])^(a[118] & b[108])^(a[117] & b[109])^(a[116] & b[110])^(a[115] & b[111])^(a[114] & b[112])^(a[113] & b[113])^(a[112] & b[114])^(a[111] & b[115])^(a[110] & b[116])^(a[109] & b[117])^(a[108] & b[118])^(a[107] & b[119])^(a[106] & b[120])^(a[105] & b[121])^(a[104] & b[122])^(a[103] & b[123])^(a[102] & b[124])^(a[101] & b[125])^(a[100] & b[126])^(a[99] & b[127])^(a[98] & b[128])^(a[97] & b[129])^(a[96] & b[130])^(a[95] & b[131])^(a[94] & b[132])^(a[93] & b[133])^(a[92] & b[134])^(a[91] & b[135])^(a[90] & b[136])^(a[89] & b[137])^(a[88] & b[138])^(a[87] & b[139])^(a[86] & b[140])^(a[85] & b[141])^(a[84] & b[142])^(a[83] & b[143])^(a[82] & b[144])^(a[81] & b[145])^(a[80] & b[146])^(a[79] & b[147])^(a[78] & b[148])^(a[77] & b[149])^(a[76] & b[150])^(a[75] & b[151])^(a[74] & b[152])^(a[73] & b[153])^(a[72] & b[154])^(a[71] & b[155])^(a[70] & b[156])^(a[69] & b[157])^(a[68] & b[158])^(a[67] & b[159])^(a[66] & b[160])^(a[65] & b[161])^(a[64] & b[162]);
assign y[227] = (a[162] & b[65])^(a[161] & b[66])^(a[160] & b[67])^(a[159] & b[68])^(a[158] & b[69])^(a[157] & b[70])^(a[156] & b[71])^(a[155] & b[72])^(a[154] & b[73])^(a[153] & b[74])^(a[152] & b[75])^(a[151] & b[76])^(a[150] & b[77])^(a[149] & b[78])^(a[148] & b[79])^(a[147] & b[80])^(a[146] & b[81])^(a[145] & b[82])^(a[144] & b[83])^(a[143] & b[84])^(a[142] & b[85])^(a[141] & b[86])^(a[140] & b[87])^(a[139] & b[88])^(a[138] & b[89])^(a[137] & b[90])^(a[136] & b[91])^(a[135] & b[92])^(a[134] & b[93])^(a[133] & b[94])^(a[132] & b[95])^(a[131] & b[96])^(a[130] & b[97])^(a[129] & b[98])^(a[128] & b[99])^(a[127] & b[100])^(a[126] & b[101])^(a[125] & b[102])^(a[124] & b[103])^(a[123] & b[104])^(a[122] & b[105])^(a[121] & b[106])^(a[120] & b[107])^(a[119] & b[108])^(a[118] & b[109])^(a[117] & b[110])^(a[116] & b[111])^(a[115] & b[112])^(a[114] & b[113])^(a[113] & b[114])^(a[112] & b[115])^(a[111] & b[116])^(a[110] & b[117])^(a[109] & b[118])^(a[108] & b[119])^(a[107] & b[120])^(a[106] & b[121])^(a[105] & b[122])^(a[104] & b[123])^(a[103] & b[124])^(a[102] & b[125])^(a[101] & b[126])^(a[100] & b[127])^(a[99] & b[128])^(a[98] & b[129])^(a[97] & b[130])^(a[96] & b[131])^(a[95] & b[132])^(a[94] & b[133])^(a[93] & b[134])^(a[92] & b[135])^(a[91] & b[136])^(a[90] & b[137])^(a[89] & b[138])^(a[88] & b[139])^(a[87] & b[140])^(a[86] & b[141])^(a[85] & b[142])^(a[84] & b[143])^(a[83] & b[144])^(a[82] & b[145])^(a[81] & b[146])^(a[80] & b[147])^(a[79] & b[148])^(a[78] & b[149])^(a[77] & b[150])^(a[76] & b[151])^(a[75] & b[152])^(a[74] & b[153])^(a[73] & b[154])^(a[72] & b[155])^(a[71] & b[156])^(a[70] & b[157])^(a[69] & b[158])^(a[68] & b[159])^(a[67] & b[160])^(a[66] & b[161])^(a[65] & b[162]);
assign y[228] = (a[162] & b[66])^(a[161] & b[67])^(a[160] & b[68])^(a[159] & b[69])^(a[158] & b[70])^(a[157] & b[71])^(a[156] & b[72])^(a[155] & b[73])^(a[154] & b[74])^(a[153] & b[75])^(a[152] & b[76])^(a[151] & b[77])^(a[150] & b[78])^(a[149] & b[79])^(a[148] & b[80])^(a[147] & b[81])^(a[146] & b[82])^(a[145] & b[83])^(a[144] & b[84])^(a[143] & b[85])^(a[142] & b[86])^(a[141] & b[87])^(a[140] & b[88])^(a[139] & b[89])^(a[138] & b[90])^(a[137] & b[91])^(a[136] & b[92])^(a[135] & b[93])^(a[134] & b[94])^(a[133] & b[95])^(a[132] & b[96])^(a[131] & b[97])^(a[130] & b[98])^(a[129] & b[99])^(a[128] & b[100])^(a[127] & b[101])^(a[126] & b[102])^(a[125] & b[103])^(a[124] & b[104])^(a[123] & b[105])^(a[122] & b[106])^(a[121] & b[107])^(a[120] & b[108])^(a[119] & b[109])^(a[118] & b[110])^(a[117] & b[111])^(a[116] & b[112])^(a[115] & b[113])^(a[114] & b[114])^(a[113] & b[115])^(a[112] & b[116])^(a[111] & b[117])^(a[110] & b[118])^(a[109] & b[119])^(a[108] & b[120])^(a[107] & b[121])^(a[106] & b[122])^(a[105] & b[123])^(a[104] & b[124])^(a[103] & b[125])^(a[102] & b[126])^(a[101] & b[127])^(a[100] & b[128])^(a[99] & b[129])^(a[98] & b[130])^(a[97] & b[131])^(a[96] & b[132])^(a[95] & b[133])^(a[94] & b[134])^(a[93] & b[135])^(a[92] & b[136])^(a[91] & b[137])^(a[90] & b[138])^(a[89] & b[139])^(a[88] & b[140])^(a[87] & b[141])^(a[86] & b[142])^(a[85] & b[143])^(a[84] & b[144])^(a[83] & b[145])^(a[82] & b[146])^(a[81] & b[147])^(a[80] & b[148])^(a[79] & b[149])^(a[78] & b[150])^(a[77] & b[151])^(a[76] & b[152])^(a[75] & b[153])^(a[74] & b[154])^(a[73] & b[155])^(a[72] & b[156])^(a[71] & b[157])^(a[70] & b[158])^(a[69] & b[159])^(a[68] & b[160])^(a[67] & b[161])^(a[66] & b[162]);
assign y[229] = (a[162] & b[67])^(a[161] & b[68])^(a[160] & b[69])^(a[159] & b[70])^(a[158] & b[71])^(a[157] & b[72])^(a[156] & b[73])^(a[155] & b[74])^(a[154] & b[75])^(a[153] & b[76])^(a[152] & b[77])^(a[151] & b[78])^(a[150] & b[79])^(a[149] & b[80])^(a[148] & b[81])^(a[147] & b[82])^(a[146] & b[83])^(a[145] & b[84])^(a[144] & b[85])^(a[143] & b[86])^(a[142] & b[87])^(a[141] & b[88])^(a[140] & b[89])^(a[139] & b[90])^(a[138] & b[91])^(a[137] & b[92])^(a[136] & b[93])^(a[135] & b[94])^(a[134] & b[95])^(a[133] & b[96])^(a[132] & b[97])^(a[131] & b[98])^(a[130] & b[99])^(a[129] & b[100])^(a[128] & b[101])^(a[127] & b[102])^(a[126] & b[103])^(a[125] & b[104])^(a[124] & b[105])^(a[123] & b[106])^(a[122] & b[107])^(a[121] & b[108])^(a[120] & b[109])^(a[119] & b[110])^(a[118] & b[111])^(a[117] & b[112])^(a[116] & b[113])^(a[115] & b[114])^(a[114] & b[115])^(a[113] & b[116])^(a[112] & b[117])^(a[111] & b[118])^(a[110] & b[119])^(a[109] & b[120])^(a[108] & b[121])^(a[107] & b[122])^(a[106] & b[123])^(a[105] & b[124])^(a[104] & b[125])^(a[103] & b[126])^(a[102] & b[127])^(a[101] & b[128])^(a[100] & b[129])^(a[99] & b[130])^(a[98] & b[131])^(a[97] & b[132])^(a[96] & b[133])^(a[95] & b[134])^(a[94] & b[135])^(a[93] & b[136])^(a[92] & b[137])^(a[91] & b[138])^(a[90] & b[139])^(a[89] & b[140])^(a[88] & b[141])^(a[87] & b[142])^(a[86] & b[143])^(a[85] & b[144])^(a[84] & b[145])^(a[83] & b[146])^(a[82] & b[147])^(a[81] & b[148])^(a[80] & b[149])^(a[79] & b[150])^(a[78] & b[151])^(a[77] & b[152])^(a[76] & b[153])^(a[75] & b[154])^(a[74] & b[155])^(a[73] & b[156])^(a[72] & b[157])^(a[71] & b[158])^(a[70] & b[159])^(a[69] & b[160])^(a[68] & b[161])^(a[67] & b[162]);
assign y[230] = (a[162] & b[68])^(a[161] & b[69])^(a[160] & b[70])^(a[159] & b[71])^(a[158] & b[72])^(a[157] & b[73])^(a[156] & b[74])^(a[155] & b[75])^(a[154] & b[76])^(a[153] & b[77])^(a[152] & b[78])^(a[151] & b[79])^(a[150] & b[80])^(a[149] & b[81])^(a[148] & b[82])^(a[147] & b[83])^(a[146] & b[84])^(a[145] & b[85])^(a[144] & b[86])^(a[143] & b[87])^(a[142] & b[88])^(a[141] & b[89])^(a[140] & b[90])^(a[139] & b[91])^(a[138] & b[92])^(a[137] & b[93])^(a[136] & b[94])^(a[135] & b[95])^(a[134] & b[96])^(a[133] & b[97])^(a[132] & b[98])^(a[131] & b[99])^(a[130] & b[100])^(a[129] & b[101])^(a[128] & b[102])^(a[127] & b[103])^(a[126] & b[104])^(a[125] & b[105])^(a[124] & b[106])^(a[123] & b[107])^(a[122] & b[108])^(a[121] & b[109])^(a[120] & b[110])^(a[119] & b[111])^(a[118] & b[112])^(a[117] & b[113])^(a[116] & b[114])^(a[115] & b[115])^(a[114] & b[116])^(a[113] & b[117])^(a[112] & b[118])^(a[111] & b[119])^(a[110] & b[120])^(a[109] & b[121])^(a[108] & b[122])^(a[107] & b[123])^(a[106] & b[124])^(a[105] & b[125])^(a[104] & b[126])^(a[103] & b[127])^(a[102] & b[128])^(a[101] & b[129])^(a[100] & b[130])^(a[99] & b[131])^(a[98] & b[132])^(a[97] & b[133])^(a[96] & b[134])^(a[95] & b[135])^(a[94] & b[136])^(a[93] & b[137])^(a[92] & b[138])^(a[91] & b[139])^(a[90] & b[140])^(a[89] & b[141])^(a[88] & b[142])^(a[87] & b[143])^(a[86] & b[144])^(a[85] & b[145])^(a[84] & b[146])^(a[83] & b[147])^(a[82] & b[148])^(a[81] & b[149])^(a[80] & b[150])^(a[79] & b[151])^(a[78] & b[152])^(a[77] & b[153])^(a[76] & b[154])^(a[75] & b[155])^(a[74] & b[156])^(a[73] & b[157])^(a[72] & b[158])^(a[71] & b[159])^(a[70] & b[160])^(a[69] & b[161])^(a[68] & b[162]);
assign y[231] = (a[162] & b[69])^(a[161] & b[70])^(a[160] & b[71])^(a[159] & b[72])^(a[158] & b[73])^(a[157] & b[74])^(a[156] & b[75])^(a[155] & b[76])^(a[154] & b[77])^(a[153] & b[78])^(a[152] & b[79])^(a[151] & b[80])^(a[150] & b[81])^(a[149] & b[82])^(a[148] & b[83])^(a[147] & b[84])^(a[146] & b[85])^(a[145] & b[86])^(a[144] & b[87])^(a[143] & b[88])^(a[142] & b[89])^(a[141] & b[90])^(a[140] & b[91])^(a[139] & b[92])^(a[138] & b[93])^(a[137] & b[94])^(a[136] & b[95])^(a[135] & b[96])^(a[134] & b[97])^(a[133] & b[98])^(a[132] & b[99])^(a[131] & b[100])^(a[130] & b[101])^(a[129] & b[102])^(a[128] & b[103])^(a[127] & b[104])^(a[126] & b[105])^(a[125] & b[106])^(a[124] & b[107])^(a[123] & b[108])^(a[122] & b[109])^(a[121] & b[110])^(a[120] & b[111])^(a[119] & b[112])^(a[118] & b[113])^(a[117] & b[114])^(a[116] & b[115])^(a[115] & b[116])^(a[114] & b[117])^(a[113] & b[118])^(a[112] & b[119])^(a[111] & b[120])^(a[110] & b[121])^(a[109] & b[122])^(a[108] & b[123])^(a[107] & b[124])^(a[106] & b[125])^(a[105] & b[126])^(a[104] & b[127])^(a[103] & b[128])^(a[102] & b[129])^(a[101] & b[130])^(a[100] & b[131])^(a[99] & b[132])^(a[98] & b[133])^(a[97] & b[134])^(a[96] & b[135])^(a[95] & b[136])^(a[94] & b[137])^(a[93] & b[138])^(a[92] & b[139])^(a[91] & b[140])^(a[90] & b[141])^(a[89] & b[142])^(a[88] & b[143])^(a[87] & b[144])^(a[86] & b[145])^(a[85] & b[146])^(a[84] & b[147])^(a[83] & b[148])^(a[82] & b[149])^(a[81] & b[150])^(a[80] & b[151])^(a[79] & b[152])^(a[78] & b[153])^(a[77] & b[154])^(a[76] & b[155])^(a[75] & b[156])^(a[74] & b[157])^(a[73] & b[158])^(a[72] & b[159])^(a[71] & b[160])^(a[70] & b[161])^(a[69] & b[162]);
assign y[232] = (a[162] & b[70])^(a[161] & b[71])^(a[160] & b[72])^(a[159] & b[73])^(a[158] & b[74])^(a[157] & b[75])^(a[156] & b[76])^(a[155] & b[77])^(a[154] & b[78])^(a[153] & b[79])^(a[152] & b[80])^(a[151] & b[81])^(a[150] & b[82])^(a[149] & b[83])^(a[148] & b[84])^(a[147] & b[85])^(a[146] & b[86])^(a[145] & b[87])^(a[144] & b[88])^(a[143] & b[89])^(a[142] & b[90])^(a[141] & b[91])^(a[140] & b[92])^(a[139] & b[93])^(a[138] & b[94])^(a[137] & b[95])^(a[136] & b[96])^(a[135] & b[97])^(a[134] & b[98])^(a[133] & b[99])^(a[132] & b[100])^(a[131] & b[101])^(a[130] & b[102])^(a[129] & b[103])^(a[128] & b[104])^(a[127] & b[105])^(a[126] & b[106])^(a[125] & b[107])^(a[124] & b[108])^(a[123] & b[109])^(a[122] & b[110])^(a[121] & b[111])^(a[120] & b[112])^(a[119] & b[113])^(a[118] & b[114])^(a[117] & b[115])^(a[116] & b[116])^(a[115] & b[117])^(a[114] & b[118])^(a[113] & b[119])^(a[112] & b[120])^(a[111] & b[121])^(a[110] & b[122])^(a[109] & b[123])^(a[108] & b[124])^(a[107] & b[125])^(a[106] & b[126])^(a[105] & b[127])^(a[104] & b[128])^(a[103] & b[129])^(a[102] & b[130])^(a[101] & b[131])^(a[100] & b[132])^(a[99] & b[133])^(a[98] & b[134])^(a[97] & b[135])^(a[96] & b[136])^(a[95] & b[137])^(a[94] & b[138])^(a[93] & b[139])^(a[92] & b[140])^(a[91] & b[141])^(a[90] & b[142])^(a[89] & b[143])^(a[88] & b[144])^(a[87] & b[145])^(a[86] & b[146])^(a[85] & b[147])^(a[84] & b[148])^(a[83] & b[149])^(a[82] & b[150])^(a[81] & b[151])^(a[80] & b[152])^(a[79] & b[153])^(a[78] & b[154])^(a[77] & b[155])^(a[76] & b[156])^(a[75] & b[157])^(a[74] & b[158])^(a[73] & b[159])^(a[72] & b[160])^(a[71] & b[161])^(a[70] & b[162]);
assign y[233] = (a[162] & b[71])^(a[161] & b[72])^(a[160] & b[73])^(a[159] & b[74])^(a[158] & b[75])^(a[157] & b[76])^(a[156] & b[77])^(a[155] & b[78])^(a[154] & b[79])^(a[153] & b[80])^(a[152] & b[81])^(a[151] & b[82])^(a[150] & b[83])^(a[149] & b[84])^(a[148] & b[85])^(a[147] & b[86])^(a[146] & b[87])^(a[145] & b[88])^(a[144] & b[89])^(a[143] & b[90])^(a[142] & b[91])^(a[141] & b[92])^(a[140] & b[93])^(a[139] & b[94])^(a[138] & b[95])^(a[137] & b[96])^(a[136] & b[97])^(a[135] & b[98])^(a[134] & b[99])^(a[133] & b[100])^(a[132] & b[101])^(a[131] & b[102])^(a[130] & b[103])^(a[129] & b[104])^(a[128] & b[105])^(a[127] & b[106])^(a[126] & b[107])^(a[125] & b[108])^(a[124] & b[109])^(a[123] & b[110])^(a[122] & b[111])^(a[121] & b[112])^(a[120] & b[113])^(a[119] & b[114])^(a[118] & b[115])^(a[117] & b[116])^(a[116] & b[117])^(a[115] & b[118])^(a[114] & b[119])^(a[113] & b[120])^(a[112] & b[121])^(a[111] & b[122])^(a[110] & b[123])^(a[109] & b[124])^(a[108] & b[125])^(a[107] & b[126])^(a[106] & b[127])^(a[105] & b[128])^(a[104] & b[129])^(a[103] & b[130])^(a[102] & b[131])^(a[101] & b[132])^(a[100] & b[133])^(a[99] & b[134])^(a[98] & b[135])^(a[97] & b[136])^(a[96] & b[137])^(a[95] & b[138])^(a[94] & b[139])^(a[93] & b[140])^(a[92] & b[141])^(a[91] & b[142])^(a[90] & b[143])^(a[89] & b[144])^(a[88] & b[145])^(a[87] & b[146])^(a[86] & b[147])^(a[85] & b[148])^(a[84] & b[149])^(a[83] & b[150])^(a[82] & b[151])^(a[81] & b[152])^(a[80] & b[153])^(a[79] & b[154])^(a[78] & b[155])^(a[77] & b[156])^(a[76] & b[157])^(a[75] & b[158])^(a[74] & b[159])^(a[73] & b[160])^(a[72] & b[161])^(a[71] & b[162]);
assign y[234] = (a[162] & b[72])^(a[161] & b[73])^(a[160] & b[74])^(a[159] & b[75])^(a[158] & b[76])^(a[157] & b[77])^(a[156] & b[78])^(a[155] & b[79])^(a[154] & b[80])^(a[153] & b[81])^(a[152] & b[82])^(a[151] & b[83])^(a[150] & b[84])^(a[149] & b[85])^(a[148] & b[86])^(a[147] & b[87])^(a[146] & b[88])^(a[145] & b[89])^(a[144] & b[90])^(a[143] & b[91])^(a[142] & b[92])^(a[141] & b[93])^(a[140] & b[94])^(a[139] & b[95])^(a[138] & b[96])^(a[137] & b[97])^(a[136] & b[98])^(a[135] & b[99])^(a[134] & b[100])^(a[133] & b[101])^(a[132] & b[102])^(a[131] & b[103])^(a[130] & b[104])^(a[129] & b[105])^(a[128] & b[106])^(a[127] & b[107])^(a[126] & b[108])^(a[125] & b[109])^(a[124] & b[110])^(a[123] & b[111])^(a[122] & b[112])^(a[121] & b[113])^(a[120] & b[114])^(a[119] & b[115])^(a[118] & b[116])^(a[117] & b[117])^(a[116] & b[118])^(a[115] & b[119])^(a[114] & b[120])^(a[113] & b[121])^(a[112] & b[122])^(a[111] & b[123])^(a[110] & b[124])^(a[109] & b[125])^(a[108] & b[126])^(a[107] & b[127])^(a[106] & b[128])^(a[105] & b[129])^(a[104] & b[130])^(a[103] & b[131])^(a[102] & b[132])^(a[101] & b[133])^(a[100] & b[134])^(a[99] & b[135])^(a[98] & b[136])^(a[97] & b[137])^(a[96] & b[138])^(a[95] & b[139])^(a[94] & b[140])^(a[93] & b[141])^(a[92] & b[142])^(a[91] & b[143])^(a[90] & b[144])^(a[89] & b[145])^(a[88] & b[146])^(a[87] & b[147])^(a[86] & b[148])^(a[85] & b[149])^(a[84] & b[150])^(a[83] & b[151])^(a[82] & b[152])^(a[81] & b[153])^(a[80] & b[154])^(a[79] & b[155])^(a[78] & b[156])^(a[77] & b[157])^(a[76] & b[158])^(a[75] & b[159])^(a[74] & b[160])^(a[73] & b[161])^(a[72] & b[162]);
assign y[235] = (a[162] & b[73])^(a[161] & b[74])^(a[160] & b[75])^(a[159] & b[76])^(a[158] & b[77])^(a[157] & b[78])^(a[156] & b[79])^(a[155] & b[80])^(a[154] & b[81])^(a[153] & b[82])^(a[152] & b[83])^(a[151] & b[84])^(a[150] & b[85])^(a[149] & b[86])^(a[148] & b[87])^(a[147] & b[88])^(a[146] & b[89])^(a[145] & b[90])^(a[144] & b[91])^(a[143] & b[92])^(a[142] & b[93])^(a[141] & b[94])^(a[140] & b[95])^(a[139] & b[96])^(a[138] & b[97])^(a[137] & b[98])^(a[136] & b[99])^(a[135] & b[100])^(a[134] & b[101])^(a[133] & b[102])^(a[132] & b[103])^(a[131] & b[104])^(a[130] & b[105])^(a[129] & b[106])^(a[128] & b[107])^(a[127] & b[108])^(a[126] & b[109])^(a[125] & b[110])^(a[124] & b[111])^(a[123] & b[112])^(a[122] & b[113])^(a[121] & b[114])^(a[120] & b[115])^(a[119] & b[116])^(a[118] & b[117])^(a[117] & b[118])^(a[116] & b[119])^(a[115] & b[120])^(a[114] & b[121])^(a[113] & b[122])^(a[112] & b[123])^(a[111] & b[124])^(a[110] & b[125])^(a[109] & b[126])^(a[108] & b[127])^(a[107] & b[128])^(a[106] & b[129])^(a[105] & b[130])^(a[104] & b[131])^(a[103] & b[132])^(a[102] & b[133])^(a[101] & b[134])^(a[100] & b[135])^(a[99] & b[136])^(a[98] & b[137])^(a[97] & b[138])^(a[96] & b[139])^(a[95] & b[140])^(a[94] & b[141])^(a[93] & b[142])^(a[92] & b[143])^(a[91] & b[144])^(a[90] & b[145])^(a[89] & b[146])^(a[88] & b[147])^(a[87] & b[148])^(a[86] & b[149])^(a[85] & b[150])^(a[84] & b[151])^(a[83] & b[152])^(a[82] & b[153])^(a[81] & b[154])^(a[80] & b[155])^(a[79] & b[156])^(a[78] & b[157])^(a[77] & b[158])^(a[76] & b[159])^(a[75] & b[160])^(a[74] & b[161])^(a[73] & b[162]);
assign y[236] = (a[162] & b[74])^(a[161] & b[75])^(a[160] & b[76])^(a[159] & b[77])^(a[158] & b[78])^(a[157] & b[79])^(a[156] & b[80])^(a[155] & b[81])^(a[154] & b[82])^(a[153] & b[83])^(a[152] & b[84])^(a[151] & b[85])^(a[150] & b[86])^(a[149] & b[87])^(a[148] & b[88])^(a[147] & b[89])^(a[146] & b[90])^(a[145] & b[91])^(a[144] & b[92])^(a[143] & b[93])^(a[142] & b[94])^(a[141] & b[95])^(a[140] & b[96])^(a[139] & b[97])^(a[138] & b[98])^(a[137] & b[99])^(a[136] & b[100])^(a[135] & b[101])^(a[134] & b[102])^(a[133] & b[103])^(a[132] & b[104])^(a[131] & b[105])^(a[130] & b[106])^(a[129] & b[107])^(a[128] & b[108])^(a[127] & b[109])^(a[126] & b[110])^(a[125] & b[111])^(a[124] & b[112])^(a[123] & b[113])^(a[122] & b[114])^(a[121] & b[115])^(a[120] & b[116])^(a[119] & b[117])^(a[118] & b[118])^(a[117] & b[119])^(a[116] & b[120])^(a[115] & b[121])^(a[114] & b[122])^(a[113] & b[123])^(a[112] & b[124])^(a[111] & b[125])^(a[110] & b[126])^(a[109] & b[127])^(a[108] & b[128])^(a[107] & b[129])^(a[106] & b[130])^(a[105] & b[131])^(a[104] & b[132])^(a[103] & b[133])^(a[102] & b[134])^(a[101] & b[135])^(a[100] & b[136])^(a[99] & b[137])^(a[98] & b[138])^(a[97] & b[139])^(a[96] & b[140])^(a[95] & b[141])^(a[94] & b[142])^(a[93] & b[143])^(a[92] & b[144])^(a[91] & b[145])^(a[90] & b[146])^(a[89] & b[147])^(a[88] & b[148])^(a[87] & b[149])^(a[86] & b[150])^(a[85] & b[151])^(a[84] & b[152])^(a[83] & b[153])^(a[82] & b[154])^(a[81] & b[155])^(a[80] & b[156])^(a[79] & b[157])^(a[78] & b[158])^(a[77] & b[159])^(a[76] & b[160])^(a[75] & b[161])^(a[74] & b[162]);
assign y[237] = (a[162] & b[75])^(a[161] & b[76])^(a[160] & b[77])^(a[159] & b[78])^(a[158] & b[79])^(a[157] & b[80])^(a[156] & b[81])^(a[155] & b[82])^(a[154] & b[83])^(a[153] & b[84])^(a[152] & b[85])^(a[151] & b[86])^(a[150] & b[87])^(a[149] & b[88])^(a[148] & b[89])^(a[147] & b[90])^(a[146] & b[91])^(a[145] & b[92])^(a[144] & b[93])^(a[143] & b[94])^(a[142] & b[95])^(a[141] & b[96])^(a[140] & b[97])^(a[139] & b[98])^(a[138] & b[99])^(a[137] & b[100])^(a[136] & b[101])^(a[135] & b[102])^(a[134] & b[103])^(a[133] & b[104])^(a[132] & b[105])^(a[131] & b[106])^(a[130] & b[107])^(a[129] & b[108])^(a[128] & b[109])^(a[127] & b[110])^(a[126] & b[111])^(a[125] & b[112])^(a[124] & b[113])^(a[123] & b[114])^(a[122] & b[115])^(a[121] & b[116])^(a[120] & b[117])^(a[119] & b[118])^(a[118] & b[119])^(a[117] & b[120])^(a[116] & b[121])^(a[115] & b[122])^(a[114] & b[123])^(a[113] & b[124])^(a[112] & b[125])^(a[111] & b[126])^(a[110] & b[127])^(a[109] & b[128])^(a[108] & b[129])^(a[107] & b[130])^(a[106] & b[131])^(a[105] & b[132])^(a[104] & b[133])^(a[103] & b[134])^(a[102] & b[135])^(a[101] & b[136])^(a[100] & b[137])^(a[99] & b[138])^(a[98] & b[139])^(a[97] & b[140])^(a[96] & b[141])^(a[95] & b[142])^(a[94] & b[143])^(a[93] & b[144])^(a[92] & b[145])^(a[91] & b[146])^(a[90] & b[147])^(a[89] & b[148])^(a[88] & b[149])^(a[87] & b[150])^(a[86] & b[151])^(a[85] & b[152])^(a[84] & b[153])^(a[83] & b[154])^(a[82] & b[155])^(a[81] & b[156])^(a[80] & b[157])^(a[79] & b[158])^(a[78] & b[159])^(a[77] & b[160])^(a[76] & b[161])^(a[75] & b[162]);
assign y[238] = (a[162] & b[76])^(a[161] & b[77])^(a[160] & b[78])^(a[159] & b[79])^(a[158] & b[80])^(a[157] & b[81])^(a[156] & b[82])^(a[155] & b[83])^(a[154] & b[84])^(a[153] & b[85])^(a[152] & b[86])^(a[151] & b[87])^(a[150] & b[88])^(a[149] & b[89])^(a[148] & b[90])^(a[147] & b[91])^(a[146] & b[92])^(a[145] & b[93])^(a[144] & b[94])^(a[143] & b[95])^(a[142] & b[96])^(a[141] & b[97])^(a[140] & b[98])^(a[139] & b[99])^(a[138] & b[100])^(a[137] & b[101])^(a[136] & b[102])^(a[135] & b[103])^(a[134] & b[104])^(a[133] & b[105])^(a[132] & b[106])^(a[131] & b[107])^(a[130] & b[108])^(a[129] & b[109])^(a[128] & b[110])^(a[127] & b[111])^(a[126] & b[112])^(a[125] & b[113])^(a[124] & b[114])^(a[123] & b[115])^(a[122] & b[116])^(a[121] & b[117])^(a[120] & b[118])^(a[119] & b[119])^(a[118] & b[120])^(a[117] & b[121])^(a[116] & b[122])^(a[115] & b[123])^(a[114] & b[124])^(a[113] & b[125])^(a[112] & b[126])^(a[111] & b[127])^(a[110] & b[128])^(a[109] & b[129])^(a[108] & b[130])^(a[107] & b[131])^(a[106] & b[132])^(a[105] & b[133])^(a[104] & b[134])^(a[103] & b[135])^(a[102] & b[136])^(a[101] & b[137])^(a[100] & b[138])^(a[99] & b[139])^(a[98] & b[140])^(a[97] & b[141])^(a[96] & b[142])^(a[95] & b[143])^(a[94] & b[144])^(a[93] & b[145])^(a[92] & b[146])^(a[91] & b[147])^(a[90] & b[148])^(a[89] & b[149])^(a[88] & b[150])^(a[87] & b[151])^(a[86] & b[152])^(a[85] & b[153])^(a[84] & b[154])^(a[83] & b[155])^(a[82] & b[156])^(a[81] & b[157])^(a[80] & b[158])^(a[79] & b[159])^(a[78] & b[160])^(a[77] & b[161])^(a[76] & b[162]);
assign y[239] = (a[162] & b[77])^(a[161] & b[78])^(a[160] & b[79])^(a[159] & b[80])^(a[158] & b[81])^(a[157] & b[82])^(a[156] & b[83])^(a[155] & b[84])^(a[154] & b[85])^(a[153] & b[86])^(a[152] & b[87])^(a[151] & b[88])^(a[150] & b[89])^(a[149] & b[90])^(a[148] & b[91])^(a[147] & b[92])^(a[146] & b[93])^(a[145] & b[94])^(a[144] & b[95])^(a[143] & b[96])^(a[142] & b[97])^(a[141] & b[98])^(a[140] & b[99])^(a[139] & b[100])^(a[138] & b[101])^(a[137] & b[102])^(a[136] & b[103])^(a[135] & b[104])^(a[134] & b[105])^(a[133] & b[106])^(a[132] & b[107])^(a[131] & b[108])^(a[130] & b[109])^(a[129] & b[110])^(a[128] & b[111])^(a[127] & b[112])^(a[126] & b[113])^(a[125] & b[114])^(a[124] & b[115])^(a[123] & b[116])^(a[122] & b[117])^(a[121] & b[118])^(a[120] & b[119])^(a[119] & b[120])^(a[118] & b[121])^(a[117] & b[122])^(a[116] & b[123])^(a[115] & b[124])^(a[114] & b[125])^(a[113] & b[126])^(a[112] & b[127])^(a[111] & b[128])^(a[110] & b[129])^(a[109] & b[130])^(a[108] & b[131])^(a[107] & b[132])^(a[106] & b[133])^(a[105] & b[134])^(a[104] & b[135])^(a[103] & b[136])^(a[102] & b[137])^(a[101] & b[138])^(a[100] & b[139])^(a[99] & b[140])^(a[98] & b[141])^(a[97] & b[142])^(a[96] & b[143])^(a[95] & b[144])^(a[94] & b[145])^(a[93] & b[146])^(a[92] & b[147])^(a[91] & b[148])^(a[90] & b[149])^(a[89] & b[150])^(a[88] & b[151])^(a[87] & b[152])^(a[86] & b[153])^(a[85] & b[154])^(a[84] & b[155])^(a[83] & b[156])^(a[82] & b[157])^(a[81] & b[158])^(a[80] & b[159])^(a[79] & b[160])^(a[78] & b[161])^(a[77] & b[162]);
assign y[240] = (a[162] & b[78])^(a[161] & b[79])^(a[160] & b[80])^(a[159] & b[81])^(a[158] & b[82])^(a[157] & b[83])^(a[156] & b[84])^(a[155] & b[85])^(a[154] & b[86])^(a[153] & b[87])^(a[152] & b[88])^(a[151] & b[89])^(a[150] & b[90])^(a[149] & b[91])^(a[148] & b[92])^(a[147] & b[93])^(a[146] & b[94])^(a[145] & b[95])^(a[144] & b[96])^(a[143] & b[97])^(a[142] & b[98])^(a[141] & b[99])^(a[140] & b[100])^(a[139] & b[101])^(a[138] & b[102])^(a[137] & b[103])^(a[136] & b[104])^(a[135] & b[105])^(a[134] & b[106])^(a[133] & b[107])^(a[132] & b[108])^(a[131] & b[109])^(a[130] & b[110])^(a[129] & b[111])^(a[128] & b[112])^(a[127] & b[113])^(a[126] & b[114])^(a[125] & b[115])^(a[124] & b[116])^(a[123] & b[117])^(a[122] & b[118])^(a[121] & b[119])^(a[120] & b[120])^(a[119] & b[121])^(a[118] & b[122])^(a[117] & b[123])^(a[116] & b[124])^(a[115] & b[125])^(a[114] & b[126])^(a[113] & b[127])^(a[112] & b[128])^(a[111] & b[129])^(a[110] & b[130])^(a[109] & b[131])^(a[108] & b[132])^(a[107] & b[133])^(a[106] & b[134])^(a[105] & b[135])^(a[104] & b[136])^(a[103] & b[137])^(a[102] & b[138])^(a[101] & b[139])^(a[100] & b[140])^(a[99] & b[141])^(a[98] & b[142])^(a[97] & b[143])^(a[96] & b[144])^(a[95] & b[145])^(a[94] & b[146])^(a[93] & b[147])^(a[92] & b[148])^(a[91] & b[149])^(a[90] & b[150])^(a[89] & b[151])^(a[88] & b[152])^(a[87] & b[153])^(a[86] & b[154])^(a[85] & b[155])^(a[84] & b[156])^(a[83] & b[157])^(a[82] & b[158])^(a[81] & b[159])^(a[80] & b[160])^(a[79] & b[161])^(a[78] & b[162]);
assign y[241] = (a[162] & b[79])^(a[161] & b[80])^(a[160] & b[81])^(a[159] & b[82])^(a[158] & b[83])^(a[157] & b[84])^(a[156] & b[85])^(a[155] & b[86])^(a[154] & b[87])^(a[153] & b[88])^(a[152] & b[89])^(a[151] & b[90])^(a[150] & b[91])^(a[149] & b[92])^(a[148] & b[93])^(a[147] & b[94])^(a[146] & b[95])^(a[145] & b[96])^(a[144] & b[97])^(a[143] & b[98])^(a[142] & b[99])^(a[141] & b[100])^(a[140] & b[101])^(a[139] & b[102])^(a[138] & b[103])^(a[137] & b[104])^(a[136] & b[105])^(a[135] & b[106])^(a[134] & b[107])^(a[133] & b[108])^(a[132] & b[109])^(a[131] & b[110])^(a[130] & b[111])^(a[129] & b[112])^(a[128] & b[113])^(a[127] & b[114])^(a[126] & b[115])^(a[125] & b[116])^(a[124] & b[117])^(a[123] & b[118])^(a[122] & b[119])^(a[121] & b[120])^(a[120] & b[121])^(a[119] & b[122])^(a[118] & b[123])^(a[117] & b[124])^(a[116] & b[125])^(a[115] & b[126])^(a[114] & b[127])^(a[113] & b[128])^(a[112] & b[129])^(a[111] & b[130])^(a[110] & b[131])^(a[109] & b[132])^(a[108] & b[133])^(a[107] & b[134])^(a[106] & b[135])^(a[105] & b[136])^(a[104] & b[137])^(a[103] & b[138])^(a[102] & b[139])^(a[101] & b[140])^(a[100] & b[141])^(a[99] & b[142])^(a[98] & b[143])^(a[97] & b[144])^(a[96] & b[145])^(a[95] & b[146])^(a[94] & b[147])^(a[93] & b[148])^(a[92] & b[149])^(a[91] & b[150])^(a[90] & b[151])^(a[89] & b[152])^(a[88] & b[153])^(a[87] & b[154])^(a[86] & b[155])^(a[85] & b[156])^(a[84] & b[157])^(a[83] & b[158])^(a[82] & b[159])^(a[81] & b[160])^(a[80] & b[161])^(a[79] & b[162]);
assign y[242] = (a[162] & b[80])^(a[161] & b[81])^(a[160] & b[82])^(a[159] & b[83])^(a[158] & b[84])^(a[157] & b[85])^(a[156] & b[86])^(a[155] & b[87])^(a[154] & b[88])^(a[153] & b[89])^(a[152] & b[90])^(a[151] & b[91])^(a[150] & b[92])^(a[149] & b[93])^(a[148] & b[94])^(a[147] & b[95])^(a[146] & b[96])^(a[145] & b[97])^(a[144] & b[98])^(a[143] & b[99])^(a[142] & b[100])^(a[141] & b[101])^(a[140] & b[102])^(a[139] & b[103])^(a[138] & b[104])^(a[137] & b[105])^(a[136] & b[106])^(a[135] & b[107])^(a[134] & b[108])^(a[133] & b[109])^(a[132] & b[110])^(a[131] & b[111])^(a[130] & b[112])^(a[129] & b[113])^(a[128] & b[114])^(a[127] & b[115])^(a[126] & b[116])^(a[125] & b[117])^(a[124] & b[118])^(a[123] & b[119])^(a[122] & b[120])^(a[121] & b[121])^(a[120] & b[122])^(a[119] & b[123])^(a[118] & b[124])^(a[117] & b[125])^(a[116] & b[126])^(a[115] & b[127])^(a[114] & b[128])^(a[113] & b[129])^(a[112] & b[130])^(a[111] & b[131])^(a[110] & b[132])^(a[109] & b[133])^(a[108] & b[134])^(a[107] & b[135])^(a[106] & b[136])^(a[105] & b[137])^(a[104] & b[138])^(a[103] & b[139])^(a[102] & b[140])^(a[101] & b[141])^(a[100] & b[142])^(a[99] & b[143])^(a[98] & b[144])^(a[97] & b[145])^(a[96] & b[146])^(a[95] & b[147])^(a[94] & b[148])^(a[93] & b[149])^(a[92] & b[150])^(a[91] & b[151])^(a[90] & b[152])^(a[89] & b[153])^(a[88] & b[154])^(a[87] & b[155])^(a[86] & b[156])^(a[85] & b[157])^(a[84] & b[158])^(a[83] & b[159])^(a[82] & b[160])^(a[81] & b[161])^(a[80] & b[162]);
assign y[243] = (a[162] & b[81])^(a[161] & b[82])^(a[160] & b[83])^(a[159] & b[84])^(a[158] & b[85])^(a[157] & b[86])^(a[156] & b[87])^(a[155] & b[88])^(a[154] & b[89])^(a[153] & b[90])^(a[152] & b[91])^(a[151] & b[92])^(a[150] & b[93])^(a[149] & b[94])^(a[148] & b[95])^(a[147] & b[96])^(a[146] & b[97])^(a[145] & b[98])^(a[144] & b[99])^(a[143] & b[100])^(a[142] & b[101])^(a[141] & b[102])^(a[140] & b[103])^(a[139] & b[104])^(a[138] & b[105])^(a[137] & b[106])^(a[136] & b[107])^(a[135] & b[108])^(a[134] & b[109])^(a[133] & b[110])^(a[132] & b[111])^(a[131] & b[112])^(a[130] & b[113])^(a[129] & b[114])^(a[128] & b[115])^(a[127] & b[116])^(a[126] & b[117])^(a[125] & b[118])^(a[124] & b[119])^(a[123] & b[120])^(a[122] & b[121])^(a[121] & b[122])^(a[120] & b[123])^(a[119] & b[124])^(a[118] & b[125])^(a[117] & b[126])^(a[116] & b[127])^(a[115] & b[128])^(a[114] & b[129])^(a[113] & b[130])^(a[112] & b[131])^(a[111] & b[132])^(a[110] & b[133])^(a[109] & b[134])^(a[108] & b[135])^(a[107] & b[136])^(a[106] & b[137])^(a[105] & b[138])^(a[104] & b[139])^(a[103] & b[140])^(a[102] & b[141])^(a[101] & b[142])^(a[100] & b[143])^(a[99] & b[144])^(a[98] & b[145])^(a[97] & b[146])^(a[96] & b[147])^(a[95] & b[148])^(a[94] & b[149])^(a[93] & b[150])^(a[92] & b[151])^(a[91] & b[152])^(a[90] & b[153])^(a[89] & b[154])^(a[88] & b[155])^(a[87] & b[156])^(a[86] & b[157])^(a[85] & b[158])^(a[84] & b[159])^(a[83] & b[160])^(a[82] & b[161])^(a[81] & b[162]);
assign y[244] = (a[162] & b[82])^(a[161] & b[83])^(a[160] & b[84])^(a[159] & b[85])^(a[158] & b[86])^(a[157] & b[87])^(a[156] & b[88])^(a[155] & b[89])^(a[154] & b[90])^(a[153] & b[91])^(a[152] & b[92])^(a[151] & b[93])^(a[150] & b[94])^(a[149] & b[95])^(a[148] & b[96])^(a[147] & b[97])^(a[146] & b[98])^(a[145] & b[99])^(a[144] & b[100])^(a[143] & b[101])^(a[142] & b[102])^(a[141] & b[103])^(a[140] & b[104])^(a[139] & b[105])^(a[138] & b[106])^(a[137] & b[107])^(a[136] & b[108])^(a[135] & b[109])^(a[134] & b[110])^(a[133] & b[111])^(a[132] & b[112])^(a[131] & b[113])^(a[130] & b[114])^(a[129] & b[115])^(a[128] & b[116])^(a[127] & b[117])^(a[126] & b[118])^(a[125] & b[119])^(a[124] & b[120])^(a[123] & b[121])^(a[122] & b[122])^(a[121] & b[123])^(a[120] & b[124])^(a[119] & b[125])^(a[118] & b[126])^(a[117] & b[127])^(a[116] & b[128])^(a[115] & b[129])^(a[114] & b[130])^(a[113] & b[131])^(a[112] & b[132])^(a[111] & b[133])^(a[110] & b[134])^(a[109] & b[135])^(a[108] & b[136])^(a[107] & b[137])^(a[106] & b[138])^(a[105] & b[139])^(a[104] & b[140])^(a[103] & b[141])^(a[102] & b[142])^(a[101] & b[143])^(a[100] & b[144])^(a[99] & b[145])^(a[98] & b[146])^(a[97] & b[147])^(a[96] & b[148])^(a[95] & b[149])^(a[94] & b[150])^(a[93] & b[151])^(a[92] & b[152])^(a[91] & b[153])^(a[90] & b[154])^(a[89] & b[155])^(a[88] & b[156])^(a[87] & b[157])^(a[86] & b[158])^(a[85] & b[159])^(a[84] & b[160])^(a[83] & b[161])^(a[82] & b[162]);
assign y[245] = (a[162] & b[83])^(a[161] & b[84])^(a[160] & b[85])^(a[159] & b[86])^(a[158] & b[87])^(a[157] & b[88])^(a[156] & b[89])^(a[155] & b[90])^(a[154] & b[91])^(a[153] & b[92])^(a[152] & b[93])^(a[151] & b[94])^(a[150] & b[95])^(a[149] & b[96])^(a[148] & b[97])^(a[147] & b[98])^(a[146] & b[99])^(a[145] & b[100])^(a[144] & b[101])^(a[143] & b[102])^(a[142] & b[103])^(a[141] & b[104])^(a[140] & b[105])^(a[139] & b[106])^(a[138] & b[107])^(a[137] & b[108])^(a[136] & b[109])^(a[135] & b[110])^(a[134] & b[111])^(a[133] & b[112])^(a[132] & b[113])^(a[131] & b[114])^(a[130] & b[115])^(a[129] & b[116])^(a[128] & b[117])^(a[127] & b[118])^(a[126] & b[119])^(a[125] & b[120])^(a[124] & b[121])^(a[123] & b[122])^(a[122] & b[123])^(a[121] & b[124])^(a[120] & b[125])^(a[119] & b[126])^(a[118] & b[127])^(a[117] & b[128])^(a[116] & b[129])^(a[115] & b[130])^(a[114] & b[131])^(a[113] & b[132])^(a[112] & b[133])^(a[111] & b[134])^(a[110] & b[135])^(a[109] & b[136])^(a[108] & b[137])^(a[107] & b[138])^(a[106] & b[139])^(a[105] & b[140])^(a[104] & b[141])^(a[103] & b[142])^(a[102] & b[143])^(a[101] & b[144])^(a[100] & b[145])^(a[99] & b[146])^(a[98] & b[147])^(a[97] & b[148])^(a[96] & b[149])^(a[95] & b[150])^(a[94] & b[151])^(a[93] & b[152])^(a[92] & b[153])^(a[91] & b[154])^(a[90] & b[155])^(a[89] & b[156])^(a[88] & b[157])^(a[87] & b[158])^(a[86] & b[159])^(a[85] & b[160])^(a[84] & b[161])^(a[83] & b[162]);
assign y[246] = (a[162] & b[84])^(a[161] & b[85])^(a[160] & b[86])^(a[159] & b[87])^(a[158] & b[88])^(a[157] & b[89])^(a[156] & b[90])^(a[155] & b[91])^(a[154] & b[92])^(a[153] & b[93])^(a[152] & b[94])^(a[151] & b[95])^(a[150] & b[96])^(a[149] & b[97])^(a[148] & b[98])^(a[147] & b[99])^(a[146] & b[100])^(a[145] & b[101])^(a[144] & b[102])^(a[143] & b[103])^(a[142] & b[104])^(a[141] & b[105])^(a[140] & b[106])^(a[139] & b[107])^(a[138] & b[108])^(a[137] & b[109])^(a[136] & b[110])^(a[135] & b[111])^(a[134] & b[112])^(a[133] & b[113])^(a[132] & b[114])^(a[131] & b[115])^(a[130] & b[116])^(a[129] & b[117])^(a[128] & b[118])^(a[127] & b[119])^(a[126] & b[120])^(a[125] & b[121])^(a[124] & b[122])^(a[123] & b[123])^(a[122] & b[124])^(a[121] & b[125])^(a[120] & b[126])^(a[119] & b[127])^(a[118] & b[128])^(a[117] & b[129])^(a[116] & b[130])^(a[115] & b[131])^(a[114] & b[132])^(a[113] & b[133])^(a[112] & b[134])^(a[111] & b[135])^(a[110] & b[136])^(a[109] & b[137])^(a[108] & b[138])^(a[107] & b[139])^(a[106] & b[140])^(a[105] & b[141])^(a[104] & b[142])^(a[103] & b[143])^(a[102] & b[144])^(a[101] & b[145])^(a[100] & b[146])^(a[99] & b[147])^(a[98] & b[148])^(a[97] & b[149])^(a[96] & b[150])^(a[95] & b[151])^(a[94] & b[152])^(a[93] & b[153])^(a[92] & b[154])^(a[91] & b[155])^(a[90] & b[156])^(a[89] & b[157])^(a[88] & b[158])^(a[87] & b[159])^(a[86] & b[160])^(a[85] & b[161])^(a[84] & b[162]);
assign y[247] = (a[162] & b[85])^(a[161] & b[86])^(a[160] & b[87])^(a[159] & b[88])^(a[158] & b[89])^(a[157] & b[90])^(a[156] & b[91])^(a[155] & b[92])^(a[154] & b[93])^(a[153] & b[94])^(a[152] & b[95])^(a[151] & b[96])^(a[150] & b[97])^(a[149] & b[98])^(a[148] & b[99])^(a[147] & b[100])^(a[146] & b[101])^(a[145] & b[102])^(a[144] & b[103])^(a[143] & b[104])^(a[142] & b[105])^(a[141] & b[106])^(a[140] & b[107])^(a[139] & b[108])^(a[138] & b[109])^(a[137] & b[110])^(a[136] & b[111])^(a[135] & b[112])^(a[134] & b[113])^(a[133] & b[114])^(a[132] & b[115])^(a[131] & b[116])^(a[130] & b[117])^(a[129] & b[118])^(a[128] & b[119])^(a[127] & b[120])^(a[126] & b[121])^(a[125] & b[122])^(a[124] & b[123])^(a[123] & b[124])^(a[122] & b[125])^(a[121] & b[126])^(a[120] & b[127])^(a[119] & b[128])^(a[118] & b[129])^(a[117] & b[130])^(a[116] & b[131])^(a[115] & b[132])^(a[114] & b[133])^(a[113] & b[134])^(a[112] & b[135])^(a[111] & b[136])^(a[110] & b[137])^(a[109] & b[138])^(a[108] & b[139])^(a[107] & b[140])^(a[106] & b[141])^(a[105] & b[142])^(a[104] & b[143])^(a[103] & b[144])^(a[102] & b[145])^(a[101] & b[146])^(a[100] & b[147])^(a[99] & b[148])^(a[98] & b[149])^(a[97] & b[150])^(a[96] & b[151])^(a[95] & b[152])^(a[94] & b[153])^(a[93] & b[154])^(a[92] & b[155])^(a[91] & b[156])^(a[90] & b[157])^(a[89] & b[158])^(a[88] & b[159])^(a[87] & b[160])^(a[86] & b[161])^(a[85] & b[162]);
assign y[248] = (a[162] & b[86])^(a[161] & b[87])^(a[160] & b[88])^(a[159] & b[89])^(a[158] & b[90])^(a[157] & b[91])^(a[156] & b[92])^(a[155] & b[93])^(a[154] & b[94])^(a[153] & b[95])^(a[152] & b[96])^(a[151] & b[97])^(a[150] & b[98])^(a[149] & b[99])^(a[148] & b[100])^(a[147] & b[101])^(a[146] & b[102])^(a[145] & b[103])^(a[144] & b[104])^(a[143] & b[105])^(a[142] & b[106])^(a[141] & b[107])^(a[140] & b[108])^(a[139] & b[109])^(a[138] & b[110])^(a[137] & b[111])^(a[136] & b[112])^(a[135] & b[113])^(a[134] & b[114])^(a[133] & b[115])^(a[132] & b[116])^(a[131] & b[117])^(a[130] & b[118])^(a[129] & b[119])^(a[128] & b[120])^(a[127] & b[121])^(a[126] & b[122])^(a[125] & b[123])^(a[124] & b[124])^(a[123] & b[125])^(a[122] & b[126])^(a[121] & b[127])^(a[120] & b[128])^(a[119] & b[129])^(a[118] & b[130])^(a[117] & b[131])^(a[116] & b[132])^(a[115] & b[133])^(a[114] & b[134])^(a[113] & b[135])^(a[112] & b[136])^(a[111] & b[137])^(a[110] & b[138])^(a[109] & b[139])^(a[108] & b[140])^(a[107] & b[141])^(a[106] & b[142])^(a[105] & b[143])^(a[104] & b[144])^(a[103] & b[145])^(a[102] & b[146])^(a[101] & b[147])^(a[100] & b[148])^(a[99] & b[149])^(a[98] & b[150])^(a[97] & b[151])^(a[96] & b[152])^(a[95] & b[153])^(a[94] & b[154])^(a[93] & b[155])^(a[92] & b[156])^(a[91] & b[157])^(a[90] & b[158])^(a[89] & b[159])^(a[88] & b[160])^(a[87] & b[161])^(a[86] & b[162]);
assign y[249] = (a[162] & b[87])^(a[161] & b[88])^(a[160] & b[89])^(a[159] & b[90])^(a[158] & b[91])^(a[157] & b[92])^(a[156] & b[93])^(a[155] & b[94])^(a[154] & b[95])^(a[153] & b[96])^(a[152] & b[97])^(a[151] & b[98])^(a[150] & b[99])^(a[149] & b[100])^(a[148] & b[101])^(a[147] & b[102])^(a[146] & b[103])^(a[145] & b[104])^(a[144] & b[105])^(a[143] & b[106])^(a[142] & b[107])^(a[141] & b[108])^(a[140] & b[109])^(a[139] & b[110])^(a[138] & b[111])^(a[137] & b[112])^(a[136] & b[113])^(a[135] & b[114])^(a[134] & b[115])^(a[133] & b[116])^(a[132] & b[117])^(a[131] & b[118])^(a[130] & b[119])^(a[129] & b[120])^(a[128] & b[121])^(a[127] & b[122])^(a[126] & b[123])^(a[125] & b[124])^(a[124] & b[125])^(a[123] & b[126])^(a[122] & b[127])^(a[121] & b[128])^(a[120] & b[129])^(a[119] & b[130])^(a[118] & b[131])^(a[117] & b[132])^(a[116] & b[133])^(a[115] & b[134])^(a[114] & b[135])^(a[113] & b[136])^(a[112] & b[137])^(a[111] & b[138])^(a[110] & b[139])^(a[109] & b[140])^(a[108] & b[141])^(a[107] & b[142])^(a[106] & b[143])^(a[105] & b[144])^(a[104] & b[145])^(a[103] & b[146])^(a[102] & b[147])^(a[101] & b[148])^(a[100] & b[149])^(a[99] & b[150])^(a[98] & b[151])^(a[97] & b[152])^(a[96] & b[153])^(a[95] & b[154])^(a[94] & b[155])^(a[93] & b[156])^(a[92] & b[157])^(a[91] & b[158])^(a[90] & b[159])^(a[89] & b[160])^(a[88] & b[161])^(a[87] & b[162]);
assign y[250] = (a[162] & b[88])^(a[161] & b[89])^(a[160] & b[90])^(a[159] & b[91])^(a[158] & b[92])^(a[157] & b[93])^(a[156] & b[94])^(a[155] & b[95])^(a[154] & b[96])^(a[153] & b[97])^(a[152] & b[98])^(a[151] & b[99])^(a[150] & b[100])^(a[149] & b[101])^(a[148] & b[102])^(a[147] & b[103])^(a[146] & b[104])^(a[145] & b[105])^(a[144] & b[106])^(a[143] & b[107])^(a[142] & b[108])^(a[141] & b[109])^(a[140] & b[110])^(a[139] & b[111])^(a[138] & b[112])^(a[137] & b[113])^(a[136] & b[114])^(a[135] & b[115])^(a[134] & b[116])^(a[133] & b[117])^(a[132] & b[118])^(a[131] & b[119])^(a[130] & b[120])^(a[129] & b[121])^(a[128] & b[122])^(a[127] & b[123])^(a[126] & b[124])^(a[125] & b[125])^(a[124] & b[126])^(a[123] & b[127])^(a[122] & b[128])^(a[121] & b[129])^(a[120] & b[130])^(a[119] & b[131])^(a[118] & b[132])^(a[117] & b[133])^(a[116] & b[134])^(a[115] & b[135])^(a[114] & b[136])^(a[113] & b[137])^(a[112] & b[138])^(a[111] & b[139])^(a[110] & b[140])^(a[109] & b[141])^(a[108] & b[142])^(a[107] & b[143])^(a[106] & b[144])^(a[105] & b[145])^(a[104] & b[146])^(a[103] & b[147])^(a[102] & b[148])^(a[101] & b[149])^(a[100] & b[150])^(a[99] & b[151])^(a[98] & b[152])^(a[97] & b[153])^(a[96] & b[154])^(a[95] & b[155])^(a[94] & b[156])^(a[93] & b[157])^(a[92] & b[158])^(a[91] & b[159])^(a[90] & b[160])^(a[89] & b[161])^(a[88] & b[162]);
assign y[251] = (a[162] & b[89])^(a[161] & b[90])^(a[160] & b[91])^(a[159] & b[92])^(a[158] & b[93])^(a[157] & b[94])^(a[156] & b[95])^(a[155] & b[96])^(a[154] & b[97])^(a[153] & b[98])^(a[152] & b[99])^(a[151] & b[100])^(a[150] & b[101])^(a[149] & b[102])^(a[148] & b[103])^(a[147] & b[104])^(a[146] & b[105])^(a[145] & b[106])^(a[144] & b[107])^(a[143] & b[108])^(a[142] & b[109])^(a[141] & b[110])^(a[140] & b[111])^(a[139] & b[112])^(a[138] & b[113])^(a[137] & b[114])^(a[136] & b[115])^(a[135] & b[116])^(a[134] & b[117])^(a[133] & b[118])^(a[132] & b[119])^(a[131] & b[120])^(a[130] & b[121])^(a[129] & b[122])^(a[128] & b[123])^(a[127] & b[124])^(a[126] & b[125])^(a[125] & b[126])^(a[124] & b[127])^(a[123] & b[128])^(a[122] & b[129])^(a[121] & b[130])^(a[120] & b[131])^(a[119] & b[132])^(a[118] & b[133])^(a[117] & b[134])^(a[116] & b[135])^(a[115] & b[136])^(a[114] & b[137])^(a[113] & b[138])^(a[112] & b[139])^(a[111] & b[140])^(a[110] & b[141])^(a[109] & b[142])^(a[108] & b[143])^(a[107] & b[144])^(a[106] & b[145])^(a[105] & b[146])^(a[104] & b[147])^(a[103] & b[148])^(a[102] & b[149])^(a[101] & b[150])^(a[100] & b[151])^(a[99] & b[152])^(a[98] & b[153])^(a[97] & b[154])^(a[96] & b[155])^(a[95] & b[156])^(a[94] & b[157])^(a[93] & b[158])^(a[92] & b[159])^(a[91] & b[160])^(a[90] & b[161])^(a[89] & b[162]);
assign y[252] = (a[162] & b[90])^(a[161] & b[91])^(a[160] & b[92])^(a[159] & b[93])^(a[158] & b[94])^(a[157] & b[95])^(a[156] & b[96])^(a[155] & b[97])^(a[154] & b[98])^(a[153] & b[99])^(a[152] & b[100])^(a[151] & b[101])^(a[150] & b[102])^(a[149] & b[103])^(a[148] & b[104])^(a[147] & b[105])^(a[146] & b[106])^(a[145] & b[107])^(a[144] & b[108])^(a[143] & b[109])^(a[142] & b[110])^(a[141] & b[111])^(a[140] & b[112])^(a[139] & b[113])^(a[138] & b[114])^(a[137] & b[115])^(a[136] & b[116])^(a[135] & b[117])^(a[134] & b[118])^(a[133] & b[119])^(a[132] & b[120])^(a[131] & b[121])^(a[130] & b[122])^(a[129] & b[123])^(a[128] & b[124])^(a[127] & b[125])^(a[126] & b[126])^(a[125] & b[127])^(a[124] & b[128])^(a[123] & b[129])^(a[122] & b[130])^(a[121] & b[131])^(a[120] & b[132])^(a[119] & b[133])^(a[118] & b[134])^(a[117] & b[135])^(a[116] & b[136])^(a[115] & b[137])^(a[114] & b[138])^(a[113] & b[139])^(a[112] & b[140])^(a[111] & b[141])^(a[110] & b[142])^(a[109] & b[143])^(a[108] & b[144])^(a[107] & b[145])^(a[106] & b[146])^(a[105] & b[147])^(a[104] & b[148])^(a[103] & b[149])^(a[102] & b[150])^(a[101] & b[151])^(a[100] & b[152])^(a[99] & b[153])^(a[98] & b[154])^(a[97] & b[155])^(a[96] & b[156])^(a[95] & b[157])^(a[94] & b[158])^(a[93] & b[159])^(a[92] & b[160])^(a[91] & b[161])^(a[90] & b[162]);
assign y[253] = (a[162] & b[91])^(a[161] & b[92])^(a[160] & b[93])^(a[159] & b[94])^(a[158] & b[95])^(a[157] & b[96])^(a[156] & b[97])^(a[155] & b[98])^(a[154] & b[99])^(a[153] & b[100])^(a[152] & b[101])^(a[151] & b[102])^(a[150] & b[103])^(a[149] & b[104])^(a[148] & b[105])^(a[147] & b[106])^(a[146] & b[107])^(a[145] & b[108])^(a[144] & b[109])^(a[143] & b[110])^(a[142] & b[111])^(a[141] & b[112])^(a[140] & b[113])^(a[139] & b[114])^(a[138] & b[115])^(a[137] & b[116])^(a[136] & b[117])^(a[135] & b[118])^(a[134] & b[119])^(a[133] & b[120])^(a[132] & b[121])^(a[131] & b[122])^(a[130] & b[123])^(a[129] & b[124])^(a[128] & b[125])^(a[127] & b[126])^(a[126] & b[127])^(a[125] & b[128])^(a[124] & b[129])^(a[123] & b[130])^(a[122] & b[131])^(a[121] & b[132])^(a[120] & b[133])^(a[119] & b[134])^(a[118] & b[135])^(a[117] & b[136])^(a[116] & b[137])^(a[115] & b[138])^(a[114] & b[139])^(a[113] & b[140])^(a[112] & b[141])^(a[111] & b[142])^(a[110] & b[143])^(a[109] & b[144])^(a[108] & b[145])^(a[107] & b[146])^(a[106] & b[147])^(a[105] & b[148])^(a[104] & b[149])^(a[103] & b[150])^(a[102] & b[151])^(a[101] & b[152])^(a[100] & b[153])^(a[99] & b[154])^(a[98] & b[155])^(a[97] & b[156])^(a[96] & b[157])^(a[95] & b[158])^(a[94] & b[159])^(a[93] & b[160])^(a[92] & b[161])^(a[91] & b[162]);
assign y[254] = (a[162] & b[92])^(a[161] & b[93])^(a[160] & b[94])^(a[159] & b[95])^(a[158] & b[96])^(a[157] & b[97])^(a[156] & b[98])^(a[155] & b[99])^(a[154] & b[100])^(a[153] & b[101])^(a[152] & b[102])^(a[151] & b[103])^(a[150] & b[104])^(a[149] & b[105])^(a[148] & b[106])^(a[147] & b[107])^(a[146] & b[108])^(a[145] & b[109])^(a[144] & b[110])^(a[143] & b[111])^(a[142] & b[112])^(a[141] & b[113])^(a[140] & b[114])^(a[139] & b[115])^(a[138] & b[116])^(a[137] & b[117])^(a[136] & b[118])^(a[135] & b[119])^(a[134] & b[120])^(a[133] & b[121])^(a[132] & b[122])^(a[131] & b[123])^(a[130] & b[124])^(a[129] & b[125])^(a[128] & b[126])^(a[127] & b[127])^(a[126] & b[128])^(a[125] & b[129])^(a[124] & b[130])^(a[123] & b[131])^(a[122] & b[132])^(a[121] & b[133])^(a[120] & b[134])^(a[119] & b[135])^(a[118] & b[136])^(a[117] & b[137])^(a[116] & b[138])^(a[115] & b[139])^(a[114] & b[140])^(a[113] & b[141])^(a[112] & b[142])^(a[111] & b[143])^(a[110] & b[144])^(a[109] & b[145])^(a[108] & b[146])^(a[107] & b[147])^(a[106] & b[148])^(a[105] & b[149])^(a[104] & b[150])^(a[103] & b[151])^(a[102] & b[152])^(a[101] & b[153])^(a[100] & b[154])^(a[99] & b[155])^(a[98] & b[156])^(a[97] & b[157])^(a[96] & b[158])^(a[95] & b[159])^(a[94] & b[160])^(a[93] & b[161])^(a[92] & b[162]);
assign y[255] = (a[162] & b[93])^(a[161] & b[94])^(a[160] & b[95])^(a[159] & b[96])^(a[158] & b[97])^(a[157] & b[98])^(a[156] & b[99])^(a[155] & b[100])^(a[154] & b[101])^(a[153] & b[102])^(a[152] & b[103])^(a[151] & b[104])^(a[150] & b[105])^(a[149] & b[106])^(a[148] & b[107])^(a[147] & b[108])^(a[146] & b[109])^(a[145] & b[110])^(a[144] & b[111])^(a[143] & b[112])^(a[142] & b[113])^(a[141] & b[114])^(a[140] & b[115])^(a[139] & b[116])^(a[138] & b[117])^(a[137] & b[118])^(a[136] & b[119])^(a[135] & b[120])^(a[134] & b[121])^(a[133] & b[122])^(a[132] & b[123])^(a[131] & b[124])^(a[130] & b[125])^(a[129] & b[126])^(a[128] & b[127])^(a[127] & b[128])^(a[126] & b[129])^(a[125] & b[130])^(a[124] & b[131])^(a[123] & b[132])^(a[122] & b[133])^(a[121] & b[134])^(a[120] & b[135])^(a[119] & b[136])^(a[118] & b[137])^(a[117] & b[138])^(a[116] & b[139])^(a[115] & b[140])^(a[114] & b[141])^(a[113] & b[142])^(a[112] & b[143])^(a[111] & b[144])^(a[110] & b[145])^(a[109] & b[146])^(a[108] & b[147])^(a[107] & b[148])^(a[106] & b[149])^(a[105] & b[150])^(a[104] & b[151])^(a[103] & b[152])^(a[102] & b[153])^(a[101] & b[154])^(a[100] & b[155])^(a[99] & b[156])^(a[98] & b[157])^(a[97] & b[158])^(a[96] & b[159])^(a[95] & b[160])^(a[94] & b[161])^(a[93] & b[162]);
assign y[256] = (a[162] & b[94])^(a[161] & b[95])^(a[160] & b[96])^(a[159] & b[97])^(a[158] & b[98])^(a[157] & b[99])^(a[156] & b[100])^(a[155] & b[101])^(a[154] & b[102])^(a[153] & b[103])^(a[152] & b[104])^(a[151] & b[105])^(a[150] & b[106])^(a[149] & b[107])^(a[148] & b[108])^(a[147] & b[109])^(a[146] & b[110])^(a[145] & b[111])^(a[144] & b[112])^(a[143] & b[113])^(a[142] & b[114])^(a[141] & b[115])^(a[140] & b[116])^(a[139] & b[117])^(a[138] & b[118])^(a[137] & b[119])^(a[136] & b[120])^(a[135] & b[121])^(a[134] & b[122])^(a[133] & b[123])^(a[132] & b[124])^(a[131] & b[125])^(a[130] & b[126])^(a[129] & b[127])^(a[128] & b[128])^(a[127] & b[129])^(a[126] & b[130])^(a[125] & b[131])^(a[124] & b[132])^(a[123] & b[133])^(a[122] & b[134])^(a[121] & b[135])^(a[120] & b[136])^(a[119] & b[137])^(a[118] & b[138])^(a[117] & b[139])^(a[116] & b[140])^(a[115] & b[141])^(a[114] & b[142])^(a[113] & b[143])^(a[112] & b[144])^(a[111] & b[145])^(a[110] & b[146])^(a[109] & b[147])^(a[108] & b[148])^(a[107] & b[149])^(a[106] & b[150])^(a[105] & b[151])^(a[104] & b[152])^(a[103] & b[153])^(a[102] & b[154])^(a[101] & b[155])^(a[100] & b[156])^(a[99] & b[157])^(a[98] & b[158])^(a[97] & b[159])^(a[96] & b[160])^(a[95] & b[161])^(a[94] & b[162]);
assign y[257] = (a[162] & b[95])^(a[161] & b[96])^(a[160] & b[97])^(a[159] & b[98])^(a[158] & b[99])^(a[157] & b[100])^(a[156] & b[101])^(a[155] & b[102])^(a[154] & b[103])^(a[153] & b[104])^(a[152] & b[105])^(a[151] & b[106])^(a[150] & b[107])^(a[149] & b[108])^(a[148] & b[109])^(a[147] & b[110])^(a[146] & b[111])^(a[145] & b[112])^(a[144] & b[113])^(a[143] & b[114])^(a[142] & b[115])^(a[141] & b[116])^(a[140] & b[117])^(a[139] & b[118])^(a[138] & b[119])^(a[137] & b[120])^(a[136] & b[121])^(a[135] & b[122])^(a[134] & b[123])^(a[133] & b[124])^(a[132] & b[125])^(a[131] & b[126])^(a[130] & b[127])^(a[129] & b[128])^(a[128] & b[129])^(a[127] & b[130])^(a[126] & b[131])^(a[125] & b[132])^(a[124] & b[133])^(a[123] & b[134])^(a[122] & b[135])^(a[121] & b[136])^(a[120] & b[137])^(a[119] & b[138])^(a[118] & b[139])^(a[117] & b[140])^(a[116] & b[141])^(a[115] & b[142])^(a[114] & b[143])^(a[113] & b[144])^(a[112] & b[145])^(a[111] & b[146])^(a[110] & b[147])^(a[109] & b[148])^(a[108] & b[149])^(a[107] & b[150])^(a[106] & b[151])^(a[105] & b[152])^(a[104] & b[153])^(a[103] & b[154])^(a[102] & b[155])^(a[101] & b[156])^(a[100] & b[157])^(a[99] & b[158])^(a[98] & b[159])^(a[97] & b[160])^(a[96] & b[161])^(a[95] & b[162]);
assign y[258] = (a[162] & b[96])^(a[161] & b[97])^(a[160] & b[98])^(a[159] & b[99])^(a[158] & b[100])^(a[157] & b[101])^(a[156] & b[102])^(a[155] & b[103])^(a[154] & b[104])^(a[153] & b[105])^(a[152] & b[106])^(a[151] & b[107])^(a[150] & b[108])^(a[149] & b[109])^(a[148] & b[110])^(a[147] & b[111])^(a[146] & b[112])^(a[145] & b[113])^(a[144] & b[114])^(a[143] & b[115])^(a[142] & b[116])^(a[141] & b[117])^(a[140] & b[118])^(a[139] & b[119])^(a[138] & b[120])^(a[137] & b[121])^(a[136] & b[122])^(a[135] & b[123])^(a[134] & b[124])^(a[133] & b[125])^(a[132] & b[126])^(a[131] & b[127])^(a[130] & b[128])^(a[129] & b[129])^(a[128] & b[130])^(a[127] & b[131])^(a[126] & b[132])^(a[125] & b[133])^(a[124] & b[134])^(a[123] & b[135])^(a[122] & b[136])^(a[121] & b[137])^(a[120] & b[138])^(a[119] & b[139])^(a[118] & b[140])^(a[117] & b[141])^(a[116] & b[142])^(a[115] & b[143])^(a[114] & b[144])^(a[113] & b[145])^(a[112] & b[146])^(a[111] & b[147])^(a[110] & b[148])^(a[109] & b[149])^(a[108] & b[150])^(a[107] & b[151])^(a[106] & b[152])^(a[105] & b[153])^(a[104] & b[154])^(a[103] & b[155])^(a[102] & b[156])^(a[101] & b[157])^(a[100] & b[158])^(a[99] & b[159])^(a[98] & b[160])^(a[97] & b[161])^(a[96] & b[162]);
assign y[259] = (a[162] & b[97])^(a[161] & b[98])^(a[160] & b[99])^(a[159] & b[100])^(a[158] & b[101])^(a[157] & b[102])^(a[156] & b[103])^(a[155] & b[104])^(a[154] & b[105])^(a[153] & b[106])^(a[152] & b[107])^(a[151] & b[108])^(a[150] & b[109])^(a[149] & b[110])^(a[148] & b[111])^(a[147] & b[112])^(a[146] & b[113])^(a[145] & b[114])^(a[144] & b[115])^(a[143] & b[116])^(a[142] & b[117])^(a[141] & b[118])^(a[140] & b[119])^(a[139] & b[120])^(a[138] & b[121])^(a[137] & b[122])^(a[136] & b[123])^(a[135] & b[124])^(a[134] & b[125])^(a[133] & b[126])^(a[132] & b[127])^(a[131] & b[128])^(a[130] & b[129])^(a[129] & b[130])^(a[128] & b[131])^(a[127] & b[132])^(a[126] & b[133])^(a[125] & b[134])^(a[124] & b[135])^(a[123] & b[136])^(a[122] & b[137])^(a[121] & b[138])^(a[120] & b[139])^(a[119] & b[140])^(a[118] & b[141])^(a[117] & b[142])^(a[116] & b[143])^(a[115] & b[144])^(a[114] & b[145])^(a[113] & b[146])^(a[112] & b[147])^(a[111] & b[148])^(a[110] & b[149])^(a[109] & b[150])^(a[108] & b[151])^(a[107] & b[152])^(a[106] & b[153])^(a[105] & b[154])^(a[104] & b[155])^(a[103] & b[156])^(a[102] & b[157])^(a[101] & b[158])^(a[100] & b[159])^(a[99] & b[160])^(a[98] & b[161])^(a[97] & b[162]);
assign y[260] = (a[162] & b[98])^(a[161] & b[99])^(a[160] & b[100])^(a[159] & b[101])^(a[158] & b[102])^(a[157] & b[103])^(a[156] & b[104])^(a[155] & b[105])^(a[154] & b[106])^(a[153] & b[107])^(a[152] & b[108])^(a[151] & b[109])^(a[150] & b[110])^(a[149] & b[111])^(a[148] & b[112])^(a[147] & b[113])^(a[146] & b[114])^(a[145] & b[115])^(a[144] & b[116])^(a[143] & b[117])^(a[142] & b[118])^(a[141] & b[119])^(a[140] & b[120])^(a[139] & b[121])^(a[138] & b[122])^(a[137] & b[123])^(a[136] & b[124])^(a[135] & b[125])^(a[134] & b[126])^(a[133] & b[127])^(a[132] & b[128])^(a[131] & b[129])^(a[130] & b[130])^(a[129] & b[131])^(a[128] & b[132])^(a[127] & b[133])^(a[126] & b[134])^(a[125] & b[135])^(a[124] & b[136])^(a[123] & b[137])^(a[122] & b[138])^(a[121] & b[139])^(a[120] & b[140])^(a[119] & b[141])^(a[118] & b[142])^(a[117] & b[143])^(a[116] & b[144])^(a[115] & b[145])^(a[114] & b[146])^(a[113] & b[147])^(a[112] & b[148])^(a[111] & b[149])^(a[110] & b[150])^(a[109] & b[151])^(a[108] & b[152])^(a[107] & b[153])^(a[106] & b[154])^(a[105] & b[155])^(a[104] & b[156])^(a[103] & b[157])^(a[102] & b[158])^(a[101] & b[159])^(a[100] & b[160])^(a[99] & b[161])^(a[98] & b[162]);
assign y[261] = (a[162] & b[99])^(a[161] & b[100])^(a[160] & b[101])^(a[159] & b[102])^(a[158] & b[103])^(a[157] & b[104])^(a[156] & b[105])^(a[155] & b[106])^(a[154] & b[107])^(a[153] & b[108])^(a[152] & b[109])^(a[151] & b[110])^(a[150] & b[111])^(a[149] & b[112])^(a[148] & b[113])^(a[147] & b[114])^(a[146] & b[115])^(a[145] & b[116])^(a[144] & b[117])^(a[143] & b[118])^(a[142] & b[119])^(a[141] & b[120])^(a[140] & b[121])^(a[139] & b[122])^(a[138] & b[123])^(a[137] & b[124])^(a[136] & b[125])^(a[135] & b[126])^(a[134] & b[127])^(a[133] & b[128])^(a[132] & b[129])^(a[131] & b[130])^(a[130] & b[131])^(a[129] & b[132])^(a[128] & b[133])^(a[127] & b[134])^(a[126] & b[135])^(a[125] & b[136])^(a[124] & b[137])^(a[123] & b[138])^(a[122] & b[139])^(a[121] & b[140])^(a[120] & b[141])^(a[119] & b[142])^(a[118] & b[143])^(a[117] & b[144])^(a[116] & b[145])^(a[115] & b[146])^(a[114] & b[147])^(a[113] & b[148])^(a[112] & b[149])^(a[111] & b[150])^(a[110] & b[151])^(a[109] & b[152])^(a[108] & b[153])^(a[107] & b[154])^(a[106] & b[155])^(a[105] & b[156])^(a[104] & b[157])^(a[103] & b[158])^(a[102] & b[159])^(a[101] & b[160])^(a[100] & b[161])^(a[99] & b[162]);
assign y[262] = (a[162] & b[100])^(a[161] & b[101])^(a[160] & b[102])^(a[159] & b[103])^(a[158] & b[104])^(a[157] & b[105])^(a[156] & b[106])^(a[155] & b[107])^(a[154] & b[108])^(a[153] & b[109])^(a[152] & b[110])^(a[151] & b[111])^(a[150] & b[112])^(a[149] & b[113])^(a[148] & b[114])^(a[147] & b[115])^(a[146] & b[116])^(a[145] & b[117])^(a[144] & b[118])^(a[143] & b[119])^(a[142] & b[120])^(a[141] & b[121])^(a[140] & b[122])^(a[139] & b[123])^(a[138] & b[124])^(a[137] & b[125])^(a[136] & b[126])^(a[135] & b[127])^(a[134] & b[128])^(a[133] & b[129])^(a[132] & b[130])^(a[131] & b[131])^(a[130] & b[132])^(a[129] & b[133])^(a[128] & b[134])^(a[127] & b[135])^(a[126] & b[136])^(a[125] & b[137])^(a[124] & b[138])^(a[123] & b[139])^(a[122] & b[140])^(a[121] & b[141])^(a[120] & b[142])^(a[119] & b[143])^(a[118] & b[144])^(a[117] & b[145])^(a[116] & b[146])^(a[115] & b[147])^(a[114] & b[148])^(a[113] & b[149])^(a[112] & b[150])^(a[111] & b[151])^(a[110] & b[152])^(a[109] & b[153])^(a[108] & b[154])^(a[107] & b[155])^(a[106] & b[156])^(a[105] & b[157])^(a[104] & b[158])^(a[103] & b[159])^(a[102] & b[160])^(a[101] & b[161])^(a[100] & b[162]);
assign y[263] = (a[162] & b[101])^(a[161] & b[102])^(a[160] & b[103])^(a[159] & b[104])^(a[158] & b[105])^(a[157] & b[106])^(a[156] & b[107])^(a[155] & b[108])^(a[154] & b[109])^(a[153] & b[110])^(a[152] & b[111])^(a[151] & b[112])^(a[150] & b[113])^(a[149] & b[114])^(a[148] & b[115])^(a[147] & b[116])^(a[146] & b[117])^(a[145] & b[118])^(a[144] & b[119])^(a[143] & b[120])^(a[142] & b[121])^(a[141] & b[122])^(a[140] & b[123])^(a[139] & b[124])^(a[138] & b[125])^(a[137] & b[126])^(a[136] & b[127])^(a[135] & b[128])^(a[134] & b[129])^(a[133] & b[130])^(a[132] & b[131])^(a[131] & b[132])^(a[130] & b[133])^(a[129] & b[134])^(a[128] & b[135])^(a[127] & b[136])^(a[126] & b[137])^(a[125] & b[138])^(a[124] & b[139])^(a[123] & b[140])^(a[122] & b[141])^(a[121] & b[142])^(a[120] & b[143])^(a[119] & b[144])^(a[118] & b[145])^(a[117] & b[146])^(a[116] & b[147])^(a[115] & b[148])^(a[114] & b[149])^(a[113] & b[150])^(a[112] & b[151])^(a[111] & b[152])^(a[110] & b[153])^(a[109] & b[154])^(a[108] & b[155])^(a[107] & b[156])^(a[106] & b[157])^(a[105] & b[158])^(a[104] & b[159])^(a[103] & b[160])^(a[102] & b[161])^(a[101] & b[162]);
assign y[264] = (a[162] & b[102])^(a[161] & b[103])^(a[160] & b[104])^(a[159] & b[105])^(a[158] & b[106])^(a[157] & b[107])^(a[156] & b[108])^(a[155] & b[109])^(a[154] & b[110])^(a[153] & b[111])^(a[152] & b[112])^(a[151] & b[113])^(a[150] & b[114])^(a[149] & b[115])^(a[148] & b[116])^(a[147] & b[117])^(a[146] & b[118])^(a[145] & b[119])^(a[144] & b[120])^(a[143] & b[121])^(a[142] & b[122])^(a[141] & b[123])^(a[140] & b[124])^(a[139] & b[125])^(a[138] & b[126])^(a[137] & b[127])^(a[136] & b[128])^(a[135] & b[129])^(a[134] & b[130])^(a[133] & b[131])^(a[132] & b[132])^(a[131] & b[133])^(a[130] & b[134])^(a[129] & b[135])^(a[128] & b[136])^(a[127] & b[137])^(a[126] & b[138])^(a[125] & b[139])^(a[124] & b[140])^(a[123] & b[141])^(a[122] & b[142])^(a[121] & b[143])^(a[120] & b[144])^(a[119] & b[145])^(a[118] & b[146])^(a[117] & b[147])^(a[116] & b[148])^(a[115] & b[149])^(a[114] & b[150])^(a[113] & b[151])^(a[112] & b[152])^(a[111] & b[153])^(a[110] & b[154])^(a[109] & b[155])^(a[108] & b[156])^(a[107] & b[157])^(a[106] & b[158])^(a[105] & b[159])^(a[104] & b[160])^(a[103] & b[161])^(a[102] & b[162]);
assign y[265] = (a[162] & b[103])^(a[161] & b[104])^(a[160] & b[105])^(a[159] & b[106])^(a[158] & b[107])^(a[157] & b[108])^(a[156] & b[109])^(a[155] & b[110])^(a[154] & b[111])^(a[153] & b[112])^(a[152] & b[113])^(a[151] & b[114])^(a[150] & b[115])^(a[149] & b[116])^(a[148] & b[117])^(a[147] & b[118])^(a[146] & b[119])^(a[145] & b[120])^(a[144] & b[121])^(a[143] & b[122])^(a[142] & b[123])^(a[141] & b[124])^(a[140] & b[125])^(a[139] & b[126])^(a[138] & b[127])^(a[137] & b[128])^(a[136] & b[129])^(a[135] & b[130])^(a[134] & b[131])^(a[133] & b[132])^(a[132] & b[133])^(a[131] & b[134])^(a[130] & b[135])^(a[129] & b[136])^(a[128] & b[137])^(a[127] & b[138])^(a[126] & b[139])^(a[125] & b[140])^(a[124] & b[141])^(a[123] & b[142])^(a[122] & b[143])^(a[121] & b[144])^(a[120] & b[145])^(a[119] & b[146])^(a[118] & b[147])^(a[117] & b[148])^(a[116] & b[149])^(a[115] & b[150])^(a[114] & b[151])^(a[113] & b[152])^(a[112] & b[153])^(a[111] & b[154])^(a[110] & b[155])^(a[109] & b[156])^(a[108] & b[157])^(a[107] & b[158])^(a[106] & b[159])^(a[105] & b[160])^(a[104] & b[161])^(a[103] & b[162]);
assign y[266] = (a[162] & b[104])^(a[161] & b[105])^(a[160] & b[106])^(a[159] & b[107])^(a[158] & b[108])^(a[157] & b[109])^(a[156] & b[110])^(a[155] & b[111])^(a[154] & b[112])^(a[153] & b[113])^(a[152] & b[114])^(a[151] & b[115])^(a[150] & b[116])^(a[149] & b[117])^(a[148] & b[118])^(a[147] & b[119])^(a[146] & b[120])^(a[145] & b[121])^(a[144] & b[122])^(a[143] & b[123])^(a[142] & b[124])^(a[141] & b[125])^(a[140] & b[126])^(a[139] & b[127])^(a[138] & b[128])^(a[137] & b[129])^(a[136] & b[130])^(a[135] & b[131])^(a[134] & b[132])^(a[133] & b[133])^(a[132] & b[134])^(a[131] & b[135])^(a[130] & b[136])^(a[129] & b[137])^(a[128] & b[138])^(a[127] & b[139])^(a[126] & b[140])^(a[125] & b[141])^(a[124] & b[142])^(a[123] & b[143])^(a[122] & b[144])^(a[121] & b[145])^(a[120] & b[146])^(a[119] & b[147])^(a[118] & b[148])^(a[117] & b[149])^(a[116] & b[150])^(a[115] & b[151])^(a[114] & b[152])^(a[113] & b[153])^(a[112] & b[154])^(a[111] & b[155])^(a[110] & b[156])^(a[109] & b[157])^(a[108] & b[158])^(a[107] & b[159])^(a[106] & b[160])^(a[105] & b[161])^(a[104] & b[162]);
assign y[267] = (a[162] & b[105])^(a[161] & b[106])^(a[160] & b[107])^(a[159] & b[108])^(a[158] & b[109])^(a[157] & b[110])^(a[156] & b[111])^(a[155] & b[112])^(a[154] & b[113])^(a[153] & b[114])^(a[152] & b[115])^(a[151] & b[116])^(a[150] & b[117])^(a[149] & b[118])^(a[148] & b[119])^(a[147] & b[120])^(a[146] & b[121])^(a[145] & b[122])^(a[144] & b[123])^(a[143] & b[124])^(a[142] & b[125])^(a[141] & b[126])^(a[140] & b[127])^(a[139] & b[128])^(a[138] & b[129])^(a[137] & b[130])^(a[136] & b[131])^(a[135] & b[132])^(a[134] & b[133])^(a[133] & b[134])^(a[132] & b[135])^(a[131] & b[136])^(a[130] & b[137])^(a[129] & b[138])^(a[128] & b[139])^(a[127] & b[140])^(a[126] & b[141])^(a[125] & b[142])^(a[124] & b[143])^(a[123] & b[144])^(a[122] & b[145])^(a[121] & b[146])^(a[120] & b[147])^(a[119] & b[148])^(a[118] & b[149])^(a[117] & b[150])^(a[116] & b[151])^(a[115] & b[152])^(a[114] & b[153])^(a[113] & b[154])^(a[112] & b[155])^(a[111] & b[156])^(a[110] & b[157])^(a[109] & b[158])^(a[108] & b[159])^(a[107] & b[160])^(a[106] & b[161])^(a[105] & b[162]);
assign y[268] = (a[162] & b[106])^(a[161] & b[107])^(a[160] & b[108])^(a[159] & b[109])^(a[158] & b[110])^(a[157] & b[111])^(a[156] & b[112])^(a[155] & b[113])^(a[154] & b[114])^(a[153] & b[115])^(a[152] & b[116])^(a[151] & b[117])^(a[150] & b[118])^(a[149] & b[119])^(a[148] & b[120])^(a[147] & b[121])^(a[146] & b[122])^(a[145] & b[123])^(a[144] & b[124])^(a[143] & b[125])^(a[142] & b[126])^(a[141] & b[127])^(a[140] & b[128])^(a[139] & b[129])^(a[138] & b[130])^(a[137] & b[131])^(a[136] & b[132])^(a[135] & b[133])^(a[134] & b[134])^(a[133] & b[135])^(a[132] & b[136])^(a[131] & b[137])^(a[130] & b[138])^(a[129] & b[139])^(a[128] & b[140])^(a[127] & b[141])^(a[126] & b[142])^(a[125] & b[143])^(a[124] & b[144])^(a[123] & b[145])^(a[122] & b[146])^(a[121] & b[147])^(a[120] & b[148])^(a[119] & b[149])^(a[118] & b[150])^(a[117] & b[151])^(a[116] & b[152])^(a[115] & b[153])^(a[114] & b[154])^(a[113] & b[155])^(a[112] & b[156])^(a[111] & b[157])^(a[110] & b[158])^(a[109] & b[159])^(a[108] & b[160])^(a[107] & b[161])^(a[106] & b[162]);
assign y[269] = (a[162] & b[107])^(a[161] & b[108])^(a[160] & b[109])^(a[159] & b[110])^(a[158] & b[111])^(a[157] & b[112])^(a[156] & b[113])^(a[155] & b[114])^(a[154] & b[115])^(a[153] & b[116])^(a[152] & b[117])^(a[151] & b[118])^(a[150] & b[119])^(a[149] & b[120])^(a[148] & b[121])^(a[147] & b[122])^(a[146] & b[123])^(a[145] & b[124])^(a[144] & b[125])^(a[143] & b[126])^(a[142] & b[127])^(a[141] & b[128])^(a[140] & b[129])^(a[139] & b[130])^(a[138] & b[131])^(a[137] & b[132])^(a[136] & b[133])^(a[135] & b[134])^(a[134] & b[135])^(a[133] & b[136])^(a[132] & b[137])^(a[131] & b[138])^(a[130] & b[139])^(a[129] & b[140])^(a[128] & b[141])^(a[127] & b[142])^(a[126] & b[143])^(a[125] & b[144])^(a[124] & b[145])^(a[123] & b[146])^(a[122] & b[147])^(a[121] & b[148])^(a[120] & b[149])^(a[119] & b[150])^(a[118] & b[151])^(a[117] & b[152])^(a[116] & b[153])^(a[115] & b[154])^(a[114] & b[155])^(a[113] & b[156])^(a[112] & b[157])^(a[111] & b[158])^(a[110] & b[159])^(a[109] & b[160])^(a[108] & b[161])^(a[107] & b[162]);
assign y[270] = (a[162] & b[108])^(a[161] & b[109])^(a[160] & b[110])^(a[159] & b[111])^(a[158] & b[112])^(a[157] & b[113])^(a[156] & b[114])^(a[155] & b[115])^(a[154] & b[116])^(a[153] & b[117])^(a[152] & b[118])^(a[151] & b[119])^(a[150] & b[120])^(a[149] & b[121])^(a[148] & b[122])^(a[147] & b[123])^(a[146] & b[124])^(a[145] & b[125])^(a[144] & b[126])^(a[143] & b[127])^(a[142] & b[128])^(a[141] & b[129])^(a[140] & b[130])^(a[139] & b[131])^(a[138] & b[132])^(a[137] & b[133])^(a[136] & b[134])^(a[135] & b[135])^(a[134] & b[136])^(a[133] & b[137])^(a[132] & b[138])^(a[131] & b[139])^(a[130] & b[140])^(a[129] & b[141])^(a[128] & b[142])^(a[127] & b[143])^(a[126] & b[144])^(a[125] & b[145])^(a[124] & b[146])^(a[123] & b[147])^(a[122] & b[148])^(a[121] & b[149])^(a[120] & b[150])^(a[119] & b[151])^(a[118] & b[152])^(a[117] & b[153])^(a[116] & b[154])^(a[115] & b[155])^(a[114] & b[156])^(a[113] & b[157])^(a[112] & b[158])^(a[111] & b[159])^(a[110] & b[160])^(a[109] & b[161])^(a[108] & b[162]);
assign y[271] = (a[162] & b[109])^(a[161] & b[110])^(a[160] & b[111])^(a[159] & b[112])^(a[158] & b[113])^(a[157] & b[114])^(a[156] & b[115])^(a[155] & b[116])^(a[154] & b[117])^(a[153] & b[118])^(a[152] & b[119])^(a[151] & b[120])^(a[150] & b[121])^(a[149] & b[122])^(a[148] & b[123])^(a[147] & b[124])^(a[146] & b[125])^(a[145] & b[126])^(a[144] & b[127])^(a[143] & b[128])^(a[142] & b[129])^(a[141] & b[130])^(a[140] & b[131])^(a[139] & b[132])^(a[138] & b[133])^(a[137] & b[134])^(a[136] & b[135])^(a[135] & b[136])^(a[134] & b[137])^(a[133] & b[138])^(a[132] & b[139])^(a[131] & b[140])^(a[130] & b[141])^(a[129] & b[142])^(a[128] & b[143])^(a[127] & b[144])^(a[126] & b[145])^(a[125] & b[146])^(a[124] & b[147])^(a[123] & b[148])^(a[122] & b[149])^(a[121] & b[150])^(a[120] & b[151])^(a[119] & b[152])^(a[118] & b[153])^(a[117] & b[154])^(a[116] & b[155])^(a[115] & b[156])^(a[114] & b[157])^(a[113] & b[158])^(a[112] & b[159])^(a[111] & b[160])^(a[110] & b[161])^(a[109] & b[162]);
assign y[272] = (a[162] & b[110])^(a[161] & b[111])^(a[160] & b[112])^(a[159] & b[113])^(a[158] & b[114])^(a[157] & b[115])^(a[156] & b[116])^(a[155] & b[117])^(a[154] & b[118])^(a[153] & b[119])^(a[152] & b[120])^(a[151] & b[121])^(a[150] & b[122])^(a[149] & b[123])^(a[148] & b[124])^(a[147] & b[125])^(a[146] & b[126])^(a[145] & b[127])^(a[144] & b[128])^(a[143] & b[129])^(a[142] & b[130])^(a[141] & b[131])^(a[140] & b[132])^(a[139] & b[133])^(a[138] & b[134])^(a[137] & b[135])^(a[136] & b[136])^(a[135] & b[137])^(a[134] & b[138])^(a[133] & b[139])^(a[132] & b[140])^(a[131] & b[141])^(a[130] & b[142])^(a[129] & b[143])^(a[128] & b[144])^(a[127] & b[145])^(a[126] & b[146])^(a[125] & b[147])^(a[124] & b[148])^(a[123] & b[149])^(a[122] & b[150])^(a[121] & b[151])^(a[120] & b[152])^(a[119] & b[153])^(a[118] & b[154])^(a[117] & b[155])^(a[116] & b[156])^(a[115] & b[157])^(a[114] & b[158])^(a[113] & b[159])^(a[112] & b[160])^(a[111] & b[161])^(a[110] & b[162]);
assign y[273] = (a[162] & b[111])^(a[161] & b[112])^(a[160] & b[113])^(a[159] & b[114])^(a[158] & b[115])^(a[157] & b[116])^(a[156] & b[117])^(a[155] & b[118])^(a[154] & b[119])^(a[153] & b[120])^(a[152] & b[121])^(a[151] & b[122])^(a[150] & b[123])^(a[149] & b[124])^(a[148] & b[125])^(a[147] & b[126])^(a[146] & b[127])^(a[145] & b[128])^(a[144] & b[129])^(a[143] & b[130])^(a[142] & b[131])^(a[141] & b[132])^(a[140] & b[133])^(a[139] & b[134])^(a[138] & b[135])^(a[137] & b[136])^(a[136] & b[137])^(a[135] & b[138])^(a[134] & b[139])^(a[133] & b[140])^(a[132] & b[141])^(a[131] & b[142])^(a[130] & b[143])^(a[129] & b[144])^(a[128] & b[145])^(a[127] & b[146])^(a[126] & b[147])^(a[125] & b[148])^(a[124] & b[149])^(a[123] & b[150])^(a[122] & b[151])^(a[121] & b[152])^(a[120] & b[153])^(a[119] & b[154])^(a[118] & b[155])^(a[117] & b[156])^(a[116] & b[157])^(a[115] & b[158])^(a[114] & b[159])^(a[113] & b[160])^(a[112] & b[161])^(a[111] & b[162]);
assign y[274] = (a[162] & b[112])^(a[161] & b[113])^(a[160] & b[114])^(a[159] & b[115])^(a[158] & b[116])^(a[157] & b[117])^(a[156] & b[118])^(a[155] & b[119])^(a[154] & b[120])^(a[153] & b[121])^(a[152] & b[122])^(a[151] & b[123])^(a[150] & b[124])^(a[149] & b[125])^(a[148] & b[126])^(a[147] & b[127])^(a[146] & b[128])^(a[145] & b[129])^(a[144] & b[130])^(a[143] & b[131])^(a[142] & b[132])^(a[141] & b[133])^(a[140] & b[134])^(a[139] & b[135])^(a[138] & b[136])^(a[137] & b[137])^(a[136] & b[138])^(a[135] & b[139])^(a[134] & b[140])^(a[133] & b[141])^(a[132] & b[142])^(a[131] & b[143])^(a[130] & b[144])^(a[129] & b[145])^(a[128] & b[146])^(a[127] & b[147])^(a[126] & b[148])^(a[125] & b[149])^(a[124] & b[150])^(a[123] & b[151])^(a[122] & b[152])^(a[121] & b[153])^(a[120] & b[154])^(a[119] & b[155])^(a[118] & b[156])^(a[117] & b[157])^(a[116] & b[158])^(a[115] & b[159])^(a[114] & b[160])^(a[113] & b[161])^(a[112] & b[162]);
assign y[275] = (a[162] & b[113])^(a[161] & b[114])^(a[160] & b[115])^(a[159] & b[116])^(a[158] & b[117])^(a[157] & b[118])^(a[156] & b[119])^(a[155] & b[120])^(a[154] & b[121])^(a[153] & b[122])^(a[152] & b[123])^(a[151] & b[124])^(a[150] & b[125])^(a[149] & b[126])^(a[148] & b[127])^(a[147] & b[128])^(a[146] & b[129])^(a[145] & b[130])^(a[144] & b[131])^(a[143] & b[132])^(a[142] & b[133])^(a[141] & b[134])^(a[140] & b[135])^(a[139] & b[136])^(a[138] & b[137])^(a[137] & b[138])^(a[136] & b[139])^(a[135] & b[140])^(a[134] & b[141])^(a[133] & b[142])^(a[132] & b[143])^(a[131] & b[144])^(a[130] & b[145])^(a[129] & b[146])^(a[128] & b[147])^(a[127] & b[148])^(a[126] & b[149])^(a[125] & b[150])^(a[124] & b[151])^(a[123] & b[152])^(a[122] & b[153])^(a[121] & b[154])^(a[120] & b[155])^(a[119] & b[156])^(a[118] & b[157])^(a[117] & b[158])^(a[116] & b[159])^(a[115] & b[160])^(a[114] & b[161])^(a[113] & b[162]);
assign y[276] = (a[162] & b[114])^(a[161] & b[115])^(a[160] & b[116])^(a[159] & b[117])^(a[158] & b[118])^(a[157] & b[119])^(a[156] & b[120])^(a[155] & b[121])^(a[154] & b[122])^(a[153] & b[123])^(a[152] & b[124])^(a[151] & b[125])^(a[150] & b[126])^(a[149] & b[127])^(a[148] & b[128])^(a[147] & b[129])^(a[146] & b[130])^(a[145] & b[131])^(a[144] & b[132])^(a[143] & b[133])^(a[142] & b[134])^(a[141] & b[135])^(a[140] & b[136])^(a[139] & b[137])^(a[138] & b[138])^(a[137] & b[139])^(a[136] & b[140])^(a[135] & b[141])^(a[134] & b[142])^(a[133] & b[143])^(a[132] & b[144])^(a[131] & b[145])^(a[130] & b[146])^(a[129] & b[147])^(a[128] & b[148])^(a[127] & b[149])^(a[126] & b[150])^(a[125] & b[151])^(a[124] & b[152])^(a[123] & b[153])^(a[122] & b[154])^(a[121] & b[155])^(a[120] & b[156])^(a[119] & b[157])^(a[118] & b[158])^(a[117] & b[159])^(a[116] & b[160])^(a[115] & b[161])^(a[114] & b[162]);
assign y[277] = (a[162] & b[115])^(a[161] & b[116])^(a[160] & b[117])^(a[159] & b[118])^(a[158] & b[119])^(a[157] & b[120])^(a[156] & b[121])^(a[155] & b[122])^(a[154] & b[123])^(a[153] & b[124])^(a[152] & b[125])^(a[151] & b[126])^(a[150] & b[127])^(a[149] & b[128])^(a[148] & b[129])^(a[147] & b[130])^(a[146] & b[131])^(a[145] & b[132])^(a[144] & b[133])^(a[143] & b[134])^(a[142] & b[135])^(a[141] & b[136])^(a[140] & b[137])^(a[139] & b[138])^(a[138] & b[139])^(a[137] & b[140])^(a[136] & b[141])^(a[135] & b[142])^(a[134] & b[143])^(a[133] & b[144])^(a[132] & b[145])^(a[131] & b[146])^(a[130] & b[147])^(a[129] & b[148])^(a[128] & b[149])^(a[127] & b[150])^(a[126] & b[151])^(a[125] & b[152])^(a[124] & b[153])^(a[123] & b[154])^(a[122] & b[155])^(a[121] & b[156])^(a[120] & b[157])^(a[119] & b[158])^(a[118] & b[159])^(a[117] & b[160])^(a[116] & b[161])^(a[115] & b[162]);
assign y[278] = (a[162] & b[116])^(a[161] & b[117])^(a[160] & b[118])^(a[159] & b[119])^(a[158] & b[120])^(a[157] & b[121])^(a[156] & b[122])^(a[155] & b[123])^(a[154] & b[124])^(a[153] & b[125])^(a[152] & b[126])^(a[151] & b[127])^(a[150] & b[128])^(a[149] & b[129])^(a[148] & b[130])^(a[147] & b[131])^(a[146] & b[132])^(a[145] & b[133])^(a[144] & b[134])^(a[143] & b[135])^(a[142] & b[136])^(a[141] & b[137])^(a[140] & b[138])^(a[139] & b[139])^(a[138] & b[140])^(a[137] & b[141])^(a[136] & b[142])^(a[135] & b[143])^(a[134] & b[144])^(a[133] & b[145])^(a[132] & b[146])^(a[131] & b[147])^(a[130] & b[148])^(a[129] & b[149])^(a[128] & b[150])^(a[127] & b[151])^(a[126] & b[152])^(a[125] & b[153])^(a[124] & b[154])^(a[123] & b[155])^(a[122] & b[156])^(a[121] & b[157])^(a[120] & b[158])^(a[119] & b[159])^(a[118] & b[160])^(a[117] & b[161])^(a[116] & b[162]);
assign y[279] = (a[162] & b[117])^(a[161] & b[118])^(a[160] & b[119])^(a[159] & b[120])^(a[158] & b[121])^(a[157] & b[122])^(a[156] & b[123])^(a[155] & b[124])^(a[154] & b[125])^(a[153] & b[126])^(a[152] & b[127])^(a[151] & b[128])^(a[150] & b[129])^(a[149] & b[130])^(a[148] & b[131])^(a[147] & b[132])^(a[146] & b[133])^(a[145] & b[134])^(a[144] & b[135])^(a[143] & b[136])^(a[142] & b[137])^(a[141] & b[138])^(a[140] & b[139])^(a[139] & b[140])^(a[138] & b[141])^(a[137] & b[142])^(a[136] & b[143])^(a[135] & b[144])^(a[134] & b[145])^(a[133] & b[146])^(a[132] & b[147])^(a[131] & b[148])^(a[130] & b[149])^(a[129] & b[150])^(a[128] & b[151])^(a[127] & b[152])^(a[126] & b[153])^(a[125] & b[154])^(a[124] & b[155])^(a[123] & b[156])^(a[122] & b[157])^(a[121] & b[158])^(a[120] & b[159])^(a[119] & b[160])^(a[118] & b[161])^(a[117] & b[162]);
assign y[280] = (a[162] & b[118])^(a[161] & b[119])^(a[160] & b[120])^(a[159] & b[121])^(a[158] & b[122])^(a[157] & b[123])^(a[156] & b[124])^(a[155] & b[125])^(a[154] & b[126])^(a[153] & b[127])^(a[152] & b[128])^(a[151] & b[129])^(a[150] & b[130])^(a[149] & b[131])^(a[148] & b[132])^(a[147] & b[133])^(a[146] & b[134])^(a[145] & b[135])^(a[144] & b[136])^(a[143] & b[137])^(a[142] & b[138])^(a[141] & b[139])^(a[140] & b[140])^(a[139] & b[141])^(a[138] & b[142])^(a[137] & b[143])^(a[136] & b[144])^(a[135] & b[145])^(a[134] & b[146])^(a[133] & b[147])^(a[132] & b[148])^(a[131] & b[149])^(a[130] & b[150])^(a[129] & b[151])^(a[128] & b[152])^(a[127] & b[153])^(a[126] & b[154])^(a[125] & b[155])^(a[124] & b[156])^(a[123] & b[157])^(a[122] & b[158])^(a[121] & b[159])^(a[120] & b[160])^(a[119] & b[161])^(a[118] & b[162]);
assign y[281] = (a[162] & b[119])^(a[161] & b[120])^(a[160] & b[121])^(a[159] & b[122])^(a[158] & b[123])^(a[157] & b[124])^(a[156] & b[125])^(a[155] & b[126])^(a[154] & b[127])^(a[153] & b[128])^(a[152] & b[129])^(a[151] & b[130])^(a[150] & b[131])^(a[149] & b[132])^(a[148] & b[133])^(a[147] & b[134])^(a[146] & b[135])^(a[145] & b[136])^(a[144] & b[137])^(a[143] & b[138])^(a[142] & b[139])^(a[141] & b[140])^(a[140] & b[141])^(a[139] & b[142])^(a[138] & b[143])^(a[137] & b[144])^(a[136] & b[145])^(a[135] & b[146])^(a[134] & b[147])^(a[133] & b[148])^(a[132] & b[149])^(a[131] & b[150])^(a[130] & b[151])^(a[129] & b[152])^(a[128] & b[153])^(a[127] & b[154])^(a[126] & b[155])^(a[125] & b[156])^(a[124] & b[157])^(a[123] & b[158])^(a[122] & b[159])^(a[121] & b[160])^(a[120] & b[161])^(a[119] & b[162]);
assign y[282] = (a[162] & b[120])^(a[161] & b[121])^(a[160] & b[122])^(a[159] & b[123])^(a[158] & b[124])^(a[157] & b[125])^(a[156] & b[126])^(a[155] & b[127])^(a[154] & b[128])^(a[153] & b[129])^(a[152] & b[130])^(a[151] & b[131])^(a[150] & b[132])^(a[149] & b[133])^(a[148] & b[134])^(a[147] & b[135])^(a[146] & b[136])^(a[145] & b[137])^(a[144] & b[138])^(a[143] & b[139])^(a[142] & b[140])^(a[141] & b[141])^(a[140] & b[142])^(a[139] & b[143])^(a[138] & b[144])^(a[137] & b[145])^(a[136] & b[146])^(a[135] & b[147])^(a[134] & b[148])^(a[133] & b[149])^(a[132] & b[150])^(a[131] & b[151])^(a[130] & b[152])^(a[129] & b[153])^(a[128] & b[154])^(a[127] & b[155])^(a[126] & b[156])^(a[125] & b[157])^(a[124] & b[158])^(a[123] & b[159])^(a[122] & b[160])^(a[121] & b[161])^(a[120] & b[162]);
assign y[283] = (a[162] & b[121])^(a[161] & b[122])^(a[160] & b[123])^(a[159] & b[124])^(a[158] & b[125])^(a[157] & b[126])^(a[156] & b[127])^(a[155] & b[128])^(a[154] & b[129])^(a[153] & b[130])^(a[152] & b[131])^(a[151] & b[132])^(a[150] & b[133])^(a[149] & b[134])^(a[148] & b[135])^(a[147] & b[136])^(a[146] & b[137])^(a[145] & b[138])^(a[144] & b[139])^(a[143] & b[140])^(a[142] & b[141])^(a[141] & b[142])^(a[140] & b[143])^(a[139] & b[144])^(a[138] & b[145])^(a[137] & b[146])^(a[136] & b[147])^(a[135] & b[148])^(a[134] & b[149])^(a[133] & b[150])^(a[132] & b[151])^(a[131] & b[152])^(a[130] & b[153])^(a[129] & b[154])^(a[128] & b[155])^(a[127] & b[156])^(a[126] & b[157])^(a[125] & b[158])^(a[124] & b[159])^(a[123] & b[160])^(a[122] & b[161])^(a[121] & b[162]);
assign y[284] = (a[162] & b[122])^(a[161] & b[123])^(a[160] & b[124])^(a[159] & b[125])^(a[158] & b[126])^(a[157] & b[127])^(a[156] & b[128])^(a[155] & b[129])^(a[154] & b[130])^(a[153] & b[131])^(a[152] & b[132])^(a[151] & b[133])^(a[150] & b[134])^(a[149] & b[135])^(a[148] & b[136])^(a[147] & b[137])^(a[146] & b[138])^(a[145] & b[139])^(a[144] & b[140])^(a[143] & b[141])^(a[142] & b[142])^(a[141] & b[143])^(a[140] & b[144])^(a[139] & b[145])^(a[138] & b[146])^(a[137] & b[147])^(a[136] & b[148])^(a[135] & b[149])^(a[134] & b[150])^(a[133] & b[151])^(a[132] & b[152])^(a[131] & b[153])^(a[130] & b[154])^(a[129] & b[155])^(a[128] & b[156])^(a[127] & b[157])^(a[126] & b[158])^(a[125] & b[159])^(a[124] & b[160])^(a[123] & b[161])^(a[122] & b[162]);
assign y[285] = (a[162] & b[123])^(a[161] & b[124])^(a[160] & b[125])^(a[159] & b[126])^(a[158] & b[127])^(a[157] & b[128])^(a[156] & b[129])^(a[155] & b[130])^(a[154] & b[131])^(a[153] & b[132])^(a[152] & b[133])^(a[151] & b[134])^(a[150] & b[135])^(a[149] & b[136])^(a[148] & b[137])^(a[147] & b[138])^(a[146] & b[139])^(a[145] & b[140])^(a[144] & b[141])^(a[143] & b[142])^(a[142] & b[143])^(a[141] & b[144])^(a[140] & b[145])^(a[139] & b[146])^(a[138] & b[147])^(a[137] & b[148])^(a[136] & b[149])^(a[135] & b[150])^(a[134] & b[151])^(a[133] & b[152])^(a[132] & b[153])^(a[131] & b[154])^(a[130] & b[155])^(a[129] & b[156])^(a[128] & b[157])^(a[127] & b[158])^(a[126] & b[159])^(a[125] & b[160])^(a[124] & b[161])^(a[123] & b[162]);
assign y[286] = (a[162] & b[124])^(a[161] & b[125])^(a[160] & b[126])^(a[159] & b[127])^(a[158] & b[128])^(a[157] & b[129])^(a[156] & b[130])^(a[155] & b[131])^(a[154] & b[132])^(a[153] & b[133])^(a[152] & b[134])^(a[151] & b[135])^(a[150] & b[136])^(a[149] & b[137])^(a[148] & b[138])^(a[147] & b[139])^(a[146] & b[140])^(a[145] & b[141])^(a[144] & b[142])^(a[143] & b[143])^(a[142] & b[144])^(a[141] & b[145])^(a[140] & b[146])^(a[139] & b[147])^(a[138] & b[148])^(a[137] & b[149])^(a[136] & b[150])^(a[135] & b[151])^(a[134] & b[152])^(a[133] & b[153])^(a[132] & b[154])^(a[131] & b[155])^(a[130] & b[156])^(a[129] & b[157])^(a[128] & b[158])^(a[127] & b[159])^(a[126] & b[160])^(a[125] & b[161])^(a[124] & b[162]);
assign y[287] = (a[162] & b[125])^(a[161] & b[126])^(a[160] & b[127])^(a[159] & b[128])^(a[158] & b[129])^(a[157] & b[130])^(a[156] & b[131])^(a[155] & b[132])^(a[154] & b[133])^(a[153] & b[134])^(a[152] & b[135])^(a[151] & b[136])^(a[150] & b[137])^(a[149] & b[138])^(a[148] & b[139])^(a[147] & b[140])^(a[146] & b[141])^(a[145] & b[142])^(a[144] & b[143])^(a[143] & b[144])^(a[142] & b[145])^(a[141] & b[146])^(a[140] & b[147])^(a[139] & b[148])^(a[138] & b[149])^(a[137] & b[150])^(a[136] & b[151])^(a[135] & b[152])^(a[134] & b[153])^(a[133] & b[154])^(a[132] & b[155])^(a[131] & b[156])^(a[130] & b[157])^(a[129] & b[158])^(a[128] & b[159])^(a[127] & b[160])^(a[126] & b[161])^(a[125] & b[162]);
assign y[288] = (a[162] & b[126])^(a[161] & b[127])^(a[160] & b[128])^(a[159] & b[129])^(a[158] & b[130])^(a[157] & b[131])^(a[156] & b[132])^(a[155] & b[133])^(a[154] & b[134])^(a[153] & b[135])^(a[152] & b[136])^(a[151] & b[137])^(a[150] & b[138])^(a[149] & b[139])^(a[148] & b[140])^(a[147] & b[141])^(a[146] & b[142])^(a[145] & b[143])^(a[144] & b[144])^(a[143] & b[145])^(a[142] & b[146])^(a[141] & b[147])^(a[140] & b[148])^(a[139] & b[149])^(a[138] & b[150])^(a[137] & b[151])^(a[136] & b[152])^(a[135] & b[153])^(a[134] & b[154])^(a[133] & b[155])^(a[132] & b[156])^(a[131] & b[157])^(a[130] & b[158])^(a[129] & b[159])^(a[128] & b[160])^(a[127] & b[161])^(a[126] & b[162]);
assign y[289] = (a[162] & b[127])^(a[161] & b[128])^(a[160] & b[129])^(a[159] & b[130])^(a[158] & b[131])^(a[157] & b[132])^(a[156] & b[133])^(a[155] & b[134])^(a[154] & b[135])^(a[153] & b[136])^(a[152] & b[137])^(a[151] & b[138])^(a[150] & b[139])^(a[149] & b[140])^(a[148] & b[141])^(a[147] & b[142])^(a[146] & b[143])^(a[145] & b[144])^(a[144] & b[145])^(a[143] & b[146])^(a[142] & b[147])^(a[141] & b[148])^(a[140] & b[149])^(a[139] & b[150])^(a[138] & b[151])^(a[137] & b[152])^(a[136] & b[153])^(a[135] & b[154])^(a[134] & b[155])^(a[133] & b[156])^(a[132] & b[157])^(a[131] & b[158])^(a[130] & b[159])^(a[129] & b[160])^(a[128] & b[161])^(a[127] & b[162]);
assign y[290] = (a[162] & b[128])^(a[161] & b[129])^(a[160] & b[130])^(a[159] & b[131])^(a[158] & b[132])^(a[157] & b[133])^(a[156] & b[134])^(a[155] & b[135])^(a[154] & b[136])^(a[153] & b[137])^(a[152] & b[138])^(a[151] & b[139])^(a[150] & b[140])^(a[149] & b[141])^(a[148] & b[142])^(a[147] & b[143])^(a[146] & b[144])^(a[145] & b[145])^(a[144] & b[146])^(a[143] & b[147])^(a[142] & b[148])^(a[141] & b[149])^(a[140] & b[150])^(a[139] & b[151])^(a[138] & b[152])^(a[137] & b[153])^(a[136] & b[154])^(a[135] & b[155])^(a[134] & b[156])^(a[133] & b[157])^(a[132] & b[158])^(a[131] & b[159])^(a[130] & b[160])^(a[129] & b[161])^(a[128] & b[162]);
assign y[291] = (a[162] & b[129])^(a[161] & b[130])^(a[160] & b[131])^(a[159] & b[132])^(a[158] & b[133])^(a[157] & b[134])^(a[156] & b[135])^(a[155] & b[136])^(a[154] & b[137])^(a[153] & b[138])^(a[152] & b[139])^(a[151] & b[140])^(a[150] & b[141])^(a[149] & b[142])^(a[148] & b[143])^(a[147] & b[144])^(a[146] & b[145])^(a[145] & b[146])^(a[144] & b[147])^(a[143] & b[148])^(a[142] & b[149])^(a[141] & b[150])^(a[140] & b[151])^(a[139] & b[152])^(a[138] & b[153])^(a[137] & b[154])^(a[136] & b[155])^(a[135] & b[156])^(a[134] & b[157])^(a[133] & b[158])^(a[132] & b[159])^(a[131] & b[160])^(a[130] & b[161])^(a[129] & b[162]);
assign y[292] = (a[162] & b[130])^(a[161] & b[131])^(a[160] & b[132])^(a[159] & b[133])^(a[158] & b[134])^(a[157] & b[135])^(a[156] & b[136])^(a[155] & b[137])^(a[154] & b[138])^(a[153] & b[139])^(a[152] & b[140])^(a[151] & b[141])^(a[150] & b[142])^(a[149] & b[143])^(a[148] & b[144])^(a[147] & b[145])^(a[146] & b[146])^(a[145] & b[147])^(a[144] & b[148])^(a[143] & b[149])^(a[142] & b[150])^(a[141] & b[151])^(a[140] & b[152])^(a[139] & b[153])^(a[138] & b[154])^(a[137] & b[155])^(a[136] & b[156])^(a[135] & b[157])^(a[134] & b[158])^(a[133] & b[159])^(a[132] & b[160])^(a[131] & b[161])^(a[130] & b[162]);
assign y[293] = (a[162] & b[131])^(a[161] & b[132])^(a[160] & b[133])^(a[159] & b[134])^(a[158] & b[135])^(a[157] & b[136])^(a[156] & b[137])^(a[155] & b[138])^(a[154] & b[139])^(a[153] & b[140])^(a[152] & b[141])^(a[151] & b[142])^(a[150] & b[143])^(a[149] & b[144])^(a[148] & b[145])^(a[147] & b[146])^(a[146] & b[147])^(a[145] & b[148])^(a[144] & b[149])^(a[143] & b[150])^(a[142] & b[151])^(a[141] & b[152])^(a[140] & b[153])^(a[139] & b[154])^(a[138] & b[155])^(a[137] & b[156])^(a[136] & b[157])^(a[135] & b[158])^(a[134] & b[159])^(a[133] & b[160])^(a[132] & b[161])^(a[131] & b[162]);
assign y[294] = (a[162] & b[132])^(a[161] & b[133])^(a[160] & b[134])^(a[159] & b[135])^(a[158] & b[136])^(a[157] & b[137])^(a[156] & b[138])^(a[155] & b[139])^(a[154] & b[140])^(a[153] & b[141])^(a[152] & b[142])^(a[151] & b[143])^(a[150] & b[144])^(a[149] & b[145])^(a[148] & b[146])^(a[147] & b[147])^(a[146] & b[148])^(a[145] & b[149])^(a[144] & b[150])^(a[143] & b[151])^(a[142] & b[152])^(a[141] & b[153])^(a[140] & b[154])^(a[139] & b[155])^(a[138] & b[156])^(a[137] & b[157])^(a[136] & b[158])^(a[135] & b[159])^(a[134] & b[160])^(a[133] & b[161])^(a[132] & b[162]);
assign y[295] = (a[162] & b[133])^(a[161] & b[134])^(a[160] & b[135])^(a[159] & b[136])^(a[158] & b[137])^(a[157] & b[138])^(a[156] & b[139])^(a[155] & b[140])^(a[154] & b[141])^(a[153] & b[142])^(a[152] & b[143])^(a[151] & b[144])^(a[150] & b[145])^(a[149] & b[146])^(a[148] & b[147])^(a[147] & b[148])^(a[146] & b[149])^(a[145] & b[150])^(a[144] & b[151])^(a[143] & b[152])^(a[142] & b[153])^(a[141] & b[154])^(a[140] & b[155])^(a[139] & b[156])^(a[138] & b[157])^(a[137] & b[158])^(a[136] & b[159])^(a[135] & b[160])^(a[134] & b[161])^(a[133] & b[162]);
assign y[296] = (a[162] & b[134])^(a[161] & b[135])^(a[160] & b[136])^(a[159] & b[137])^(a[158] & b[138])^(a[157] & b[139])^(a[156] & b[140])^(a[155] & b[141])^(a[154] & b[142])^(a[153] & b[143])^(a[152] & b[144])^(a[151] & b[145])^(a[150] & b[146])^(a[149] & b[147])^(a[148] & b[148])^(a[147] & b[149])^(a[146] & b[150])^(a[145] & b[151])^(a[144] & b[152])^(a[143] & b[153])^(a[142] & b[154])^(a[141] & b[155])^(a[140] & b[156])^(a[139] & b[157])^(a[138] & b[158])^(a[137] & b[159])^(a[136] & b[160])^(a[135] & b[161])^(a[134] & b[162]);
assign y[297] = (a[162] & b[135])^(a[161] & b[136])^(a[160] & b[137])^(a[159] & b[138])^(a[158] & b[139])^(a[157] & b[140])^(a[156] & b[141])^(a[155] & b[142])^(a[154] & b[143])^(a[153] & b[144])^(a[152] & b[145])^(a[151] & b[146])^(a[150] & b[147])^(a[149] & b[148])^(a[148] & b[149])^(a[147] & b[150])^(a[146] & b[151])^(a[145] & b[152])^(a[144] & b[153])^(a[143] & b[154])^(a[142] & b[155])^(a[141] & b[156])^(a[140] & b[157])^(a[139] & b[158])^(a[138] & b[159])^(a[137] & b[160])^(a[136] & b[161])^(a[135] & b[162]);
assign y[298] = (a[162] & b[136])^(a[161] & b[137])^(a[160] & b[138])^(a[159] & b[139])^(a[158] & b[140])^(a[157] & b[141])^(a[156] & b[142])^(a[155] & b[143])^(a[154] & b[144])^(a[153] & b[145])^(a[152] & b[146])^(a[151] & b[147])^(a[150] & b[148])^(a[149] & b[149])^(a[148] & b[150])^(a[147] & b[151])^(a[146] & b[152])^(a[145] & b[153])^(a[144] & b[154])^(a[143] & b[155])^(a[142] & b[156])^(a[141] & b[157])^(a[140] & b[158])^(a[139] & b[159])^(a[138] & b[160])^(a[137] & b[161])^(a[136] & b[162]);
assign y[299] = (a[162] & b[137])^(a[161] & b[138])^(a[160] & b[139])^(a[159] & b[140])^(a[158] & b[141])^(a[157] & b[142])^(a[156] & b[143])^(a[155] & b[144])^(a[154] & b[145])^(a[153] & b[146])^(a[152] & b[147])^(a[151] & b[148])^(a[150] & b[149])^(a[149] & b[150])^(a[148] & b[151])^(a[147] & b[152])^(a[146] & b[153])^(a[145] & b[154])^(a[144] & b[155])^(a[143] & b[156])^(a[142] & b[157])^(a[141] & b[158])^(a[140] & b[159])^(a[139] & b[160])^(a[138] & b[161])^(a[137] & b[162]);
assign y[300] = (a[162] & b[138])^(a[161] & b[139])^(a[160] & b[140])^(a[159] & b[141])^(a[158] & b[142])^(a[157] & b[143])^(a[156] & b[144])^(a[155] & b[145])^(a[154] & b[146])^(a[153] & b[147])^(a[152] & b[148])^(a[151] & b[149])^(a[150] & b[150])^(a[149] & b[151])^(a[148] & b[152])^(a[147] & b[153])^(a[146] & b[154])^(a[145] & b[155])^(a[144] & b[156])^(a[143] & b[157])^(a[142] & b[158])^(a[141] & b[159])^(a[140] & b[160])^(a[139] & b[161])^(a[138] & b[162]);
assign y[301] = (a[162] & b[139])^(a[161] & b[140])^(a[160] & b[141])^(a[159] & b[142])^(a[158] & b[143])^(a[157] & b[144])^(a[156] & b[145])^(a[155] & b[146])^(a[154] & b[147])^(a[153] & b[148])^(a[152] & b[149])^(a[151] & b[150])^(a[150] & b[151])^(a[149] & b[152])^(a[148] & b[153])^(a[147] & b[154])^(a[146] & b[155])^(a[145] & b[156])^(a[144] & b[157])^(a[143] & b[158])^(a[142] & b[159])^(a[141] & b[160])^(a[140] & b[161])^(a[139] & b[162]);
assign y[302] = (a[162] & b[140])^(a[161] & b[141])^(a[160] & b[142])^(a[159] & b[143])^(a[158] & b[144])^(a[157] & b[145])^(a[156] & b[146])^(a[155] & b[147])^(a[154] & b[148])^(a[153] & b[149])^(a[152] & b[150])^(a[151] & b[151])^(a[150] & b[152])^(a[149] & b[153])^(a[148] & b[154])^(a[147] & b[155])^(a[146] & b[156])^(a[145] & b[157])^(a[144] & b[158])^(a[143] & b[159])^(a[142] & b[160])^(a[141] & b[161])^(a[140] & b[162]);
assign y[303] = (a[162] & b[141])^(a[161] & b[142])^(a[160] & b[143])^(a[159] & b[144])^(a[158] & b[145])^(a[157] & b[146])^(a[156] & b[147])^(a[155] & b[148])^(a[154] & b[149])^(a[153] & b[150])^(a[152] & b[151])^(a[151] & b[152])^(a[150] & b[153])^(a[149] & b[154])^(a[148] & b[155])^(a[147] & b[156])^(a[146] & b[157])^(a[145] & b[158])^(a[144] & b[159])^(a[143] & b[160])^(a[142] & b[161])^(a[141] & b[162]);
assign y[304] = (a[162] & b[142])^(a[161] & b[143])^(a[160] & b[144])^(a[159] & b[145])^(a[158] & b[146])^(a[157] & b[147])^(a[156] & b[148])^(a[155] & b[149])^(a[154] & b[150])^(a[153] & b[151])^(a[152] & b[152])^(a[151] & b[153])^(a[150] & b[154])^(a[149] & b[155])^(a[148] & b[156])^(a[147] & b[157])^(a[146] & b[158])^(a[145] & b[159])^(a[144] & b[160])^(a[143] & b[161])^(a[142] & b[162]);
assign y[305] = (a[162] & b[143])^(a[161] & b[144])^(a[160] & b[145])^(a[159] & b[146])^(a[158] & b[147])^(a[157] & b[148])^(a[156] & b[149])^(a[155] & b[150])^(a[154] & b[151])^(a[153] & b[152])^(a[152] & b[153])^(a[151] & b[154])^(a[150] & b[155])^(a[149] & b[156])^(a[148] & b[157])^(a[147] & b[158])^(a[146] & b[159])^(a[145] & b[160])^(a[144] & b[161])^(a[143] & b[162]);
assign y[306] = (a[162] & b[144])^(a[161] & b[145])^(a[160] & b[146])^(a[159] & b[147])^(a[158] & b[148])^(a[157] & b[149])^(a[156] & b[150])^(a[155] & b[151])^(a[154] & b[152])^(a[153] & b[153])^(a[152] & b[154])^(a[151] & b[155])^(a[150] & b[156])^(a[149] & b[157])^(a[148] & b[158])^(a[147] & b[159])^(a[146] & b[160])^(a[145] & b[161])^(a[144] & b[162]);
assign y[307] = (a[162] & b[145])^(a[161] & b[146])^(a[160] & b[147])^(a[159] & b[148])^(a[158] & b[149])^(a[157] & b[150])^(a[156] & b[151])^(a[155] & b[152])^(a[154] & b[153])^(a[153] & b[154])^(a[152] & b[155])^(a[151] & b[156])^(a[150] & b[157])^(a[149] & b[158])^(a[148] & b[159])^(a[147] & b[160])^(a[146] & b[161])^(a[145] & b[162]);
assign y[308] = (a[162] & b[146])^(a[161] & b[147])^(a[160] & b[148])^(a[159] & b[149])^(a[158] & b[150])^(a[157] & b[151])^(a[156] & b[152])^(a[155] & b[153])^(a[154] & b[154])^(a[153] & b[155])^(a[152] & b[156])^(a[151] & b[157])^(a[150] & b[158])^(a[149] & b[159])^(a[148] & b[160])^(a[147] & b[161])^(a[146] & b[162]);
assign y[309] = (a[162] & b[147])^(a[161] & b[148])^(a[160] & b[149])^(a[159] & b[150])^(a[158] & b[151])^(a[157] & b[152])^(a[156] & b[153])^(a[155] & b[154])^(a[154] & b[155])^(a[153] & b[156])^(a[152] & b[157])^(a[151] & b[158])^(a[150] & b[159])^(a[149] & b[160])^(a[148] & b[161])^(a[147] & b[162]);
assign y[310] = (a[162] & b[148])^(a[161] & b[149])^(a[160] & b[150])^(a[159] & b[151])^(a[158] & b[152])^(a[157] & b[153])^(a[156] & b[154])^(a[155] & b[155])^(a[154] & b[156])^(a[153] & b[157])^(a[152] & b[158])^(a[151] & b[159])^(a[150] & b[160])^(a[149] & b[161])^(a[148] & b[162]);
assign y[311] = (a[162] & b[149])^(a[161] & b[150])^(a[160] & b[151])^(a[159] & b[152])^(a[158] & b[153])^(a[157] & b[154])^(a[156] & b[155])^(a[155] & b[156])^(a[154] & b[157])^(a[153] & b[158])^(a[152] & b[159])^(a[151] & b[160])^(a[150] & b[161])^(a[149] & b[162]);
assign y[312] = (a[162] & b[150])^(a[161] & b[151])^(a[160] & b[152])^(a[159] & b[153])^(a[158] & b[154])^(a[157] & b[155])^(a[156] & b[156])^(a[155] & b[157])^(a[154] & b[158])^(a[153] & b[159])^(a[152] & b[160])^(a[151] & b[161])^(a[150] & b[162]);
assign y[313] = (a[162] & b[151])^(a[161] & b[152])^(a[160] & b[153])^(a[159] & b[154])^(a[158] & b[155])^(a[157] & b[156])^(a[156] & b[157])^(a[155] & b[158])^(a[154] & b[159])^(a[153] & b[160])^(a[152] & b[161])^(a[151] & b[162]);
assign y[314] = (a[162] & b[152])^(a[161] & b[153])^(a[160] & b[154])^(a[159] & b[155])^(a[158] & b[156])^(a[157] & b[157])^(a[156] & b[158])^(a[155] & b[159])^(a[154] & b[160])^(a[153] & b[161])^(a[152] & b[162]);
assign y[315] = (a[162] & b[153])^(a[161] & b[154])^(a[160] & b[155])^(a[159] & b[156])^(a[158] & b[157])^(a[157] & b[158])^(a[156] & b[159])^(a[155] & b[160])^(a[154] & b[161])^(a[153] & b[162]);
assign y[316] = (a[162] & b[154])^(a[161] & b[155])^(a[160] & b[156])^(a[159] & b[157])^(a[158] & b[158])^(a[157] & b[159])^(a[156] & b[160])^(a[155] & b[161])^(a[154] & b[162]);
assign y[317] = (a[162] & b[155])^(a[161] & b[156])^(a[160] & b[157])^(a[159] & b[158])^(a[158] & b[159])^(a[157] & b[160])^(a[156] & b[161])^(a[155] & b[162]);
assign y[318] = (a[162] & b[156])^(a[161] & b[157])^(a[160] & b[158])^(a[159] & b[159])^(a[158] & b[160])^(a[157] & b[161])^(a[156] & b[162]);
assign y[319] = (a[162] & b[157])^(a[161] & b[158])^(a[160] & b[159])^(a[159] & b[160])^(a[158] & b[161])^(a[157] & b[162]);
assign y[320] = (a[162] & b[158])^(a[161] & b[159])^(a[160] & b[160])^(a[159] & b[161])^(a[158] & b[162]);
assign y[321] = (a[162] & b[159])^(a[161] & b[160])^(a[160] & b[161])^(a[159] & b[162]);
assign y[322] = (a[162] & b[160])^(a[161] & b[161])^(a[160] & b[162]);
assign y[323] = (a[162] & b[161])^(a[161] & b[162]);
assign y[324] = (a[162] & b[162]);


endmodule
